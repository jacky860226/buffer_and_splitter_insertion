module c5315(G1, G10, G100, G101, G102, G103, G104, G105, G106, G107, G108, G109, G11, G110, G111, G112, G113, G114, G115, G116, G117, G118, G119, G12, G120, G121, G122, G123, G124, G125, G126, G127, G128, G129, G13, G130, G131, G132, G133, G134, G135, G136, G137, G138, G139, G14, G140, G141, G142, G143, G144, G145, G146, G147, G148, G149, G15, G150, G151, G152, G153, G154, G155, G156, G157, G158, G159, G16, G160, G161, G162, G163, G164, G165, G166, G167, G168, G169, G17, G170, G171, G172, G173, G174, G175, G176, G177, G178, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G42, G43, G44, G45, G46, G47, G48, G49, G5, G50, G51, G5193, G5194, G5195, G5196, G5197, G5198, G5199, G52, G5200, G5201, G5202, G5203, G5204, G5205, G5206, G5207, G5208, G5209, G5210, G5211, G5212, G5213, G5214, G5215, G5216, G5217, G5218, G5219, G5220, G5221, G5222, G5223, G5224, G5225, G5226, G5227, G5228, G5229, G5230, G5231, G5232, G5233, G5234, G5235, G5236, G5237, G5238, G5239, G5240, G5241, G5242, G5243, G5244, G5245, G5246, G5247, G5248, G5249, G5250, G5251, G5252, G5253, G5254, G5255, G5256, G5257, G5258, G5259, G5260, G5261, G5262, G5263, G5264, G5265, G5266, G5267, G5268, G5269, G5270, G5271, G5272, G5273, G5274, G5275, G5276, G5277, G5278, G5279, G5280, G5281, G5282, G5283, G5284, G5285, G5286, G5287, G5288, G5289, G5290, G5291, G5292, G5293, G5294, G5295, G5296, G5297, G5298, G5299, G53, G5300, G5301, G5302, G5303, G5304, G5305, G5306, G5307, G5308, G5309, G5310, G5311, G5312, G5313, G5314, G5315, G54, G55, G56, G57, G58, G59, G6, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G7, G70, G71, G72, G73, G74, G75, G76, G77, G78, G79, G8, G80, G81, G82, G83, G84, G85, G86, G87, G88, G89, G9, G90, G91, G92, G93, G94, G95, G96, G97, G98, G99);
	wire new_net_5273;
	wire new_net_6137;
	wire new_net_6755;
	wire new_net_5485;
	wire new_net_7197;
	wire new_net_5730;
	wire new_net_6927;
	wire new_net_4677;
	wire new_net_6476;
	wire _0022_;
	wire _0232_;
	wire new_net_3041;
	wire new_net_1330;
	wire new_net_2256;
	wire _0946_;
	wire _0442_;
	wire new_net_287;
	wire new_net_323;
	wire _0736_;
	wire new_net_7011;
	wire new_net_7924;
	wire new_net_7844;
	wire new_net_6949;
	wire new_net_183;
	wire new_net_252;
	wire new_net_1364;
	wire new_net_3612;
	wire new_net_3908;
	wire new_net_4542;
	wire new_net_4611;
	wire new_net_4629;
	wire new_net_5104;
	wire new_net_6466;
	wire new_net_7449;
	wire new_net_7532;
	wire new_net_7780;
	wire new_net_5640;
	wire new_net_5803;
	wire _0023_;
	wire _0233_;
	wire new_net_1296;
	wire _0947_;
	wire _0443_;
	wire new_net_1644;
	wire new_net_3399;
	wire new_net_2439;
	wire new_net_1224;
	wire _0737_;
	wire new_net_6638;
	wire new_net_7556;
	wire new_net_7254;
	wire new_net_8207;
	wire new_net_7471;
	wire new_net_4536;
	wire new_net_6314;
	wire new_net_1465;
	wire new_net_1432;
	wire new_net_1501;
	wire new_net_1576;
	wire new_net_2018;
	wire new_net_2093;
	wire new_net_3869;
	wire new_net_3893;
	wire new_net_5402;
	wire new_net_6388;
	wire new_net_7571;
	wire new_net_7778;
	wire new_net_5222;
	wire new_net_4298;
	wire new_net_7776;
	wire _0024_;
	wire _0234_;
	wire _0444_;
	wire _0738_;
	wire new_net_2105;
	wire new_net_1262;
	wire new_net_2162;
	wire new_net_2463;
	wire new_net_2893;
	wire _0948_;
	wire new_net_8195;
	wire new_net_184;
	wire new_net_427;
	wire new_net_898;
	wire new_net_1904;
	wire new_net_3349;
	wire new_net_5647;
	wire new_net_6243;
	wire new_net_6341;
	wire new_net_6365;
	wire new_net_6669;
	wire new_net_8134;
	wire new_net_8266;
	wire _0235_;
	wire _0025_;
	wire _0739_;
	wire new_net_3576;
	wire new_net_1297;
	wire _0949_;
	wire _0445_;
	wire new_net_1645;
	wire new_net_1225;
	wire new_net_3926;
	wire new_net_5355;
	wire new_net_324;
	wire new_net_1331;
	wire new_net_1433;
	wire new_net_1466;
	wire new_net_2772;
	wire new_net_1502;
	wire new_net_3042;
	wire new_net_4167;
	wire new_net_4267;
	wire new_net_4291;
	wire new_net_4638;
	wire new_net_6274;
	wire new_net_6272;
	wire new_net_1716;
	wire _0950_;
	wire _0236_;
	wire _0026_;
	wire _0740_;
	wire new_net_1263;
	wire new_net_2401;
	wire new_net_2913;
	wire new_net_3613;
	wire new_net_253;
	wire new_net_6368;
	wire new_net_6830;
	wire new_net_185;
	wire new_net_218;
	wire new_net_428;
	wire new_net_1741;
	wire new_net_3362;
	wire new_net_3400;
	wire new_net_3655;
	wire new_net_899;
	wire new_net_4357;
	wire new_net_4652;
	wire new_net_7041;
	wire new_net_6629;
	wire new_net_5613;
	wire _0027_;
	wire _0237_;
	wire new_net_1226;
	wire _0741_;
	wire new_net_2773;
	wire new_net_1298;
	wire _0951_;
	wire new_net_1577;
	wire _0447_;
	wire new_net_2961;
	wire new_net_5988;
	wire new_net_7307;
	wire new_net_4165;
	wire new_net_8215;
	wire new_net_3828;
	wire new_net_4225;
	wire new_net_7936;
	wire new_net_289;
	wire new_net_325;
	wire new_net_1332;
	wire new_net_1434;
	wire new_net_1467;
	wire new_net_2523;
	wire new_net_2894;
	wire new_net_1503;
	wire new_net_2883;
	wire new_net_1878;
	wire new_net_6956;
	wire _0448_;
	wire _0742_;
	wire _0028_;
	wire _0238_;
	wire new_net_1264;
	wire new_net_2163;
	wire new_net_2524;
	wire new_net_2914;
	wire new_net_3350;
	wire _0952_;
	wire new_net_8002;
	wire new_net_4052;
	wire new_net_186;
	wire new_net_219;
	wire new_net_429;
	wire new_net_900;
	wire new_net_3577;
	wire new_net_1646;
	wire new_net_3927;
	wire new_net_3951;
	wire new_net_3966;
	wire new_net_5950;
	wire new_net_6860;
	wire new_net_5250;
	wire new_net_6442;
	wire new_net_8024;
	wire _0449_;
	wire _0743_;
	wire _0239_;
	wire _0029_;
	wire new_net_1227;
	wire new_net_2417;
	wire new_net_1762;
	wire new_net_3043;
	wire _0953_;
	wire new_net_1578;
	wire new_net_6882;
	wire new_net_6794;
	wire new_net_7828;
	wire new_net_6187;
	wire new_net_7511;
	wire new_net_290;
	wire new_net_326;
	wire new_net_1717;
	wire new_net_2078;
	wire new_net_1468;
	wire new_net_2104;
	wire new_net_1504;
	wire new_net_1540;
	wire new_net_3614;
	wire new_net_3910;
	wire new_net_6354;
	wire new_net_5624;
	wire new_net_7361;
	wire new_net_5400;
	wire new_net_1367;
	wire new_net_3401;
	wire _0954_;
	wire _0240_;
	wire _0030_;
	wire _0744_;
	wire new_net_2258;
	wire _0450_;
	wire new_net_4653;
	wire new_net_5626;
	wire new_net_4963;
	wire new_net_5061;
	wire new_net_5606;
	wire new_net_4942;
	wire new_net_1299;
	wire new_net_1647;
	wire new_net_1764;
	wire new_net_3871;
	wire new_net_3895;
	wire new_net_4525;
	wire new_net_5404;
	wire new_net_6390;
	wire new_net_6445;
	wire new_net_7338;
	wire new_net_7298;
	wire new_net_7671;
	wire new_net_5032;
	wire new_net_5206;
	wire new_net_7054;
	wire new_net_6976;
	wire new_net_6565;
	wire new_net_7642;
	wire new_net_5739;
	wire new_net_6936;
	wire _0955_;
	wire _0241_;
	wire _0031_;
	wire new_net_1228;
	wire new_net_1435;
	wire _0745_;
	wire new_net_2465;
	wire new_net_2895;
	wire _0451_;
	wire new_net_6692;
	wire new_net_6074;
	wire new_net_8177;
	wire new_net_6652;
	wire new_net_7149;
	wire new_net_5710;
	wire new_net_7944;
	wire new_net_3256;
	wire new_net_3657;
	wire new_net_255;
	wire new_net_1265;
	wire new_net_1718;
	wire new_net_1469;
	wire new_net_3351;
	wire new_net_1505;
	wire new_net_2915;
	wire new_net_1541;
	wire new_net_5103;
	wire new_net_7165;
	wire new_net_6384;
	wire new_net_6306;
	wire new_net_5817;
	wire _0452_;
	wire _0032_;
	wire _0242_;
	wire new_net_1368;
	wire new_net_901;
	wire new_net_187;
	wire _0746_;
	wire new_net_220;
	wire new_net_430;
	wire new_net_2164;
	wire new_net_5778;
	wire new_net_7391;
	wire new_net_4978;
	wire new_net_6406;
	wire new_net_8015;
	wire new_net_6323;
	wire new_net_1744;
	wire new_net_1300;
	wire new_net_1579;
	wire new_net_3044;
	wire new_net_4269;
	wire new_net_4293;
	wire new_net_4358;
	wire new_net_4845;
	wire new_net_7316;
	wire new_net_8137;
	wire new_net_7819;
	wire new_net_4257;
	wire new_net_7988;
	wire new_net_6178;
	wire new_net_6713;
	wire new_net_291;
	wire _0453_;
	wire _0747_;
	wire new_net_327;
	wire _0033_;
	wire new_net_2355;
	wire new_net_1229;
	wire new_net_1436;
	wire new_net_2403;
	wire _0243_;
	wire new_net_5524;
	wire new_net_5939;
	wire new_net_6345;
	wire new_net_6595;
	wire new_net_8126;
	wire new_net_4280;
	wire new_net_6106;
	wire new_net_256;
	wire new_net_1266;
	wire new_net_3257;
	wire new_net_3402;
	wire new_net_1470;
	wire new_net_1506;
	wire new_net_3595;
	wire new_net_4654;
	wire new_net_5129;
	wire new_net_5627;
	wire new_net_8054;
	wire new_net_6907;
	wire new_net_8091;
	wire new_net_7278;
	wire new_net_6905;
	wire new_net_6456;
	wire new_net_6454;
	wire _0454_;
	wire _0748_;
	wire _0034_;
	wire new_net_1369;
	wire new_net_1648;
	wire new_net_1821;
	wire new_net_3658;
	wire new_net_902;
	wire new_net_188;
	wire new_net_221;
	wire new_net_1908;
	wire new_net_7595;
	wire new_net_8246;
	wire new_net_7802;
	wire new_net_1301;
	wire new_net_1580;
	wire new_net_2896;
	wire new_net_6693;
	wire new_net_6820;
	wire new_net_6966;
	wire new_net_7670;
	wire new_net_7800;
	wire new_net_6065;
	wire new_net_6817;
	wire new_net_7851;
	wire new_net_3365;
	wire _0959_;
	wire _0035_;
	wire _0455_;
	wire new_net_292;
	wire new_net_2963;
	wire new_net_328;
	wire new_net_1230;
	wire new_net_1719;
	wire _0749_;
	wire new_net_5674;
	wire new_net_7895;
	wire new_net_7699;
	wire new_net_6292;
	wire new_net_8158;
	wire new_net_7866;
	wire new_net_7249;
	wire new_net_1817;
	wire new_net_1267;
	wire new_net_1471;
	wire new_net_3579;
	wire new_net_3929;
	wire new_net_3953;
	wire new_net_3968;
	wire new_net_4169;
	wire new_net_5952;
	wire new_net_6797;
	wire new_net_7957;
	wire new_net_6142;
	wire new_net_5495;
	wire _0960_;
	wire _0036_;
	wire _0456_;
	wire new_net_1370;
	wire new_net_1649;
	wire _0750_;
	wire new_net_222;
	wire new_net_2165;
	wire _0246_;
	wire new_net_3045;
	wire new_net_4354;
	wire new_net_6164;
	wire new_net_3616;
	wire new_net_1335;
	wire new_net_1437;
	wire new_net_1869;
	wire new_net_2774;
	wire new_net_3912;
	wire new_net_4307;
	wire new_net_4526;
	wire new_net_4614;
	wire new_net_4633;
	wire new_net_257;
	wire _0457_;
	wire _0751_;
	wire _0961_;
	wire new_net_1543;
	wire _0037_;
	wire new_net_1231;
	wire new_net_1720;
	wire new_net_2884;
	wire new_net_1507;
	wire new_net_7092;
	wire new_net_5416;
	wire new_net_7264;
	wire new_net_7481;
	wire new_net_189;
	wire new_net_432;
	wire new_net_903;
	wire new_net_1268;
	wire new_net_1472;
	wire new_net_3873;
	wire new_net_4207;
	wire new_net_5406;
	wire new_net_6447;
	wire new_net_7340;
	wire new_net_7653;
	wire new_net_7586;
	wire new_net_8232;
	wire new_net_3852;
	wire _0458_;
	wire _0752_;
	wire _0962_;
	wire new_net_1581;
	wire new_net_2260;
	wire new_net_3751;
	wire new_net_1371;
	wire new_net_1650;
	wire _0038_;
	wire new_net_2437;
	wire new_net_6808;
	wire new_net_7431;
	wire new_net_7603;
	wire new_net_293;
	wire new_net_329;
	wire new_net_1336;
	wire new_net_1438;
	wire new_net_3366;
	wire new_net_3750;
	wire new_net_3357;
	wire new_net_4308;
	wire new_net_4394;
	wire new_net_5651;
	wire new_net_6201;
	wire new_net_6736;
	wire new_net_6734;
	wire new_net_7024;
	wire new_net_4172;
	wire new_net_7196;
	wire _0249_;
	wire new_net_1508;
	wire _0963_;
	wire _0459_;
	wire _0753_;
	wire new_net_258;
	wire new_net_2047;
	wire _0039_;
	wire new_net_1232;
	wire new_net_2885;
	wire new_net_4594;
	wire new_net_5274;
	wire new_net_6138;
	wire new_net_5486;
	wire new_net_6968;
	wire new_net_4997;
	wire new_net_5731;
	wire new_net_6928;
	wire new_net_3046;
	wire new_net_190;
	wire new_net_433;
	wire new_net_904;
	wire new_net_1269;
	wire new_net_1473;
	wire new_net_4271;
	wire new_net_4295;
	wire new_net_4675;
	wire new_net_4847;
	wire new_net_6477;
	wire new_net_7925;
	wire _0250_;
	wire new_net_1303;
	wire _0964_;
	wire new_net_3617;
	wire new_net_1582;
	wire _0460_;
	wire new_net_1372;
	wire new_net_1651;
	wire new_net_1795;
	wire _0040_;
	wire new_net_6950;
	wire new_net_5012;
	wire new_net_5804;
	wire new_net_4340;
	wire new_net_1774;
	wire new_net_294;
	wire new_net_330;
	wire new_net_1544;
	wire new_net_1995;
	wire new_net_3259;
	wire new_net_1841;
	wire new_net_4656;
	wire new_net_5629;
	wire new_net_6098;
	wire new_net_6639;
	wire new_net_7550;
	wire new_net_8208;
	wire new_net_7472;
	wire new_net_5085;
	wire new_net_6315;
	wire _0251_;
	wire new_net_2916;
	wire _0461_;
	wire _0755_;
	wire _0965_;
	wire new_net_259;
	wire new_net_1791;
	wire _0041_;
	wire new_net_1233;
	wire new_net_3874;
	wire new_net_7400;
	wire new_net_7572;
	wire new_net_7073;
	wire new_net_4894;
	wire new_net_7777;
	wire new_net_1270;
	wire new_net_1474;
	wire new_net_2898;
	wire new_net_3;
	wire new_net_224;
	wire new_net_434;
	wire new_net_905;
	wire new_net_5145;
	wire new_net_6695;
	wire new_net_6798;
	wire new_net_7071;
	wire new_net_8196;
	wire new_net_5444;
	wire _0252_;
	wire _0462_;
	wire _0756_;
	wire new_net_1337;
	wire _0966_;
	wire new_net_2000;
	wire new_net_2261;
	wire new_net_3367;
	wire _0000_;
	wire new_net_1373;
	wire new_net_4458;
	wire new_net_6604;
	wire new_net_8135;
	wire new_net_5584;
	wire new_net_3596;
	wire new_net_3581;
	wire new_net_1509;
	wire new_net_1545;
	wire new_net_3931;
	wire new_net_3970;
	wire new_net_4171;
	wire new_net_4359;
	wire new_net_4548;
	wire new_net_5954;
	wire new_net_8267;
	wire new_net_6124;
	wire new_net_4520;
	wire new_net_5356;
	wire new_net_5354;
	wire new_net_191;
	wire new_net_1234;
	wire _0757_;
	wire _0001_;
	wire _0043_;
	wire _0253_;
	wire new_net_3047;
	wire _0967_;
	wire new_net_260;
	wire _0463_;
	wire new_net_4826;
	wire new_net_7916;
	wire new_net_1475;
	wire new_net_225;
	wire new_net_435;
	wire new_net_1304;
	wire new_net_3618;
	wire new_net_1583;
	wire new_net_3896;
	wire new_net_4635;
	wire new_net_4690;
	wire new_net_5110;
	wire new_net_5661;
	wire new_net_6369;
	wire new_net_3260;
	wire new_net_1440;
	wire _0758_;
	wire new_net_2167;
	wire _0002_;
	wire _0044_;
	wire _0254_;
	wire new_net_1338;
	wire _0968_;
	wire _1158_;
	wire new_net_4082;
	wire new_net_6391;
	wire new_net_7042;
	wire new_net_1510;
	wire new_net_1546;
	wire new_net_3597;
	wire new_net_3875;
	wire new_net_4987;
	wire new_net_5408;
	wire new_net_6449;
	wire new_net_7342;
	wire new_net_7773;
	wire new_net_8163;
	wire new_net_5989;
	wire new_net_7308;
	wire new_net_8216;
	wire new_net_906;
	wire new_net_192;
	wire new_net_1235;
	wire new_net_1271;
	wire new_net_1766;
	wire new_net_2469;
	wire new_net_2899;
	wire _0465_;
	wire _0759_;
	wire _0255_;
	wire new_net_5131;
	wire new_net_5749;
	wire new_net_7153;
	wire new_net_7937;
	wire new_net_8187;
	wire new_net_4952;
	wire new_net_6011;
	wire new_net_226;
	wire new_net_436;
	wire new_net_1305;
	wire new_net_1584;
	wire new_net_3368;
	wire new_net_1653;
	wire new_net_3404;
	wire new_net_3914;
	wire new_net_5653;
	wire new_net_6249;
	wire new_net_7175;
	wire new_net_1754;
	wire _0256_;
	wire _0046_;
	wire _0004_;
	wire _0760_;
	wire new_net_3582;
	wire new_net_1830;
	wire _0970_;
	wire new_net_2262;
	wire _0466_;
	wire new_net_1547;
	wire new_net_1843;
	wire new_net_3898;
	wire new_net_4273;
	wire new_net_4297;
	wire new_net_4849;
	wire new_net_5132;
	wire new_net_7320;
	wire new_net_8025;
	wire new_net_8141;
	wire new_net_5849;
	wire new_net_6795;
	wire new_net_6883;
	wire new_net_7829;
	wire new_net_7418;
	wire new_net_907;
	wire new_net_2359;
	wire new_net_1476;
	wire new_net_1236;
	wire new_net_2407;
	wire _0971_;
	wire _0257_;
	wire _0005_;
	wire _0047_;
	wire _0761_;
	wire new_net_6188;
	wire new_net_5625;
	wire new_net_4544;
	wire new_net_1654;
	wire new_net_3261;
	wire new_net_1441;
	wire new_net_227;
	wire new_net_437;
	wire new_net_1306;
	wire new_net_3405;
	wire new_net_3660;
	wire new_net_4226;
	wire new_net_4241;
	wire new_net_6616;
	wire new_net_6544;
	wire new_net_1376;
	wire _0006_;
	wire _0048_;
	wire _0258_;
	wire new_net_2168;
	wire _0762_;
	wire new_net_1511;
	wire new_net_3598;
	wire new_net_1829;
	wire _0972_;
	wire new_net_5607;
	wire new_net_7672;
	wire new_net_7299;
	wire new_net_5207;
	wire new_net_6395;
	wire new_net_7055;
	wire new_net_4759;
	wire new_net_6977;
	wire new_net_193;
	wire new_net_262;
	wire new_net_1548;
	wire new_net_2900;
	wire new_net_3352;
	wire new_net_4142;
	wire new_net_5379;
	wire new_net_5740;
	wire new_net_6566;
	wire new_net_6697;
	wire new_net_6937;
	wire new_net_4140;
	wire new_net_8178;
	wire new_net_6075;
	wire new_net_6653;
	wire _0469_;
	wire _0763_;
	wire _0259_;
	wire _0049_;
	wire _0007_;
	wire new_net_1237;
	wire new_net_1477;
	wire _0973_;
	wire new_net_1585;
	wire new_net_3369;
	wire new_net_7945;
	wire _1152_;
	wire new_net_6385;
	wire new_net_6307;
	wire new_net_333;
	wire new_net_438;
	wire new_net_1307;
	wire new_net_1340;
	wire new_net_1442;
	wire new_net_3583;
	wire new_net_3933;
	wire new_net_3972;
	wire new_net_4173;
	wire new_net_4361;
	wire new_net_7392;
	wire new_net_298;
	wire new_net_1377;
	wire new_net_1842;
	wire new_net_2435;
	wire _0470_;
	wire _0764_;
	wire _0260_;
	wire _0050_;
	wire _0008_;
	wire new_net_1512;
	wire new_net_6324;
	wire new_net_8016;
	wire new_net_4691;
	wire new_net_4618;
	wire new_net_7820;
	wire new_net_194;
	wire new_net_263;
	wire new_net_908;
	wire new_net_1273;
	wire new_net_1549;
	wire new_net_3620;
	wire new_net_3915;
	wire new_net_4637;
	wire new_net_5112;
	wire new_net_5527;
	wire new_net_6714;
	wire new_net_6346;
	wire new_net_5940;
	wire new_net_6596;
	wire new_net_8127;
	wire _0471_;
	wire new_net_1586;
	wire new_net_1655;
	wire new_net_1882;
	wire new_net_3262;
	wire new_net_3406;
	wire new_net_3661;
	wire _0261_;
	wire _0009_;
	wire _0051_;
	wire new_net_4356;
	wire new_net_8254;
	wire new_net_8055;
	wire new_net_8053;
	wire new_net_7614;
	wire new_net_7491;
	wire new_net_6457;
	wire new_net_1880;
	wire new_net_4;
	wire new_net_334;
	wire new_net_439;
	wire new_net_1308;
	wire new_net_3599;
	wire new_net_3877;
	wire new_net_5598;
	wire new_net_5654;
	wire new_net_6372;
	wire new_net_7596;
	wire new_net_2026;
	wire _0472_;
	wire new_net_299;
	wire new_net_1378;
	wire _0976_;
	wire _0010_;
	wire _0052_;
	wire _0262_;
	wire new_net_2901;
	wire new_net_2471;
	wire new_net_8247;
	wire new_net_7801;
	wire new_net_4459;
	wire new_net_6818;
	wire new_net_7852;
	wire new_net_3370;
	wire new_net_264;
	wire new_net_909;
	wire new_net_1274;
	wire new_net_1478;
	wire new_net_1550;
	wire new_net_1789;
	wire new_net_3955;
	wire new_net_4397;
	wire new_net_4616;
	wire new_net_6985;
	wire new_net_4708;
	wire new_net_7896;
	wire new_net_5302;
	wire new_net_7240;
	wire new_net_7034;
	wire new_net_4962;
	wire new_net_6293;
	wire new_net_3961;
	wire new_net_8159;
	wire new_net_1587;
	wire new_net_229;
	wire new_net_1656;
	wire _0977_;
	wire _0263_;
	wire _0011_;
	wire _0053_;
	wire new_net_3584;
	wire new_net_1239;
	wire new_net_1443;
	wire new_net_7378;
	wire new_net_5976;
	wire new_net_7958;
	wire new_net_3354;
	wire new_net_1925;
	wire new_net_440;
	wire new_net_1840;
	wire new_net_1309;
	wire new_net_1513;
	wire new_net_4275;
	wire new_net_4678;
	wire new_net_4851;
	wire new_net_5134;
	wire new_net_6025;
	wire new_net_6165;
	wire new_net_3621;
	wire _0978_;
	wire new_net_2264;
	wire new_net_300;
	wire _0474_;
	wire _0768_;
	wire _0054_;
	wire _0012_;
	wire new_net_1379;
	wire new_net_1822;
	wire new_net_5926;
	wire new_net_1551;
	wire new_net_265;
	wire new_net_910;
	wire new_net_1275;
	wire new_net_3263;
	wire new_net_3407;
	wire new_net_1479;
	wire new_net_4660;
	wire new_net_4692;
	wire new_net_5633;
	wire new_net_7093;
	wire new_net_7265;
	wire new_net_7482;
	wire _0979_;
	wire new_net_1588;
	wire _0475_;
	wire _0769_;
	wire _0055_;
	wire _0013_;
	wire new_net_335;
	wire new_net_1657;
	wire new_net_3662;
	wire new_net_1240;
	wire new_net_3535;
	wire new_net_7654;
	wire new_net_7587;
	wire new_net_8233;
	wire new_net_2917;
	wire new_net_3048;
	wire new_net_441;
	wire new_net_1310;
	wire new_net_1514;
	wire new_net_1935;
	wire new_net_2902;
	wire new_net_4312;
	wire new_net_5957;
	wire new_net_6699;
	wire new_net_6430;
	wire new_net_6809;
	wire new_net_7432;
	wire _0266_;
	wire new_net_3371;
	wire _0980_;
	wire _0014_;
	wire _0056_;
	wire _0476_;
	wire new_net_301;
	wire new_net_1380;
	wire new_net_196;
	wire _0770_;
	wire new_net_7604;
	wire new_net_6202;
	wire new_net_6737;
	wire new_net_6735;
	wire new_net_7025;
	wire new_net_6831;
	wire new_net_8150;
	wire new_net_4661;
	wire new_net_1933;
	wire new_net_1796;
	wire new_net_1552;
	wire new_net_3585;
	wire new_net_3935;
	wire new_net_3974;
	wire new_net_4175;
	wire new_net_4617;
	wire new_net_4970;
	wire new_net_5410;
	wire new_net_4865;
	wire new_net_6759;
	wire new_net_6757;
	wire new_net_5487;
	wire new_net_2918;
	wire new_net_3049;
	wire new_net_1343;
	wire new_net_1818;
	wire _0981_;
	wire _0267_;
	wire _0057_;
	wire _0015_;
	wire _0477_;
	wire new_net_336;
	wire new_net_4998;
	wire new_net_6929;
	wire new_net_7013;
	wire new_net_7926;
	wire new_net_5790;
	wire new_net_1311;
	wire new_net_1515;
	wire new_net_3622;
	wire new_net_1924;
	wire new_net_3258;
	wire new_net_4529;
	wire new_net_4549;
	wire new_net_4639;
	wire new_net_5114;
	wire new_net_5509;
	wire new_net_7451;
	wire new_net_6015;
	wire _0268_;
	wire new_net_2265;
	wire new_net_266;
	wire _0478_;
	wire _0772_;
	wire _0982_;
	wire _0016_;
	wire new_net_302;
	wire new_net_2538;
	wire new_net_3264;
	wire new_net_3899;
	wire new_net_7558;
	wire new_net_7551;
	wire new_net_8209;
	wire new_net_7473;
	wire new_net_4797;
	wire new_net_4538;
	wire new_net_3601;
	wire new_net_1553;
	wire new_net_1589;
	wire new_net_912;
	wire new_net_1241;
	wire new_net_1277;
	wire new_net_3879;
	wire new_net_3956;
	wire new_net_6374;
	wire new_net_6453;
	wire new_net_5827;
	wire new_net_6861;
	wire new_net_7401;
	wire new_net_7573;
	wire new_net_442;
	wire _0269_;
	wire new_net_1344;
	wire _0479_;
	wire _0773_;
	wire new_net_2903;
	wire _0983_;
	wire new_net_2473;
	wire _0017_;
	wire new_net_337;
	wire new_net_5224;
	wire new_net_7074;
	wire new_net_8197;
	wire new_net_1516;
	wire new_net_1828;
	wire new_net_1312;
	wire new_net_1381;
	wire new_net_3372;
	wire new_net_2534;
	wire new_net_6351;
	wire new_net_7919;
	wire new_net_8041;
	wire new_net_5614;
	wire new_net_6605;
	wire new_net_8136;
	wire new_net_5585;
	wire new_net_2055;
	wire new_net_1481;
	wire new_net_2171;
	wire new_net_3586;
	wire _0270_;
	wire _0984_;
	wire _0480_;
	wire _0774_;
	wire _0018_;
	wire new_net_267;
	wire new_net_5960;
	wire new_net_7279;
	wire new_net_8268;
	wire new_net_2919;
	wire new_net_232;
	wire new_net_913;
	wire new_net_1242;
	wire new_net_1278;
	wire new_net_1554;
	wire new_net_1590;
	wire new_net_4277;
	wire new_net_4853;
	wire new_net_5136;
	wire new_net_4827;
	wire new_net_7917;
	wire new_net_5859;
	wire new_net_5578;
	wire new_net_1447;
	wire new_net_2411;
	wire new_net_443;
	wire new_net_2777;
	wire _0271_;
	wire new_net_1752;
	wire new_net_3623;
	wire _0985_;
	wire _0481_;
	wire _0775_;
	wire new_net_6276;
	wire new_net_7644;
	wire new_net_7227;
	wire new_net_5866;
	wire new_net_6370;
	wire new_net_1517;
	wire new_net_198;
	wire new_net_1313;
	wire new_net_1382;
	wire new_net_3265;
	wire new_net_4662;
	wire new_net_4694;
	wire new_net_5635;
	wire new_net_7198;
	wire new_net_4527;
	wire new_net_7043;
	wire _0062_;
	wire new_net_1482;
	wire _0272_;
	wire new_net_3602;
	wire _0482_;
	wire _0776_;
	wire _0986_;
	wire new_net_2266;
	wire _0020_;
	wire new_net_304;
	wire new_net_4679;
	wire new_net_5990;
	wire new_net_7309;
	wire new_net_7911;
	wire new_net_8217;
	wire new_net_1279;
	wire new_net_2904;
	wire new_net_233;
	wire new_net_914;
	wire new_net_1345;
	wire new_net_1555;
	wire new_net_2964;
	wire new_net_3663;
	wire new_net_4363;
	wire new_net_4968;
	wire new_net_7938;
	wire new_net_8188;
	wire new_net_7326;
	wire new_net_6012;
	wire new_net_6668;
	wire _0063_;
	wire _0273_;
	wire new_net_3050;
	wire _0483_;
	wire _0777_;
	wire _0987_;
	wire new_net_3373;
	wire _0021_;
	wire new_net_339;
	wire new_net_1661;
	wire new_net_5409;
	wire new_net_5326;
	wire new_net_1773;
	wire new_net_3587;
	wire new_net_1518;
	wire new_net_199;
	wire new_net_268;
	wire new_net_1314;
	wire new_net_1792;
	wire new_net_1934;
	wire new_net_3937;
	wire new_net_3976;
	wire new_net_4054;
	wire new_net_8026;
	wire new_net_6884;
	wire new_net_6796;
	wire new_net_7830;
	wire new_net_7713;
	wire new_net_6189;
	wire new_net_7513;
	wire new_net_2130;
	wire _0526_;
	wire _1030_;
	wire _1240_;
	wire new_net_3719;
	wire new_net_2193;
	wire new_net_1609;
	wire new_net_4063;
	wire new_net_4743;
	wire new_net_5149;
	wire new_net_6356;
	wire new_net_7363;
	wire new_net_357;
	wire new_net_2541;
	wire new_net_4322;
	wire new_net_4864;
	wire new_net_5006;
	wire new_net_6509;
	wire new_net_6758;
	wire new_net_8077;
	wire new_net_8180;
	wire new_net_8204;
	wire _0150_;
	wire new_net_6545;
	wire new_net_5648;
	wire new_net_5608;
	wire new_net_1987;
	wire new_net_3454;
	wire _0527_;
	wire _1031_;
	wire _1241_;
	wire new_net_76;
	wire new_net_3383;
	wire new_net_4450;
	wire new_net_4707;
	wire new_net_4974;
	wire new_net_7673;
	wire new_net_7798;
	wire new_net_7300;
	wire new_net_6143;
	wire new_net_5208;
	wire new_net_7056;
	wire new_net_6978;
	wire new_net_5380;
	wire new_net_6567;
	wire new_net_6938;
	wire new_net_3909;
	wire new_net_1893;
	wire new_net_2974;
	wire new_net_1681;
	wire new_net_4011;
	wire new_net_5275;
	wire new_net_5548;
	wire new_net_7106;
	wire new_net_7209;
	wire new_net_7360;
	wire new_net_7688;
	wire new_net_8179;
	wire new_net_6654;
	wire new_net_1610;
	wire new_net_3417;
	wire new_net_2763;
	wire _1032_;
	wire _0528_;
	wire _1242_;
	wire new_net_2511;
	wire new_net_2225;
	wire new_net_3057;
	wire new_net_5424;
	wire new_net_7946;
	wire new_net_7167;
	wire new_net_6386;
	wire new_net_358;
	wire new_net_3791;
	wire new_net_4344;
	wire new_net_4409;
	wire new_net_4431;
	wire new_net_4469;
	wire new_net_4493;
	wire new_net_5027;
	wire new_net_5745;
	wire new_net_5819;
	wire new_net_7393;
	wire new_net_5780;
	wire new_net_4977;
	wire new_net_6408;
	wire new_net_8017;
	wire new_net_6325;
	wire new_net_77;
	wire new_net_3646;
	wire new_net_2994;
	wire new_net_3681;
	wire _1033_;
	wire _0529_;
	wire _1243_;
	wire new_net_3884;
	wire new_net_3916;
	wire new_net_3989;
	wire new_net_4258;
	wire new_net_8255;
	wire new_net_7990;
	wire new_net_4000;
	wire new_net_6180;
	wire new_net_1682;
	wire new_net_3720;
	wire new_net_4064;
	wire new_net_4744;
	wire new_net_5150;
	wire new_net_5526;
	wire new_net_5528;
	wire new_net_5892;
	wire new_net_6117;
	wire new_net_6347;
	wire new_net_6715;
	wire new_net_5039;
	wire new_net_6597;
	wire new_net_8128;
	wire new_net_4282;
	wire new_net_6108;
	wire new_net_7349;
	wire new_net_1611;
	wire new_net_2058;
	wire new_net_2365;
	wire new_net_3418;
	wire new_net_2131;
	wire new_net_2625;
	wire _0530_;
	wire _1034_;
	wire _1244_;
	wire new_net_2194;
	wire new_net_8056;
	wire new_net_6909;
	wire new_net_4300;
	wire new_net_6458;
	wire new_net_4555;
	wire new_net_359;
	wire new_net_4208;
	wire new_net_4342;
	wire new_net_5072;
	wire new_net_5996;
	wire new_net_7442;
	wire new_net_7545;
	wire new_net_8078;
	wire new_net_5194;
	wire new_net_6969;
	wire new_net_8248;
	wire _1035_;
	wire new_net_78;
	wire new_net_2975;
	wire _0531_;
	wire _1245_;
	wire new_net_2540;
	wire new_net_4012;
	wire new_net_4315;
	wire new_net_5276;
	wire new_net_5549;
	wire new_net_7804;
	wire new_net_6067;
	wire new_net_6819;
	wire new_net_7853;
	wire new_net_7732;
	wire new_net_7730;
	wire new_net_2082;
	wire new_net_2006;
	wire new_net_2764;
	wire new_net_5425;
	wire new_net_5791;
	wire new_net_5973;
	wire new_net_6533;
	wire new_net_7062;
	wire new_net_7419;
	wire new_net_7955;
	wire new_net_7897;
	wire new_net_5676;
	wire new_net_7035;
	wire new_net_4961;
	wire new_net_6294;
	wire new_net_8160;
	wire new_net_5805;
	wire new_net_2226;
	wire new_net_2946;
	wire new_net_1612;
	wire _1036_;
	wire _0532_;
	wire _1246_;
	wire new_net_3792;
	wire new_net_4410;
	wire new_net_4432;
	wire new_net_4470;
	wire new_net_7379;
	wire new_net_7959;
	wire new_net_6316;
	wire new_net_2995;
	wire new_net_360;
	wire new_net_1978;
	wire new_net_3434;
	wire new_net_3682;
	wire new_net_2786;
	wire new_net_3870;
	wire new_net_3990;
	wire new_net_4191;
	wire new_net_4323;
	wire new_net_7976;
	wire new_net_6166;
	wire new_net_2447;
	wire new_net_79;
	wire new_net_1902;
	wire new_net_3384;
	wire _1037_;
	wire _0533_;
	wire new_net_1683;
	wire new_net_2535;
	wire _1247_;
	wire new_net_2787;
	wire new_net_3721;
	wire new_net_4002;
	wire new_net_3059;
	wire new_net_2626;
	wire new_net_4866;
	wire new_net_6511;
	wire new_net_6760;
	wire new_net_8182;
	wire new_net_8206;
	wire new_net_4917;
	wire new_net_4246;
	wire new_net_5418;
	wire new_net_7266;
	wire new_net_7107;
	wire new_net_7483;
	wire new_net_2195;
	wire new_net_2947;
	wire _0534_;
	wire _1038_;
	wire new_net_2433;
	wire new_net_2132;
	wire new_net_4343;
	wire new_net_5073;
	wire new_net_5997;
	wire new_net_7443;
	wire new_net_7588;
	wire new_net_8234;
	wire new_net_3854;
	wire new_net_2976;
	wire new_net_361;
	wire new_net_4721;
	wire new_net_5277;
	wire new_net_5550;
	wire new_net_7108;
	wire new_net_7211;
	wire new_net_6431;
	wire new_net_7362;
	wire new_net_7690;
	wire new_net_6810;
	wire new_net_7433;
	wire new_net_7605;
	wire _0535_;
	wire _1039_;
	wire new_net_1684;
	wire new_net_4762;
	wire new_net_5426;
	wire new_net_5670;
	wire new_net_5792;
	wire new_net_5974;
	wire new_net_6203;
	wire new_net_6534;
	wire new_net_6738;
	wire new_net_7026;
	wire new_net_4174;
	wire new_net_6832;
	wire new_net_8151;
	wire new_net_21;
	wire new_net_1613;
	wire new_net_2083;
	wire new_net_3793;
	wire new_net_4433;
	wire new_net_4471;
	wire new_net_4495;
	wire new_net_5029;
	wire new_net_5747;
	wire new_net_6489;
	wire new_net_431;
	wire new_net_6392;
	wire new_net_5488;
	wire new_net_3683;
	wire new_net_2227;
	wire _1040_;
	wire _0536_;
	wire new_net_2996;
	wire new_net_3455;
	wire new_net_3991;
	wire new_net_4192;
	wire new_net_5008;
	wire new_net_5769;
	wire new_net_7014;
	wire new_net_7927;
	wire new_net_2661;
	wire new_net_3722;
	wire new_net_2836;
	wire new_net_3647;
	wire new_net_80;
	wire new_net_3538;
	wire new_net_4066;
	wire new_net_4452;
	wire new_net_4722;
	wire new_net_4746;
	wire new_net_5918;
	wire new_net_6952;
	wire new_net_7454;
	wire new_net_7452;
	wire new_net_1857;
	wire new_net_3060;
	wire new_net_3435;
	wire _1041_;
	wire _0537_;
	wire new_net_2367;
	wire new_net_2627;
	wire new_net_4324;
	wire new_net_4867;
	wire new_net_6512;
	wire new_net_6634;
	wire new_net_7559;
	wire new_net_7552;
	wire new_net_8210;
	wire new_net_4605;
	wire new_net_7474;
	wire new_net_2183;
	wire new_net_8004;
	wire new_net_2948;
	wire new_net_1614;
	wire new_net_4347;
	wire new_net_5074;
	wire new_net_5998;
	wire new_net_3363;
	wire new_net_7444;
	wire new_net_7547;
	wire new_net_5828;
	wire new_net_261;
	wire new_net_7574;
	wire new_net_7075;
	wire new_net_2133;
	wire new_net_2196;
	wire new_net_2539;
	wire new_net_2788;
	wire _0538_;
	wire _1042_;
	wire new_net_2977;
	wire new_net_362;
	wire new_net_4411;
	wire new_net_5278;
	wire new_net_8198;
	wire new_net_81;
	wire new_net_3648;
	wire new_net_3539;
	wire new_net_1685;
	wire new_net_3419;
	wire new_net_5427;
	wire new_net_5671;
	wire new_net_5793;
	wire new_net_5975;
	wire new_net_6535;
	wire new_net_6606;
	wire new_net_5586;
	wire _0539_;
	wire _1043_;
	wire new_net_3794;
	wire new_net_4434;
	wire new_net_4472;
	wire new_net_4496;
	wire new_net_4695;
	wire new_net_4709;
	wire new_net_5030;
	wire new_net_5748;
	wire new_net_8269;
	wire new_net_4693;
	wire new_net_6126;
	wire new_net_5358;
	wire new_net_2630;
	wire new_net_3684;
	wire new_net_1615;
	wire new_net_2997;
	wire new_net_3992;
	wire new_net_4193;
	wire new_net_5009;
	wire new_net_5770;
	wire new_net_5873;
	wire new_net_6615;
	wire new_net_4828;
	wire new_net_7918;
	wire new_net_363;
	wire new_net_3723;
	wire new_net_2228;
	wire _1044_;
	wire _0540_;
	wire new_net_4067;
	wire new_net_4723;
	wire new_net_4747;
	wire new_net_5153;
	wire new_net_5529;
	wire new_net_5663;
	wire new_net_4253;
	wire new_net_6371;
	wire new_net_5882;
	wire new_net_1686;
	wire new_net_3420;
	wire new_net_3436;
	wire new_net_3061;
	wire new_net_4325;
	wire new_net_4868;
	wire new_net_6513;
	wire new_net_6762;
	wire new_net_8184;
	wire new_net_4084;
	wire new_net_7044;
	wire new_net_2169;
	wire new_net_2949;
	wire _1045_;
	wire _0541_;
	wire new_net_2628;
	wire new_net_4345;
	wire new_net_4453;
	wire new_net_5075;
	wire new_net_5999;
	wire new_net_7445;
	wire new_net_7548;
	wire new_net_5991;
	wire new_net_7310;
	wire new_net_8218;
	wire new_net_1616;
	wire new_net_2978;
	wire new_net_5279;
	wire new_net_5552;
	wire new_net_6490;
	wire new_net_6739;
	wire new_net_7110;
	wire new_net_5133;
	wire new_net_7213;
	wire new_net_7364;
	wire new_net_7155;
	wire new_net_4528;
	wire new_net_8189;
	wire new_net_7327;
	wire new_net_6013;
	wire new_net_2134;
	wire new_net_2197;
	wire _1046_;
	wire new_net_82;
	wire new_net_3649;
	wire _0542_;
	wire new_net_3540;
	wire new_net_5428;
	wire new_net_5672;
	wire new_net_5794;
	wire new_net_5117;
	wire new_net_7177;
	wire new_net_1687;
	wire new_net_2766;
	wire new_net_3795;
	wire new_net_3147;
	wire new_net_4412;
	wire new_net_4435;
	wire new_net_4473;
	wire new_net_4497;
	wire new_net_4710;
	wire new_net_5031;
	wire new_net_2998;
	wire new_net_3685;
	wire _0543_;
	wire _1047_;
	wire new_net_2076;
	wire new_net_3993;
	wire new_net_4194;
	wire new_net_5010;
	wire new_net_5771;
	wire new_net_5874;
	wire new_net_3894;
	wire new_net_6885;
	wire new_net_7420;
	wire new_net_4218;
	wire _0464_;
	wire new_net_295;
	wire new_net_3009;
	wire new_net_3724;
	wire new_net_364;
	wire new_net_1617;
	wire new_net_4068;
	wire new_net_4724;
	wire new_net_4748;
	wire new_net_5154;
	wire new_net_5530;
	wire new_net_5896;
	wire new_net_6190;
	wire new_net_7514;
	wire new_net_2483;
	wire new_net_6357;
	wire new_net_3950;
	wire new_net_4391;
	wire new_net_1148;
	wire new_net_3948;
	wire new_net_4545;
	wire new_net_2369;
	wire new_net_1979;
	wire _0544_;
	wire new_net_2229;
	wire new_net_3062;
	wire _1048_;
	wire new_net_83;
	wire new_net_2837;
	wire new_net_4029;
	wire new_net_4326;
	wire new_net_6618;
	wire new_net_5020;
	wire _0432_;
	wire new_net_6546;
	wire new_net_5649;
	wire new_net_2629;
	wire new_net_2542;
	wire new_net_2950;
	wire new_net_4346;
	wire new_net_4454;
	wire new_net_5076;
	wire new_net_5609;
	wire new_net_6000;
	wire new_net_7446;
	wire new_net_7549;
	wire new_net_7674;
	wire new_net_6144;
	wire new_net_5209;
	wire new_net_7057;
	wire new_net_2979;
	wire new_net_3456;
	wire _1049_;
	wire _0545_;
	wire new_net_4013;
	wire new_net_4761;
	wire new_net_5280;
	wire new_net_4144;
	wire new_net_5381;
	wire new_net_5553;
	wire new_net_5742;
	wire new_net_6568;
	wire new_net_6939;
	wire new_net_7645;
	wire new_net_6655;
	wire new_net_1444;
	wire new_net_3338;
	wire new_net_1618;
	wire new_net_3650;
	wire new_net_3541;
	wire new_net_3010;
	wire new_net_365;
	wire new_net_5429;
	wire new_net_5673;
	wire new_net_5977;
	wire new_net_6537;
	wire new_net_6640;
	wire new_net_7947;
	wire new_net_7168;
	wire new_net_5318;
	wire new_net_3526;
	wire new_net_6387;
	wire new_net_1688;
	wire new_net_2135;
	wire new_net_2767;
	wire new_net_2198;
	wire _1050_;
	wire _0546_;
	wire new_net_3796;
	wire new_net_4413;
	wire new_net_4474;
	wire new_net_4498;
	wire new_net_7394;
	wire new_net_4026;
	wire new_net_6411;
	wire new_net_3686;
	wire new_net_2999;
	wire new_net_3994;
	wire new_net_4195;
	wire new_net_5011;
	wire new_net_5772;
	wire new_net_5875;
	wire new_net_6409;
	wire new_net_6617;
	wire new_net_7237;
	wire new_net_6326;
	wire new_net_8018;
	wire _1051_;
	wire _0547_;
	wire new_net_2662;
	wire new_net_3725;
	wire new_net_4069;
	wire new_net_4209;
	wire new_net_4725;
	wire new_net_4749;
	wire new_net_5155;
	wire new_net_5531;
	wire new_net_6348;
	wire new_net_641;
	wire new_net_5040;
	wire new_net_6598;
	wire new_net_2423;
	wire new_net_8129;
	wire new_net_6109;
	wire new_net_7350;
	wire new_net_3063;
	wire new_net_84;
	wire new_net_1619;
	wire new_net_2789;
	wire new_net_4210;
	wire new_net_4327;
	wire new_net_4870;
	wire new_net_6764;
	wire new_net_7365;
	wire new_net_8186;
	wire new_net_6488;
	wire new_net_5551;
	wire new_net_8057;
	wire new_net_5173;
	wire new_net_7616;
	wire new_net_6910;
	wire new_net_7493;
	wire new_net_2951;
	wire _1052_;
	wire new_net_1689;
	wire _0548_;
	wire new_net_2543;
	wire new_net_2230;
	wire new_net_5077;
	wire new_net_5600;
	wire new_net_5795;
	wire new_net_6001;
	wire new_net_6459;
	wire new_net_8079;
	wire new_net_711;
	wire new_net_2980;
	wire new_net_5281;
	wire new_net_5554;
	wire new_net_5750;
	wire new_net_6492;
	wire new_net_6741;
	wire new_net_6970;
	wire new_net_7112;
	wire new_net_7215;
	wire new_net_7694;
	wire new_net_1971;
	wire new_net_7733;
	wire new_net_2077;
	wire new_net_3651;
	wire new_net_3542;
	wire new_net_366;
	wire new_net_2431;
	wire new_net_3421;
	wire _1053_;
	wire _0549_;
	wire new_net_2663;
	wire new_net_4042;
	wire new_net_6987;
	wire new_net_7900;
	wire new_net_7898;
	wire new_net_7036;
	wire new_net_4184;
	wire new_net_6958;
	wire new_net_6295;
	wire new_net_3425;
	wire new_net_2768;
	wire new_net_3437;
	wire new_net_85;
	wire new_net_3457;
	wire new_net_3797;
	wire new_net_4475;
	wire new_net_4499;
	wire new_net_5033;
	wire new_net_5806;
	wire new_net_8161;
	wire new_net_7380;
	wire new_net_5978;
	wire new_net_6641;
	wire new_net_7960;
	wire new_net_1705;
	wire new_net_1690;
	wire new_net_3000;
	wire new_net_2136;
	wire new_net_3687;
	wire _1054_;
	wire _0550_;
	wire new_net_2199;
	wire new_net_3995;
	wire new_net_4015;
	wire new_net_4196;
	wire new_net_6317;
	wire new_net_7527;
	wire new_net_3726;
	wire new_net_4030;
	wire new_net_4070;
	wire new_net_4302;
	wire new_net_4455;
	wire new_net_4726;
	wire new_net_4750;
	wire new_net_5156;
	wire new_net_5532;
	wire new_net_5898;
	wire new_net_5928;
	wire new_net_3777;
	wire new_net_3422;
	wire new_net_3064;
	wire new_net_1912;
	wire new_net_367;
	wire new_net_2371;
	wire _0551_;
	wire _1055_;
	wire new_net_3104;
	wire new_net_4328;
	wire new_net_4990;
	wire new_net_5419;
	wire new_net_7484;
	wire new_net_2544;
	wire new_net_2952;
	wire new_net_1723;
	wire new_net_86;
	wire new_net_945;
	wire new_net_2631;
	wire new_net_3438;
	wire new_net_4014;
	wire new_net_3537;
	wire new_net_5078;
	wire new_net_7280;
	wire new_net_2281;
	wire new_net_4959;
	wire new_net_3130;
	wire new_net_2231;
	wire new_net_2838;
	wire new_net_2981;
	wire new_net_1691;
	wire _0552_;
	wire _1056_;
	wire new_net_5282;
	wire new_net_5555;
	wire new_net_5751;
	wire new_net_6493;
	wire new_net_7589;
	wire new_net_8235;
	wire new_net_6811;
	wire new_net_7434;
	wire new_net_2312;
	wire new_net_2664;
	wire new_net_3543;
	wire new_net_1858;
	wire new_net_5431;
	wire new_net_5458;
	wire new_net_5675;
	wire new_net_5773;
	wire new_net_5979;
	wire new_net_6515;
	wire new_net_6642;
	wire new_net_7606;
	wire new_net_7228;
	wire new_net_1621;
	wire _1057_;
	wire _0553_;
	wire new_net_3798;
	wire new_net_4476;
	wire new_net_4500;
	wire new_net_5034;
	wire new_net_6123;
	wire new_net_6719;
	wire new_net_6049;
	wire new_net_6833;
	wire new_net_8152;
	wire new_net_6761;
	wire new_net_296;
	wire new_net_6393;
	wire new_net_87;
	wire new_net_2769;
	wire new_net_3688;
	wire new_net_3996;
	wire new_net_4197;
	wire new_net_5013;
	wire new_net_5368;
	wire new_net_5489;
	wire new_net_5877;
	wire new_net_6555;
	wire new_net_5000;
	wire new_net_4680;
	wire new_net_8064;
	wire new_net_7015;
	wire new_net_7928;
	wire new_net_1149;
	wire new_net_2200;
	wire new_net_3727;
	wire new_net_2839;
	wire new_net_1692;
	wire _1058_;
	wire _0554_;
	wire new_net_331;
	wire new_net_812;
	wire new_net_1988;
	wire new_net_2137;
	wire new_net_4546;
	wire new_net_6037;
	wire new_net_5511;
	wire new_net_6577;
	wire new_net_7939;
	wire new_net_3918;
	wire new_net_4260;
	wire new_net_4777;
	wire new_net_3965;
	wire new_net_3423;
	wire new_net_2790;
	wire new_net_3065;
	wire new_net_368;
	wire new_net_1980;
	wire new_net_3963;
	wire new_net_4872;
	wire new_net_6766;
	wire new_net_7367;
	wire new_net_7597;
	wire new_net_7560;
	wire new_net_7553;
	wire new_net_8211;
	wire new_net_7475;
	wire new_net_2632;
	wire new_net_3439;
	wire new_net_2545;
	wire new_net_2953;
	wire _0555_;
	wire _1059_;
	wire new_net_4414;
	wire new_net_4456;
	wire new_net_4540;
	wire new_net_4712;
	wire new_net_4799;
	wire new_net_8005;
	wire new_net_3364;
	wire new_net_8099;
	wire new_net_4731;
	wire new_net_1445;
	wire new_net_7575;
	wire new_net_2982;
	wire new_net_88;
	wire new_net_2536;
	wire new_net_3778;
	wire new_net_4113;
	wire new_net_5283;
	wire new_net_5556;
	wire new_net_5752;
	wire new_net_6494;
	wire new_net_7076;
	wire new_net_7782;
	wire new_net_1942;
	wire new_net_5226;
	wire new_net_5148;
	wire new_net_8199;
	wire new_net_2665;
	wire new_net_2791;
	wire new_net_2232;
	wire new_net_3385;
	wire new_net_3544;
	wire _0556_;
	wire _1060_;
	wire new_net_1693;
	wire new_net_5432;
	wire new_net_5449;
	wire new_net_5616;
	wire new_net_1292;
	wire new_net_8138;
	wire new_net_1622;
	wire new_net_369;
	wire new_net_3799;
	wire new_net_4415;
	wire new_net_4436;
	wire new_net_4477;
	wire new_net_4501;
	wire new_net_5035;
	wire new_net_5587;
	wire new_net_6720;
	wire new_net_4228;
	wire new_net_5962;
	wire new_net_2770;
	wire new_net_3689;
	wire new_net_1914;
	wire _0557_;
	wire _1061_;
	wire new_net_3997;
	wire new_net_4198;
	wire new_net_4329;
	wire new_net_5014;
	wire new_net_5359;
	wire new_net_5861;
	wire new_net_3728;
	wire new_net_2840;
	wire new_net_3386;
	wire new_net_89;
	wire new_net_4032;
	wire new_net_2184;
	wire new_net_4072;
	wire new_net_4728;
	wire new_net_4752;
	wire new_net_5158;
	wire new_net_5580;
	wire new_net_6278;
	wire new_net_5470;
	wire _0124_;
	wire new_net_1694;
	wire new_net_3424;
	wire new_net_2138;
	wire new_net_2201;
	wire new_net_2373;
	wire new_net_3066;
	wire _1062_;
	wire _0558_;
	wire new_net_6743;
	wire new_net_6767;
	wire new_net_4085;
	wire new_net_6679;
	wire _0467_;
	wire new_net_7045;
	wire new_net_3440;
	wire new_net_2954;
	wire new_net_1623;
	wire new_net_712;
	wire new_net_4457;
	wire new_net_5080;
	wire new_net_5980;
	wire new_net_6004;
	wire new_net_6643;
	wire new_net_7450;
	wire new_net_5079;
	wire new_net_5992;
	wire new_net_3656;
	wire new_net_6244;
	wire new_net_7311;
	wire new_net_8219;
	wire new_net_2983;
	wire new_net_3001;
	wire new_net_3458;
	wire _0559_;
	wire _1063_;
	wire new_net_456;
	wire new_net_3832;
	wire new_net_5284;
	wire new_net_5557;
	wire new_net_5753;
	wire new_net_5391;
	wire new_net_8190;
	wire new_net_7328;
	wire new_net_6014;
	wire new_net_2792;
	wire new_net_90;
	wire new_net_5677;
	wire new_net_5775;
	wire new_net_6517;
	wire new_net_7070;
	wire new_net_7963;
	wire new_net_6716;
	wire _1201_;
	wire new_net_5411;
	wire new_net_7178;
	wire new_net_370;
	wire new_net_1695;
	wire new_net_2233;
	wire _0560_;
	wire _1064_;
	wire new_net_3800;
	wire new_net_4416;
	wire new_net_4478;
	wire new_net_5036;
	wire new_net_1742;
	wire new_net_8256;
	wire new_net_3690;
	wire new_net_3459;
	wire new_net_3998;
	wire new_net_4199;
	wire new_net_4873;
	wire new_net_5015;
	wire new_net_5879;
	wire new_net_6621;
	wire new_net_7117;
	wire new_net_3571;
	wire new_net_6999;
	wire new_net_1404;
	wire new_net_1259;
	wire new_net_3058;
	wire new_net_6510;
	wire new_net_7421;
	wire new_net_7832;
	wire new_net_7711;
	wire new_net_2429;
	wire new_net_3013;
	wire new_net_3729;
	wire _0561_;
	wire _1065_;
	wire new_net_3387;
	wire new_net_4033;
	wire new_net_4073;
	wire new_net_4437;
	wire new_net_2170;
	wire new_net_7515;
	wire new_net_7805;
	wire new_net_6358;
	wire new_net_6532;
	wire new_net_3011;
	wire new_net_3067;
	wire new_net_91;
	wire new_net_4330;
	wire new_net_5628;
	wire new_net_6744;
	wire new_net_6768;
	wire new_net_946;
	wire new_net_7369;
	wire new_net_7599;
	wire _0264_;
	wire new_net_6619;
	wire new_net_606;
	wire new_net_8067;
	wire new_net_1624;
	wire new_net_371;
	wire new_net_1696;
	wire new_net_2139;
	wire new_net_3441;
	wire new_net_2202;
	wire new_net_2955;
	wire _1066_;
	wire _0562_;
	wire new_net_5065;
	wire new_net_5650;
	wire new_net_5891;
	wire new_net_6547;
	wire new_net_5610;
	wire new_net_4876;
	wire new_net_8089;
	wire new_net_4607;
	wire new_net_6145;
	wire new_net_2984;
	wire new_net_3780;
	wire new_net_5285;
	wire new_net_5210;
	wire new_net_5558;
	wire new_net_6125;
	wire new_net_6496;
	wire new_net_7058;
	wire new_net_7116;
	wire new_net_7219;
	wire _0084_;
	wire new_net_5087;
	wire new_net_5382;
	wire new_net_6569;
	wire new_net_6940;
	wire new_net_3911;
	wire new_net_1019;
	wire new_net_2761;
	wire new_net_2263;
	wire new_net_6656;
	wire _0563_;
	wire new_net_1981;
	wire new_net_3012;
	wire new_net_2793;
	wire _1067_;
	wire new_net_4016;
	wire new_net_4348;
	wire new_net_5678;
	wire new_net_471;
	wire new_net_5776;
	wire new_net_7948;
	wire new_net_7169;
	wire new_net_1722;
	wire _0468_;
	wire new_net_92;
	wire new_net_297;
	wire new_net_3801;
	wire new_net_4074;
	wire new_net_4349;
	wire new_net_4417;
	wire new_net_4479;
	wire new_net_5037;
	wire new_net_7097;
	wire new_net_5782;
	wire new_net_22;
	wire new_net_1625;
	wire new_net_1697;
	wire new_net_3691;
	wire new_net_3460;
	wire new_net_2234;
	wire _0564_;
	wire _1068_;
	wire new_net_3999;
	wire new_net_4200;
	wire new_net_6702;
	wire new_net_332;
	wire new_net_6410;
	wire new_net_8019;
	wire new_net_6327;
	wire new_net_7992;
	wire _0436_;
	wire new_net_3388;
	wire new_net_2666;
	wire new_net_3730;
	wire new_net_4034;
	wire new_net_4438;
	wire new_net_4714;
	wire new_net_4730;
	wire new_net_4754;
	wire new_net_5160;
	wire new_net_5799;
	wire new_net_6182;
	wire new_net_6349;
	wire _1202_;
	wire new_net_5041;
	wire new_net_6599;
	wire new_net_8130;
	wire _1069_;
	wire new_net_2375;
	wire new_net_2546;
	wire _0565_;
	wire new_net_3068;
	wire new_net_4284;
	wire new_net_4331;
	wire new_net_4350;
	wire new_net_4515;
	wire new_net_5754;
	wire new_net_6110;
	wire new_net_7351;
	wire new_net_5949;
	wire new_net_3679;
	wire new_net_4065;
	wire new_net_8058;
	wire new_net_6626;
	wire new_net_8270;
	wire new_net_7617;
	wire new_net_2956;
	wire new_net_3652;
	wire new_net_3442;
	wire new_net_93;
	wire new_net_372;
	wire new_net_1446;
	wire new_net_4502;
	wire new_net_5082;
	wire new_net_5434;
	wire new_net_5982;
	wire _0713_;
	wire new_net_6460;
	wire new_net_8080;
	wire new_net_2985;
	wire new_net_1698;
	wire new_net_3002;
	wire new_net_2140;
	wire new_net_1859;
	wire new_net_2203;
	wire new_net_2667;
	wire _1070_;
	wire _0566_;
	wire new_net_5559;
	wire new_net_6971;
	wire new_net_7879;
	wire new_net_4317;
	wire new_net_1293;
	wire new_net_5870;
	wire new_net_2547;
	wire new_net_2794;
	wire new_net_4017;
	wire new_net_5679;
	wire new_net_5777;
	wire new_net_6519;
	wire new_net_6821;
	wire new_net_7072;
	wire new_net_7734;
	wire new_net_7855;
	wire new_net_6988;
	wire _0265_;
	wire new_net_6209;
	wire new_net_7899;
	wire new_net_1725;
	wire _1071_;
	wire _0567_;
	wire new_net_3802;
	wire new_net_4418;
	wire new_net_4480;
	wire new_net_4503;
	wire new_net_6723;
	wire new_net_7037;
	wire new_net_7094;
	wire new_net_8162;
	wire new_net_5807;
	wire _0608_;
	wire new_net_7381;
	wire new_net_4986;
	wire new_net_7961;
	wire new_net_2389;
	wire new_net_3461;
	wire new_net_1626;
	wire new_net_2771;
	wire new_net_3692;
	wire new_net_94;
	wire new_net_373;
	wire new_net_4201;
	wire new_net_4875;
	wire new_net_5881;
	wire new_net_6623;
	wire new_net_5499;
	wire new_net_3872;
	wire new_net_6782;
	wire new_net_6236;
	wire new_net_7978;
	wire new_net_6168;
	wire new_net_4482;
	wire new_net_8027;
	wire new_net_4004;
	wire new_net_3928;
	wire _0106_;
	wire _0316_;
	wire _0820_;
	wire new_net_2932;
	wire new_net_3077;
	wire new_net_2298;
	wire new_net_3101;
	wire new_net_9;
	wire new_net_1168;
	wire _0610_;
	wire new_net_4719;
	wire new_net_5420;
	wire new_net_7109;
	wire new_net_7485;
	wire new_net_597;
	wire new_net_705;
	wire new_net_1026;
	wire new_net_2827;
	wire new_net_3636;
	wire new_net_2714;
	wire new_net_3835;
	wire new_net_5571;
	wire new_net_4150;
	wire new_net_5937;
	wire new_net_7281;
	wire new_net_7590;
	wire new_net_8236;
	wire _0611_;
	wire _0107_;
	wire _0317_;
	wire _0821_;
	wire new_net_3493;
	wire new_net_3132;
	wire new_net_3856;
	wire new_net_5320;
	wire new_net_6984;
	wire new_net_7709;
	wire new_net_3901;
	wire new_net_6812;
	wire new_net_7435;
	wire new_net_5459;
	wire new_net_563;
	wire new_net_1916;
	wire new_net_635;
	wire new_net_2680;
	wire new_net_2577;
	wire new_net_2061;
	wire new_net_4106;
	wire new_net_4786;
	wire new_net_5297;
	wire new_net_5445;
	wire new_net_6205;
	wire new_net_4176;
	wire new_net_8153;
	wire _0108_;
	wire _0318_;
	wire new_net_2475;
	wire _0822_;
	wire new_net_3184;
	wire new_net_495;
	wire new_net_2267;
	wire new_net_2330;
	wire _0612_;
	wire new_net_4911;
	wire new_net_6394;
	wire new_net_5490;
	wire new_net_5369;
	wire new_net_598;
	wire new_net_706;
	wire new_net_1027;
	wire new_net_2808;
	wire new_net_5094;
	wire new_net_5812;
	wire new_net_6556;
	wire new_net_6657;
	wire new_net_7756;
	wire new_net_7929;
	wire new_net_4547;
	wire _0109_;
	wire _0319_;
	wire _0823_;
	wire _0613_;
	wire new_net_2060;
	wire new_net_3553;
	wire new_net_3153;
	wire new_net_4888;
	wire new_net_5049;
	wire new_net_5712;
	wire new_net_6578;
	wire new_net_5920;
	wire new_net_5016;
	wire new_net_1169;
	wire new_net_2933;
	wire new_net_3744;
	wire new_net_3078;
	wire new_net_2578;
	wire new_net_2847;
	wire new_net_4982;
	wire new_net_5172;
	wire new_net_5691;
	wire new_net_6840;
	wire new_net_7757;
	wire new_net_7554;
	wire _0110_;
	wire _0320_;
	wire _0824_;
	wire new_net_496;
	wire new_net_1897;
	wire new_net_2828;
	wire new_net_3637;
	wire new_net_2299;
	wire new_net_2715;
	wire _0614_;
	wire new_net_6002;
	wire new_net_7576;
	wire new_net_4900;
	wire new_net_599;
	wire new_net_707;
	wire new_net_2532;
	wire new_net_1946;
	wire new_net_5321;
	wire new_net_7710;
	wire new_net_7783;
	wire new_net_8100;
	wire _0111_;
	wire _0321_;
	wire _0825_;
	wire _0615_;
	wire new_net_636;
	wire new_net_3554;
	wire new_net_4107;
	wire new_net_5446;
	wire new_net_5592;
	wire new_net_5915;
	wire new_net_5617;
	wire new_net_7598;
	wire new_net_5714;
	wire new_net_8139;
	wire new_net_3133;
	wire new_net_1170;
	wire new_net_2848;
	wire new_net_3185;
	wire new_net_5195;
	wire new_net_5298;
	wire new_net_6059;
	wire new_net_6265;
	wire new_net_5963;
	wire new_net_7613;
	wire new_net_5188;
	wire new_net_4523;
	wire new_net_5360;
	wire _0616_;
	wire _0112_;
	wire _0322_;
	wire _0826_;
	wire new_net_1028;
	wire new_net_2268;
	wire new_net_2331;
	wire new_net_3859;
	wire new_net_5095;
	wire new_net_5813;
	wire new_net_4830;
	wire new_net_7675;
	wire new_net_7920;
	wire new_net_600;
	wire new_net_3154;
	wire new_net_3566;
	wire new_net_4889;
	wire new_net_5050;
	wire new_net_5713;
	wire new_net_6279;
	wire new_net_6412;
	wire new_net_6783;
	wire new_net_5665;
	wire new_net_4254;
	wire new_net_5471;
	wire _0617_;
	wire new_net_637;
	wire _0113_;
	wire _0827_;
	wire _0323_;
	wire new_net_2934;
	wire new_net_3745;
	wire new_net_3079;
	wire new_net_2579;
	wire new_net_4556;
	wire new_net_6680;
	wire new_net_7046;
	wire new_net_1171;
	wire new_net_10;
	wire new_net_497;
	wire new_net_3472;
	wire new_net_3638;
	wire new_net_2716;
	wire new_net_3837;
	wire new_net_4045;
	wire new_net_4767;
	wire new_net_4787;
	wire new_net_4392;
	wire new_net_5993;
	wire new_net_6245;
	wire new_net_7312;
	wire new_net_7935;
	wire new_net_8220;
	wire _0828_;
	wire _0114_;
	wire _0324_;
	wire _0618_;
	wire new_net_708;
	wire new_net_1029;
	wire new_net_2300;
	wire new_net_4912;
	wire new_net_5322;
	wire new_net_6329;
	wire new_net_5135;
	wire new_net_5392;
	wire new_net_7157;
	wire new_net_8191;
	wire new_net_1954;
	wire new_net_2614;
	wire new_net_3555;
	wire new_net_4108;
	wire new_net_5447;
	wire new_net_5593;
	wire new_net_5916;
	wire new_net_6864;
	wire new_net_6888;
	wire new_net_6986;
	wire new_net_6717;
	wire new_net_5119;
	wire new_net_4382;
	wire new_net_5943;
	wire new_net_5412;
	wire new_net_7179;
	wire _0829_;
	wire _0115_;
	wire _0619_;
	wire new_net_3134;
	wire new_net_2441;
	wire new_net_2477;
	wire new_net_3186;
	wire _0325_;
	wire new_net_5196;
	wire new_net_6060;
	wire new_net_8257;
	wire new_net_4255;
	wire new_net_7118;
	wire new_net_498;
	wire new_net_1172;
	wire new_net_3473;
	wire new_net_5096;
	wire new_net_5814;
	wire new_net_6659;
	wire new_net_7758;
	wire new_net_7422;
	wire new_net_7712;
	wire _0620_;
	wire _0116_;
	wire _0326_;
	wire new_net_601;
	wire new_net_3155;
	wire new_net_3567;
	wire new_net_709;
	wire _0830_;
	wire new_net_2332;
	wire new_net_2269;
	wire new_net_6192;
	wire new_net_7516;
	wire new_net_7806;
	wire new_net_4505;
	wire new_net_6359;
	wire new_net_3952;
	wire new_net_566;
	wire new_net_638;
	wire new_net_2615;
	wire new_net_2935;
	wire new_net_3080;
	wire new_net_4981;
	wire new_net_5693;
	wire new_net_6842;
	wire new_net_7735;
	wire new_net_6620;
	wire new_net_8068;
	wire new_net_6959;
	wire new_net_2717;
	wire _0621_;
	wire _0117_;
	wire new_net_2643;
	wire new_net_2778;
	wire _0831_;
	wire _0327_;
	wire new_net_3838;
	wire new_net_4046;
	wire new_net_5174;
	wire new_net_5644;
	wire new_net_5611;
	wire new_net_8090;
	wire new_net_4608;
	wire new_net_6146;
	wire new_net_1030;
	wire new_net_1173;
	wire new_net_1951;
	wire new_net_4913;
	wire new_net_5299;
	wire new_net_5323;
	wire new_net_7059;
	wire new_net_6981;
	wire new_net_7535;
	wire new_net_5088;
	wire new_net_5383;
	wire new_net_6570;
	wire new_net_6941;
	wire new_net_6081;
	wire new_net_6079;
	wire _0832_;
	wire _0118_;
	wire new_net_2301;
	wire new_net_602;
	wire _0622_;
	wire new_net_710;
	wire _0328_;
	wire new_net_3860;
	wire new_net_4109;
	wire new_net_5448;
	wire new_net_7744;
	wire new_net_5105;
	wire new_net_7170;
	wire new_net_567;
	wire new_net_639;
	wire new_net_3135;
	wire new_net_2522;
	wire new_net_2644;
	wire new_net_3187;
	wire new_net_2809;
	wire new_net_5197;
	wire new_net_7615;
	wire new_net_7098;
	wire new_net_5783;
	wire _0833_;
	wire _0119_;
	wire new_net_1947;
	wire _0623_;
	wire new_net_3474;
	wire _0329_;
	wire new_net_499;
	wire new_net_1917;
	wire new_net_5097;
	wire new_net_5815;
	wire new_net_6413;
	wire new_net_8020;
	wire new_net_8115;
	wire new_net_6328;
	wire new_net_4622;
	wire new_net_2829;
	wire new_net_1031;
	wire new_net_1174;
	wire new_net_2531;
	wire new_net_3156;
	wire new_net_4788;
	wire new_net_4891;
	wire new_net_5052;
	wire new_net_5715;
	wire new_net_6414;
	wire new_net_6350;
	wire _0330_;
	wire new_net_2936;
	wire new_net_2270;
	wire new_net_3081;
	wire new_net_3753;
	wire _0624_;
	wire _0834_;
	wire _0120_;
	wire new_net_2333;
	wire new_net_2849;
	wire new_net_7352;
	wire new_net_7607;
	wire new_net_6740;
	wire new_net_8059;
	wire new_net_8271;
	wire new_net_7618;
	wire new_net_5883;
	wire new_net_2718;
	wire new_net_3839;
	wire new_net_4047;
	wire new_net_5175;
	wire new_net_5575;
	wire new_net_5917;
	wire new_net_5941;
	wire new_net_6461;
	wire new_net_7387;
	wire new_net_5602;
	wire new_net_8081;
	wire _0331_;
	wire new_net_500;
	wire new_net_3494;
	wire _0625_;
	wire _0121_;
	wire _0835_;
	wire new_net_1835;
	wire new_net_4914;
	wire new_net_5300;
	wire new_net_5324;
	wire new_net_6972;
	wire new_net_7141;
	wire new_net_5871;
	wire new_net_6822;
	wire new_net_1898;
	wire new_net_3502;
	wire new_net_603;
	wire new_net_1032;
	wire new_net_3754;
	wire new_net_1175;
	wire new_net_2580;
	wire new_net_2784;
	wire new_net_3861;
	wire new_net_4110;
	wire new_net_6038;
	wire new_net_4151;
	wire new_net_7902;
	wire new_net_6210;
	wire new_net_7940;
	wire new_net_5306;
	wire new_net_7038;
	wire _0332_;
	wire _0836_;
	wire _0626_;
	wire new_net_568;
	wire new_net_2302;
	wire new_net_2581;
	wire new_net_2850;
	wire new_net_640;
	wire new_net_3136;
	wire _0122_;
	wire new_net_6839;
	wire new_net_7382;
	wire new_net_5774;
	wire new_net_7962;
	wire new_net_6772;
	wire new_net_3475;
	wire new_net_2745;
	wire new_net_5098;
	wire new_net_3218;
	wire new_net_5816;
	wire new_net_4541;
	wire new_net_6266;
	wire new_net_6661;
	wire new_net_7760;
	wire new_net_4256;
	wire new_net_4031;
	wire _0333_;
	wire new_net_501;
	wire new_net_3495;
	wire new_net_3746;
	wire _0837_;
	wire _0627_;
	wire new_net_3556;
	wire _0123_;
	wire new_net_3157;
	wire new_net_4789;
	wire new_net_6169;
	wire new_net_4557;
	wire new_net_8028;
	wire new_net_5930;
	wire new_net_1033;
	wire new_net_604;
	wire new_net_2937;
	wire new_net_3082;
	wire new_net_3760;
	wire new_net_1176;
	wire new_net_5695;
	wire new_net_6844;
	wire new_net_7737;
	wire new_net_5421;
	wire new_net_713;
	wire new_net_2779;
	wire _0628_;
	wire _0838_;
	wire _0334_;
	wire new_net_2271;
	wire new_net_569;
	wire new_net_2719;
	wire new_net_3102;
	wire new_net_2334;
	wire new_net_5588;
	wire new_net_7486;
	wire new_net_7655;
	wire new_net_7282;
	wire new_net_2681;
	wire new_net_5301;
	wire new_net_5325;
	wire new_net_6062;
	wire new_net_7210;
	wire new_net_7537;
	wire new_net_7714;
	wire new_net_8104;
	wire new_net_5161;
	wire new_net_5862;
	wire new_net_6813;
	wire new_net_7436;
	wire new_net_2521;
	wire _0629_;
	wire _0839_;
	wire _0335_;
	wire new_net_502;
	wire _0125_;
	wire new_net_3862;
	wire new_net_4111;
	wire new_net_5450;
	wire new_net_5460;
	wire new_net_7232;
	wire new_net_7230;
	wire new_net_6373;
	wire new_net_4177;
	wire new_net_2646;
	wire new_net_1034;
	wire new_net_3189;
	wire new_net_605;
	wire new_net_3103;
	wire new_net_1177;
	wire new_net_3137;
	wire new_net_5199;
	wire new_net_6020;
	wire new_net_6835;
	wire new_net_8154;
	wire new_net_4869;
	wire new_net_6763;
	wire new_net_714;
	wire new_net_2303;
	wire _0630_;
	wire _0840_;
	wire new_net_3476;
	wire _0336_;
	wire new_net_570;
	wire new_net_642;
	wire _0473_;
	wire _0126_;
	wire new_net_5370;
	wire new_net_6557;
	wire new_net_7314;
	wire new_net_7930;
	wire new_net_1948;
	wire new_net_2682;
	wire new_net_3496;
	wire new_net_2830;
	wire new_net_4790;
	wire new_net_4893;
	wire new_net_5054;
	wire new_net_5576;
	wire new_net_5717;
	wire new_net_5942;
	wire new_net_6579;
	wire new_net_5921;
	wire new_net_3920;
	wire _0857_;
	wire new_net_7336;
	wire new_net_4779;
	wire new_net_7329;
	wire _0127_;
	wire _0337_;
	wire _0841_;
	wire new_net_2938;
	wire new_net_3083;
	wire _0631_;
	wire new_net_3967;
	wire new_net_4769;
	wire new_net_4915;
	wire new_net_5696;
	wire new_net_7562;
	wire new_net_7555;
	wire new_net_1950;
	wire new_net_1178;
	wire new_net_3747;
	wire new_net_2720;
	wire new_net_1991;
	wire new_net_3841;
	wire new_net_4049;
	wire new_net_5177;
	wire new_net_5919;
	wire new_net_7389;
	wire new_net_7407;
	wire new_net_7405;
	wire new_net_4733;
	wire new_net_6003;
	wire new_net_715;
	wire _0128_;
	wire _0338_;
	wire _0842_;
	wire new_net_2272;
	wire new_net_3639;
	wire new_net_571;
	wire new_net_2335;
	wire _0632_;
	wire new_net_4115;
	wire new_net_7494;
	wire new_net_7577;
	wire new_net_7784;
	wire new_net_8201;
	wire new_net_6799;
	wire new_net_503;
	wire new_net_3863;
	wire new_net_4112;
	wire new_net_5099;
	wire new_net_5451;
	wire new_net_5597;
	wire new_net_6868;
	wire new_net_6892;
	wire new_net_5618;
	wire _0633_;
	wire new_net_3138;
	wire new_net_2445;
	wire new_net_3158;
	wire _0129_;
	wire _0339_;
	wire new_net_2481;
	wire new_net_2647;
	wire _0843_;
	wire new_net_1035;
	wire new_net_8140;
	wire new_net_7366;
	wire new_net_5964;
	wire new_net_4524;
	wire new_net_643;
	wire new_net_3477;
	wire new_net_1179;
	wire new_net_5818;
	wire new_net_6268;
	wire new_net_6663;
	wire new_net_7762;
	wire new_net_4831;
	wire new_net_7676;
	wire new_net_3629;
	wire _0634_;
	wire new_net_3557;
	wire _0130_;
	wire _0340_;
	wire new_net_716;
	wire _0844_;
	wire new_net_2683;
	wire new_net_3497;
	wire new_net_572;
	wire new_net_2304;
	wire new_net_3913;
	wire new_net_8101;
	wire new_net_5472;
	wire new_net_3764;
	wire new_net_504;
	wire new_net_1852;
	wire new_net_2939;
	wire new_net_3084;
	wire new_net_4770;
	wire new_net_4916;
	wire new_net_5697;
	wire new_net_6846;
	wire new_net_7739;
	wire new_net_7949;
	wire new_net_607;
	wire new_net_1851;
	wire _0635_;
	wire _0845_;
	wire _0131_;
	wire _0341_;
	wire new_net_1036;
	wire new_net_3748;
	wire new_net_2721;
	wire new_net_3842;
	wire new_net_6681;
	wire new_net_7047;
	wire new_net_5081;
	wire new_net_5994;
	wire new_net_4393;
	wire new_net_6246;
	wire new_net_7313;
	wire new_net_8221;
	wire new_net_3836;
	wire new_net_644;
	wire new_net_3706;
	wire new_net_5303;
	wire new_net_5327;
	wire new_net_6064;
	wire new_net_7539;
	wire new_net_7716;
	wire new_net_8106;
	wire new_net_3834;
	wire new_net_6330;
	wire new_net_5393;
	wire new_net_2336;
	wire _0636_;
	wire _0132_;
	wire _0342_;
	wire new_net_2273;
	wire new_net_717;
	wire _0846_;
	wire new_net_1899;
	wire new_net_573;
	wire new_net_3864;
	wire new_net_6718;
	wire new_net_5944;
	wire new_net_5332;
	wire new_net_7180;
	wire new_net_5330;
	wire new_net_3139;
	wire new_net_2648;
	wire new_net_3191;
	wire new_net_3105;
	wire new_net_5201;
	wire new_net_5577;
	wire new_net_5718;
	wire new_net_6022;
	wire new_net_7619;
	wire new_net_8131;
	wire new_net_2582;
	wire new_net_1180;
	wire new_net_1910;
	wire _0637_;
	wire _0133_;
	wire _0847_;
	wire new_net_1037;
	wire new_net_3478;
	wire _0343_;
	wire new_net_2810;
	wire new_net_7119;
	wire new_net_7423;
	wire new_net_1990;
	wire new_net_3159;
	wire new_net_645;
	wire new_net_1989;
	wire new_net_2684;
	wire new_net_3498;
	wire new_net_2831;
	wire new_net_4792;
	wire new_net_4895;
	wire new_net_5056;
	wire new_net_7880;
	wire new_net_6193;
	wire new_net_7517;
	wire new_net_574;
	wire new_net_2305;
	wire new_net_2851;
	wire _0638_;
	wire new_net_2747;
	wire _0134_;
	wire _0848_;
	wire _0344_;
	wire new_net_505;
	wire new_net_3085;
	wire new_net_5630;
	wire new_net_8069;
	wire new_net_2583;
	wire new_net_2722;
	wire new_net_608;
	wire new_net_2530;
	wire new_net_2520;
	wire new_net_2811;
	wire new_net_3843;
	wire new_net_4051;
	wire new_net_5100;
	wire new_net_5179;
	wire new_net_5893;
	wire new_net_6960;
	wire new_net_6549;
	wire new_net_5652;
	wire new_net_5645;
	wire new_net_5612;
	wire new_net_6232;
	wire new_net_8212;
	wire new_net_1181;
	wire _0849_;
	wire _0135_;
	wire _0639_;
	wire _0345_;
	wire new_net_4609;
	wire new_net_4878;
	wire new_net_5304;
	wire new_net_5212;
	wire new_net_5328;
	wire new_net_6147;
	wire new_net_7060;
	wire new_net_6982;
	wire new_net_5089;
	wire new_net_6571;
	wire new_net_6254;
	wire new_net_646;
	wire new_net_718;
	wire new_net_3865;
	wire new_net_4114;
	wire new_net_5453;
	wire new_net_5599;
	wire new_net_6870;
	wire new_net_7745;
	wire new_net_5106;
	wire new_net_2274;
	wire new_net_575;
	wire new_net_3106;
	wire new_net_2049;
	wire new_net_2337;
	wire _0850_;
	wire _0136_;
	wire _0346_;
	wire _0640_;
	wire new_net_3140;
	wire new_net_4922;
	wire new_net_5823;
	wire new_net_5784;
	wire new_net_609;
	wire new_net_1038;
	wire new_net_3479;
	wire new_net_5820;
	wire new_net_6665;
	wire new_net_7764;
	wire new_net_4810;
	wire new_net_6704;
	wire _0347_;
	wire new_net_3499;
	wire new_net_3160;
	wire _0641_;
	wire new_net_1182;
	wire new_net_3558;
	wire _0137_;
	wire _0851_;
	wire new_net_4793;
	wire new_net_4896;
	wire new_net_7994;
	wire new_net_6184;
	wire new_net_6520;
	wire new_net_5043;
	wire new_net_647;
	wire new_net_719;
	wire new_net_3086;
	wire new_net_3755;
	wire new_net_4772;
	wire new_net_4918;
	wire new_net_5699;
	wire new_net_6112;
	wire new_net_6848;
	wire new_net_7741;
	wire new_net_7353;
	wire new_net_5951;
	wire new_net_7608;
	wire new_net_8060;
	wire new_net_5176;
	wire new_net_8272;
	wire _0348_;
	wire new_net_2812;
	wire new_net_576;
	wire new_net_2306;
	wire new_net_2584;
	wire _0642_;
	wire _0138_;
	wire new_net_2723;
	wire _0852_;
	wire new_net_3844;
	wire new_net_6913;
	wire new_net_6462;
	wire new_net_6051;
	wire new_net_2775;
	wire new_net_1039;
	wire new_net_1961;
	wire new_net_5305;
	wire new_net_5198;
	wire new_net_5329;
	wire new_net_5719;
	wire new_net_6066;
	wire new_net_7541;
	wire new_net_7718;
	wire new_net_8082;
	wire new_net_7142;
	wire _0654_;
	wire _0349_;
	wire new_net_3756;
	wire new_net_3527;
	wire _0853_;
	wire _0643_;
	wire new_net_1183;
	wire new_net_1955;
	wire new_net_2616;
	wire new_net_3559;
	wire _0139_;
	wire new_net_5872;
	wire new_net_6823;
	wire new_net_7736;
	wire new_net_7903;
	wire new_net_7941;
	wire new_net_4365;
	wire new_net_6211;
	wire new_net_3193;
	wire new_net_507;
	wire new_net_648;
	wire new_net_3107;
	wire new_net_3141;
	wire new_net_2650;
	wire new_net_5203;
	wire new_net_5579;
	wire new_net_6024;
	wire new_net_6419;
	wire new_net_5809;
	wire _0350_;
	wire new_net_2275;
	wire _0854_;
	wire new_net_577;
	wire new_net_610;
	wire new_net_2338;
	wire _0644_;
	wire _0140_;
	wire new_net_5821;
	wire new_net_6666;
	wire new_net_6690;
	wire new_net_6773;
	wire new_net_8007;
	wire new_net_6862;
	wire new_net_6784;
	wire new_net_7980;
	wire new_net_3500;
	wire new_net_3749;
	wire new_net_2832;
	wire new_net_1040;
	wire new_net_4794;
	wire new_net_4897;
	wire new_net_5946;
	wire new_net_6791;
	wire new_net_6170;
	wire new_net_7078;
	wire new_net_4484;
	wire new_net_8029;
	wire new_net_4006;
	wire new_net_3930;
	wire new_net_720;
	wire _0351_;
	wire new_net_3087;
	wire _0645_;
	wire _0855_;
	wire new_net_2765;
	wire _0141_;
	wire new_net_4773;
	wire new_net_4919;
	wire new_net_4535;
	wire new_net_1900;
	wire new_net_2813;
	wire new_net_508;
	wire new_net_649;
	wire new_net_1994;
	wire new_net_2585;
	wire new_net_1969;
	wire new_net_2748;
	wire new_net_3845;
	wire new_net_4053;
	wire new_net_4976;
	wire new_net_7111;
	wire new_net_7487;
	wire new_net_4230;
	wire new_net_7656;
	wire new_net_6499;
	wire new_net_3707;
	wire _0856_;
	wire _0352_;
	wire _0646_;
	wire _0142_;
	wire new_net_2307;
	wire new_net_2685;
	wire new_net_11;
	wire new_net_611;
	wire new_net_1962;
	wire new_net_5189;
	wire new_net_3858;
	wire new_net_4096;
	wire new_net_3903;
	wire new_net_1041;
	wire new_net_1184;
	wire new_net_1984;
	wire new_net_3867;
	wire new_net_4116;
	wire new_net_5455;
	wire new_net_5601;
	wire new_net_6271;
	wire new_net_6814;
	wire new_net_6872;
	wire new_net_7437;
	wire new_net_5461;
	wire new_net_7233;
	wire new_net_7231;
	wire new_net_6207;
	wire new_net_7700;
	wire _0143_;
	wire new_net_2449;
	wire new_net_3161;
	wire new_net_721;
	wire new_net_2485;
	wire new_net_2651;
	wire new_net_3194;
	wire new_net_3142;
	wire new_net_2749;
	wire _0353_;
	wire new_net_4663;
	wire new_net_7867;
	wire new_net_8155;
	wire new_net_5690;
	wire new_net_2686;
	wire new_net_2780;
	wire new_net_3708;
	wire new_net_578;
	wire new_net_650;
	wire new_net_4980;
	wire new_net_5822;
	wire new_net_6667;
	wire new_net_7766;
	wire new_net_6396;
	wire new_net_5371;
	wire new_net_6558;
	wire new_net_7315;
	wire _0144_;
	wire _0354_;
	wire new_net_3501;
	wire _0858_;
	wire _0648_;
	wire new_net_2276;
	wire new_net_612;
	wire new_net_2339;
	wire new_net_4795;
	wire new_net_4898;
	wire new_net_7931;
	wire new_net_5922;
	wire new_net_8111;
	wire new_net_1042;
	wire new_net_1185;
	wire new_net_3088;
	wire new_net_5701;
	wire new_net_6850;
	wire new_net_7337;
	wire new_net_7330;
	wire new_net_7743;
	wire new_net_7759;
	wire _0145_;
	wire new_net_722;
	wire _0859_;
	wire _0355_;
	wire new_net_509;
	wire new_net_2814;
	wire new_net_2586;
	wire new_net_2852;
	wire _0649_;
	wire new_net_1909;
	wire new_net_3822;
	wire new_net_7408;
	wire new_net_579;
	wire new_net_651;
	wire new_net_5058;
	wire new_net_5307;
	wire new_net_5331;
	wire new_net_4401;
	wire new_net_6068;
	wire new_net_7543;
	wire new_net_7720;
	wire new_net_8110;
	wire new_net_7578;
	wire new_net_4902;
	wire new_net_8202;
	wire _0146_;
	wire new_net_3568;
	wire _0650_;
	wire _0860_;
	wire _0356_;
	wire new_net_2308;
	wire new_net_3528;
	wire new_net_613;
	wire new_net_3868;
	wire new_net_4117;
	wire new_net_6800;
	wire new_net_5452;
	wire new_net_7600;
	wire new_net_5619;
	wire new_net_7807;
	wire new_net_2750;
	wire new_net_3143;
	wire new_net_2652;
	wire new_net_3195;
	wire new_net_1043;
	wire new_net_3109;
	wire new_net_5205;
	wire new_net_6026;
	wire new_net_6421;
	wire new_net_6610;
	wire new_net_7225;
	wire new_net_6989;
	wire new_net_5023;
	wire _0147_;
	wire new_net_3480;
	wire new_net_723;
	wire _0861_;
	wire _0651_;
	wire _0357_;
	wire new_net_510;
	wire new_net_3761;
	wire new_net_2687;
	wire new_net_4920;
	wire new_net_8281;
	wire new_net_2098;
	wire new_net_3162;
	wire new_net_3569;
	wire new_net_580;
	wire new_net_652;
	wire new_net_1918;
	wire new_net_4796;
	wire new_net_4899;
	wire new_net_5948;
	wire new_net_6793;
	wire new_net_5667;
	wire new_net_8102;
	wire new_net_4303;
	wire new_net_7950;
	wire new_net_6682;
	wire new_net_7048;
	wire new_net_2109;
	wire new_net_2537;
	wire new_net_2561;
	wire new_net_671;
	wire new_net_2172;
	wire _0400_;
	wire _1114_;
	wire _0904_;
	wire new_net_461;
	wire new_net_2235;
	wire new_net_5903;
	wire new_net_4318;
	wire new_net_6247;
	wire new_net_8222;
	wire new_net_528;
	wire new_net_846;
	wire new_net_915;
	wire new_net_990;
	wire new_net_1346;
	wire new_net_1556;
	wire new_net_1736;
	wire new_net_1097;
	wire new_net_4531;
	wire new_net_5116;
	wire new_net_6331;
	wire new_net_133;
	wire new_net_1383;
	wire new_net_1203;
	wire new_net_1416;
	wire new_net_952;
	wire new_net_1825;
	wire _0401_;
	wire _0905_;
	wire _1115_;
	wire new_net_778;
	wire new_net_5121;
	wire new_net_4384;
	wire new_net_5945;
	wire new_net_4645;
	wire new_net_7181;
	wire new_net_4984;
	wire new_net_8132;
	wire new_net_200;
	wire new_net_881;
	wire new_net_2024;
	wire new_net_3881;
	wire new_net_4130;
	wire new_net_4995;
	wire new_net_5038;
	wire new_net_5469;
	wire new_net_6139;
	wire new_net_7027;
	wire new_net_2598;
	wire new_net_2141;
	wire _0402_;
	wire _0906_;
	wire _1116_;
	wire new_net_234;
	wire new_net_462;
	wire new_net_813;
	wire new_net_4808;
	wire new_net_5017;
	wire new_net_7002;
	wire new_net_6886;
	wire new_net_5855;
	wire new_net_7424;
	wire new_net_1827;
	wire new_net_1881;
	wire new_net_916;
	wire new_net_991;
	wire new_net_1347;
	wire new_net_1557;
	wire new_net_1098;
	wire new_net_3815;
	wire new_net_4219;
	wire new_net_5343;
	wire new_net_7881;
	wire new_net_6194;
	wire new_net_7518;
	wire new_net_4574;
	wire new_net_4507;
	wire new_net_6361;
	wire new_net_3954;
	wire new_net_5631;
	wire new_net_3512;
	wire new_net_134;
	wire new_net_1384;
	wire new_net_1826;
	wire new_net_1204;
	wire new_net_1417;
	wire new_net_953;
	wire _1117_;
	wire _0403_;
	wire _0907_;
	wire new_net_5755;
	wire new_net_6622;
	wire new_net_8070;
	wire new_net_201;
	wire new_net_672;
	wire new_net_1936;
	wire new_net_4087;
	wire new_net_4972;
	wire new_net_5138;
	wire new_net_5894;
	wire new_net_6961;
	wire new_net_7635;
	wire new_net_7977;
	wire new_net_5646;
	wire new_net_5981;
	wire new_net_5291;
	wire new_net_6155;
	wire new_net_8092;
	wire new_net_6148;
	wire new_net_529;
	wire new_net_847;
	wire new_net_1931;
	wire new_net_2377;
	wire new_net_3117;
	wire new_net_2110;
	wire _0404_;
	wire _1118_;
	wire _0908_;
	wire new_net_235;
	wire new_net_5213;
	wire new_net_6983;
	wire new_net_7533;
	wire new_net_4148;
	wire new_net_5385;
	wire new_net_6572;
	wire new_net_6083;
	wire new_net_779;
	wire new_net_992;
	wire new_net_1558;
	wire new_net_6082;
	wire new_net_6908;
	wire new_net_7006;
	wire new_net_7557;
	wire new_net_8124;
	wire new_net_7746;
	wire new_net_8031;
	wire new_net_5107;
	wire _1180_;
	wire new_net_7172;
	wire new_net_882;
	wire new_net_1205;
	wire new_net_1418;
	wire _0909_;
	wire _0405_;
	wire _1119_;
	wire new_net_954;
	wire new_net_3882;
	wire new_net_4131;
	wire new_net_4996;
	wire new_net_5252;
	wire new_net_673;
	wire new_net_814;
	wire new_net_4809;
	wire new_net_5018;
	wire new_net_5219;
	wire new_net_5961;
	wire new_net_6415;
	wire new_net_6703;
	wire new_net_6705;
	wire new_net_6806;
	wire new_net_4624;
	wire new_net_1348;
	wire new_net_2032;
	wire new_net_530;
	wire new_net_1099;
	wire new_net_848;
	wire new_net_3118;
	wire new_net_917;
	wire _0910_;
	wire _0406_;
	wire _1120_;
	wire new_net_6185;
	wire new_net_7678;
	wire new_net_5533;
	wire new_net_6352;
	wire new_net_5044;
	wire new_net_1064;
	wire new_net_1559;
	wire new_net_1385;
	wire new_net_135;
	wire new_net_780;
	wire new_net_993;
	wire new_net_1758;
	wire new_net_4516;
	wire new_net_6113;
	wire new_net_6163;
	wire new_net_7354;
	wire new_net_6742;
	wire new_net_8061;
	wire new_net_8273;
	wire new_net_7620;
	wire _1121_;
	wire new_net_883;
	wire _0407_;
	wire _0911_;
	wire new_net_1206;
	wire new_net_202;
	wire new_net_955;
	wire new_net_4088;
	wire new_net_4973;
	wire new_net_5139;
	wire new_net_5885;
	wire new_net_6463;
	wire new_net_8083;
	wire new_net_0;
	wire new_net_674;
	wire new_net_815;
	wire new_net_4533;
	wire new_net_5118;
	wire new_net_4420;
	wire new_net_5836;
	wire new_net_7835;
	wire new_net_7143;
	wire new_net_4464;
	wire new_net_465;
	wire new_net_1349;
	wire new_net_2237;
	wire new_net_531;
	wire new_net_1100;
	wire _1122_;
	wire _0408_;
	wire _0912_;
	wire new_net_918;
	wire new_net_2111;
	wire new_net_6040;
	wire new_net_6824;
	wire new_net_7904;
	wire new_net_4366;
	wire new_net_6212;
	wire new_net_7942;
	wire new_net_4190;
	wire new_net_1065;
	wire new_net_1560;
	wire new_net_1386;
	wire new_net_136;
	wire new_net_781;
	wire new_net_994;
	wire new_net_1419;
	wire new_net_1983;
	wire new_net_3172;
	wire new_net_3883;
	wire new_net_6841;
	wire new_net_7966;
	wire new_net_7964;
	wire new_net_6774;
	wire new_net_2070;
	wire new_net_2700;
	wire _0409_;
	wire _1123_;
	wire _0913_;
	wire new_net_2600;
	wire new_net_1207;
	wire new_net_203;
	wire new_net_956;
	wire new_net_3173;
	wire new_net_6691;
	wire new_net_6863;
	wire new_net_5834;
	wire new_net_6785;
	wire new_net_5832;
	wire new_net_7981;
	wire new_net_237;
	wire new_net_675;
	wire new_net_849;
	wire new_net_3119;
	wire new_net_3817;
	wire new_net_4229;
	wire new_net_4551;
	wire new_net_5345;
	wire new_net_6039;
	wire new_net_7490;
	wire new_net_6171;
	wire new_net_4561;
	wire new_net_7495;
	wire new_net_6979;
	wire new_net_8030;
	wire new_net_466;
	wire new_net_532;
	wire new_net_1919;
	wire new_net_1819;
	wire _0410_;
	wire _1124_;
	wire _0914_;
	wire new_net_1350;
	wire new_net_919;
	wire new_net_2143;
	wire new_net_3108;
	wire new_net_1561;
	wire new_net_782;
	wire new_net_884;
	wire new_net_1420;
	wire new_net_4089;
	wire new_net_5140;
	wire new_net_7637;
	wire new_net_7979;
	wire new_net_8149;
	wire new_net_5590;
	wire new_net_7657;
	wire new_net_7284;
	wire new_net_6500;
	wire new_net_5190;
	wire new_net_2379;
	wire new_net_816;
	wire new_net_2701;
	wire _0411_;
	wire _0915_;
	wire _1125_;
	wire new_net_1208;
	wire new_net_204;
	wire new_net_957;
	wire new_net_4534;
	wire new_net_7212;
	wire new_net_7129;
	wire new_net_5864;
	wire new_net_3513;
	wire new_net_238;
	wire new_net_676;
	wire new_net_850;
	wire new_net_1101;
	wire new_net_4231;
	wire new_net_4552;
	wire new_net_5019;
	wire new_net_6084;
	wire new_net_6815;
	wire new_net_7438;
	wire new_net_5462;
	wire new_net_7234;
	wire new_net_7701;
	wire new_net_6375;
	wire new_net_995;
	wire new_net_2175;
	wire new_net_2238;
	wire new_net_467;
	wire new_net_1066;
	wire new_net_1351;
	wire new_net_2031;
	wire new_net_533;
	wire _1126_;
	wire _0412_;
	wire new_net_6837;
	wire new_net_8156;
	wire new_net_4871;
	wire new_net_6765;
	wire new_net_1732;
	wire new_net_1562;
	wire new_net_783;
	wire new_net_1932;
	wire new_net_885;
	wire new_net_303;
	wire new_net_2601;
	wire new_net_1743;
	wire new_net_4811;
	wire new_net_5221;
	wire new_net_6397;
	wire new_net_5372;
	wire new_net_4844;
	wire new_net_3715;
	wire new_net_7932;
	wire new_net_958;
	wire new_net_2099;
	wire new_net_1888;
	wire new_net_817;
	wire _1127_;
	wire _0413_;
	wire _0917_;
	wire new_net_3120;
	wire new_net_1209;
	wire new_net_3818;
	wire new_net_6581;
	wire new_net_5923;
	wire new_net_8112;
	wire new_net_4266;
	wire new_net_7459;
	wire new_net_4264;
	wire new_net_1811;
	wire new_net_1834;
	wire new_net_2562;
	wire new_net_3514;
	wire new_net_239;
	wire new_net_677;
	wire new_net_1102;
	wire new_net_2730;
	wire new_net_3917;
	wire new_net_3969;
	wire new_net_4781;
	wire new_net_1943;
	wire new_net_7564;
	wire new_net_1421;
	wire new_net_2144;
	wire new_net_996;
	wire new_net_1067;
	wire new_net_1352;
	wire _0918_;
	wire _1128_;
	wire _0414_;
	wire new_net_1737;
	wire new_net_138;
	wire new_net_3219;
	wire new_net_4803;
	wire new_net_6491;
	wire new_net_7409;
	wire new_net_4735;
	wire new_net_6005;
	wire new_net_205;
	wire new_net_1563;
	wire new_net_2702;
	wire new_net_3900;
	wire new_net_4220;
	wire new_net_5120;
	wire new_net_5838;
	wire new_net_7837;
	wire new_net_7120;
	wire new_net_7786;
	wire _1182_;
	wire new_net_8203;
	wire new_net_6801;
	wire new_net_959;
	wire new_net_2427;
	wire new_net_1968;
	wire _0919_;
	wire _0415_;
	wire new_net_2563;
	wire new_net_1210;
	wire _0202_;
	wire new_net_851;
	wire _1129_;
	wire new_net_5620;
	wire new_net_2731;
	wire new_net_240;
	wire new_net_468;
	wire new_net_534;
	wire new_net_678;
	wire new_net_921;
	wire new_net_3885;
	wire new_net_4134;
	wire new_net_4999;
	wire new_net_5473;
	wire new_net_8142;
	wire new_net_7368;
	wire new_net_5966;
	wire new_net_6712;
	wire new_net_886;
	wire new_net_1422;
	wire new_net_2113;
	wire new_net_2239;
	wire new_net_2176;
	wire new_net_784;
	wire new_net_1068;
	wire new_net_1353;
	wire _1130_;
	wire _0920_;
	wire new_net_1780;
	wire new_net_8164;
	wire new_net_6644;
	wire new_net_1975;
	wire new_net_206;
	wire new_net_818;
	wire new_net_3819;
	wire new_net_5347;
	wire new_net_4610;
	wire new_net_6041;
	wire new_net_7492;
	wire new_net_8048;
	wire new_net_8103;
	wire new_net_5474;
	wire new_net_1211;
	wire new_net_960;
	wire new_net_3174;
	wire new_net_1778;
	wire _1131_;
	wire _0417_;
	wire _0921_;
	wire new_net_2041;
	wire new_net_1103;
	wire new_net_3515;
	wire new_net_3234;
	wire new_net_4086;
	wire new_net_1389;
	wire new_net_2053;
	wire new_net_139;
	wire new_net_469;
	wire new_net_535;
	wire new_net_679;
	wire new_net_922;
	wire new_net_997;
	wire new_net_4091;
	wire new_net_4530;
	wire new_net_6322;
	wire new_net_6683;
	wire new_net_4395;
	wire new_net_887;
	wire new_net_2381;
	wire new_net_2145;
	wire _0922_;
	wire _1132_;
	wire _0418_;
	wire new_net_785;
	wire new_net_1069;
	wire new_net_1354;
	wire new_net_1564;
	wire new_net_8223;
	wire new_net_6332;
	wire new_net_5395;
	wire new_net_6093;
	wire new_net_1745;
	wire new_net_207;
	wire new_net_819;
	wire new_net_5021;
	wire new_net_6086;
	wire new_net_6912;
	wire new_net_7010;
	wire new_net_7283;
	wire new_net_7561;
	wire new_net_7860;
	wire new_net_5240;
	wire new_net_4385;
	wire new_net_5334;
	wire new_net_7182;
	wire new_net_853;
	wire new_net_1212;
	wire new_net_961;
	wire new_net_241;
	wire _0923_;
	wire _1133_;
	wire _0419_;
	wire new_net_1104;
	wire new_net_3886;
	wire new_net_4135;
	wire new_net_8133;
	wire new_net_7609;
	wire new_net_140;
	wire new_net_680;
	wire new_net_998;
	wire new_net_1390;
	wire new_net_1423;
	wire new_net_1790;
	wire new_net_4519;
	wire new_net_4813;
	wire new_net_5223;
	wire new_net_5965;
	wire new_net_7003;
	wire new_net_6887;
	wire new_net_7833;
	wire new_net_6514;
	wire new_net_5856;
	wire new_net_2114;
	wire new_net_1886;
	wire new_net_2177;
	wire _0420_;
	wire _1134_;
	wire _0924_;
	wire new_net_786;
	wire new_net_1070;
	wire new_net_1355;
	wire new_net_1565;
	wire new_net_7425;
	wire new_net_7715;
	wire new_net_7882;
	wire new_net_7519;
	wire new_net_4580;
	wire new_net_6362;
	wire new_net_3516;
	wire new_net_3919;
	wire new_net_5042;
	wire new_net_6167;
	wire new_net_6191;
	wire new_net_6289;
	wire new_net_6536;
	wire new_net_6684;
	wire new_net_7134;
	wire new_net_7412;
	wire new_net_5632;
	wire new_net_615;
	wire new_net_3306;
	wire new_net_8071;
	wire new_net_536;
	wire new_net_2564;
	wire new_net_1793;
	wire new_net_923;
	wire new_net_1213;
	wire new_net_242;
	wire _0421_;
	wire _1135_;
	wire _0925_;
	wire new_net_470;
	wire new_net_6962;
	wire new_net_5895;
	wire new_net_2746;
	wire new_net_3121;
	wire new_net_681;
	wire new_net_888;
	wire new_net_1424;
	wire new_net_3902;
	wire new_net_4537;
	wire new_net_4554;
	wire new_net_4606;
	wire new_net_5122;
	wire new_net_5840;
	wire new_net_6149;
	wire new_net_8093;
	wire new_net_5214;
	wire new_net_5091;
	wire new_net_6573;
	wire new_net_787;
	wire new_net_1071;
	wire new_net_1356;
	wire new_net_820;
	wire new_net_1960;
	wire new_net_1566;
	wire new_net_208;
	wire new_net_2146;
	wire _0926_;
	wire _0422_;
	wire new_net_7747;
	wire new_net_8032;
	wire new_net_7079;
	wire new_net_5108;
	wire new_net_1062;
	wire new_net_2548;
	wire new_net_7173;
	wire new_net_2565;
	wire new_net_1967;
	wire new_net_854;
	wire new_net_962;
	wire new_net_1105;
	wire new_net_3887;
	wire new_net_5001;
	wire new_net_5475;
	wire new_net_7033;
	wire new_net_4924;
	wire new_net_5253;
	wire new_net_7101;
	wire new_net_5786;
	wire new_net_1959;
	wire new_net_537;
	wire new_net_141;
	wire new_net_1391;
	wire new_net_2602;
	wire new_net_924;
	wire new_net_1214;
	wire _0927_;
	wire _0423_;
	wire _1137_;
	wire new_net_6416;
	wire new_net_4812;
	wire new_net_6706;
	wire new_net_1768;
	wire new_net_4441;
	wire new_net_2549;
	wire new_net_1926;
	wire new_net_2703;
	wire new_net_889;
	wire new_net_5349;
	wire new_net_6043;
	wire new_net_37;
	wire new_net_3739;
	wire new_net_7996;
	wire new_net_5534;
	wire new_net_4097;
	wire new_net_6522;
	wire new_net_1072;
	wire new_net_1357;
	wire new_net_1567;
	wire new_net_2241;
	wire new_net_821;
	wire new_net_2008;
	wire new_net_3517;
	wire new_net_2115;
	wire new_net_209;
	wire _0424_;
	wire new_net_4290;
	wire new_net_4288;
	wire new_net_6114;
	wire new_net_7355;
	wire new_net_5953;
	wire new_net_7534;
	wire new_net_137;
	wire new_net_8062;
	wire new_net_5178;
	wire new_net_1106;
	wire new_net_243;
	wire new_net_855;
	wire new_net_963;
	wire new_net_5022;
	wire new_net_5144;
	wire new_net_6834;
	wire new_net_7621;
	wire new_net_7641;
	wire new_net_7983;
	wire new_net_8274;
	wire new_net_6464;
	wire new_net_6053;
	wire new_net_2074;
	wire new_net_2100;
	wire new_net_538;
	wire new_net_142;
	wire new_net_1392;
	wire new_net_1215;
	wire new_net_1425;
	wire new_net_2383;
	wire _0425_;
	wire _1139_;
	wire _0929_;
	wire new_net_2776;
	wire new_net_5200;
	wire new_net_8084;
	wire new_net_6559;
	wire new_net_7144;
	wire new_net_2097;
	wire new_net_788;
	wire new_net_890;
	wire new_net_4232;
	wire new_net_6088;
	wire new_net_6914;
	wire new_net_7012;
	wire new_net_7285;
	wire new_net_7563;
	wire new_net_7862;
	wire new_net_6825;
	wire new_net_5796;
	wire new_net_7738;
	wire new_net_7244;
	wire new_net_7905;
	wire new_net_6213;
	wire _0930_;
	wire new_net_1073;
	wire new_net_1820;
	wire _0426_;
	wire _1140_;
	wire new_net_1334;
	wire new_net_2147;
	wire new_net_3888;
	wire new_net_5002;
	wire new_net_5476;
	wire new_net_6670;
	wire new_net_698;
	wire new_net_3353;
	wire new_net_5811;
	wire new_net_7967;
	wire new_net_7965;
	wire new_net_1107;
	wire new_net_1944;
	wire new_net_244;
	wire new_net_472;
	wire new_net_1738;
	wire new_net_925;
	wire new_net_964;
	wire new_net_4815;
	wire new_net_5225;
	wire new_net_5967;
	wire new_net_1777;
	wire new_net_5835;
	wire new_net_3876;
	wire new_net_6786;
	wire new_net_5833;
	wire new_net_539;
	wire new_net_143;
	wire new_net_1216;
	wire new_net_1426;
	wire _0931_;
	wire _0427_;
	wire _1141_;
	wire new_net_683;
	wire new_net_5350;
	wire new_net_6044;
	wire new_net_7982;
	wire new_net_7498;
	wire new_net_2455;
	wire new_net_6172;
	wire new_net_7496;
	wire new_net_3932;
	wire new_net_1568;
	wire new_net_2044;
	wire new_net_3518;
	wire new_net_2732;
	wire new_net_210;
	wire new_net_789;
	wire new_net_891;
	wire new_net_1358;
	wire new_net_3921;
	wire new_net_4521;
	wire new_net_3979;
	wire new_net_7808;
	wire new_net_2179;
	wire new_net_1074;
	wire new_net_2242;
	wire new_net_823;
	wire new_net_2704;
	wire _0932_;
	wire _0428_;
	wire _1142_;
	wire new_net_2116;
	wire new_net_2021;
	wire new_net_7113;
	wire new_net_338;
	wire new_net_4550;
	wire new_net_6990;
	wire new_net_1001;
	wire new_net_1393;
	wire new_net_2101;
	wire new_net_245;
	wire new_net_473;
	wire new_net_857;
	wire new_net_926;
	wire new_net_1679;
	wire new_net_3904;
	wire new_net_4539;
	wire new_net_4745;
	wire _0042_;
	wire new_net_7130;
	wire new_net_6432;
	wire new_net_684;
	wire new_net_2733;
	wire _0429_;
	wire _1143_;
	wire _0933_;
	wire new_net_1217;
	wire new_net_3820;
	wire new_net_3905;
	wire new_net_6089;
	wire new_net_6915;
	wire new_net_6816;
	wire new_net_5124;
	wire new_net_7439;
	wire new_net_5463;
	wire new_net_7235;
	wire new_net_2048;
	wire new_net_1569;
	wire new_net_2073;
	wire new_net_211;
	wire new_net_892;
	wire new_net_1359;
	wire new_net_3889;
	wire new_net_4137;
	wire new_net_5003;
	wire new_net_5477;
	wire new_net_4665;
	wire new_net_7869;
	wire new_net_6838;
	wire new_net_8157;
	wire new_net_1923;
	wire new_net_7951;
	wire new_net_5692;
	wire new_net_965;
	wire new_net_2148;
	wire new_net_1075;
	wire new_net_824;
	wire new_net_1108;
	wire new_net_2096;
	wire _0430_;
	wire _1144_;
	wire _0934_;
	wire new_net_2425;
	wire new_net_6027;
	wire new_net_6398;
	wire new_net_7317;
	wire new_net_1427;
	wire new_net_144;
	wire new_net_246;
	wire new_net_474;
	wire new_net_540;
	wire new_net_858;
	wire new_net_1002;
	wire new_net_1394;
	wire new_net_4094;
	wire new_net_5351;
	wire new_net_5513;
	wire new_net_6582;
	wire new_net_5924;
	wire new_net_8113;
	wire new_net_7460;
	wire new_net_1218;
	wire new_net_1953;
	wire new_net_685;
	wire new_net_790;
	wire new_net_2075;
	wire new_net_3519;
	wire _0935_;
	wire _0431_;
	wire _1145_;
	wire new_net_3922;
	wire new_net_7339;
	wire new_net_4782;
	wire new_net_7332;
	wire new_net_7761;
	wire new_net_7267;
	wire new_net_1807;
	wire new_net_1570;
	wire new_net_2705;
	wire new_net_212;
	wire new_net_4222;
	wire new_net_3328;
	wire new_net_5024;
	wire new_net_5146;
	wire new_net_6443;
	wire new_net_6836;
	wire new_net_7565;
	wire new_net_7410;
	wire new_net_927;
	wire new_net_2117;
	wire new_net_2385;
	wire new_net_966;
	wire new_net_2180;
	wire new_net_1733;
	wire new_net_1076;
	wire new_net_2243;
	wire new_net_1109;
	wire new_net_2566;
	wire new_net_2151;
	wire new_net_6006;
	wire new_net_4904;
	wire new_net_7121;
	wire new_net_7787;
	wire new_net_1063;
	wire new_net_2734;
	wire new_net_1428;
	wire new_net_2569;
	wire new_net_145;
	wire new_net_247;
	wire new_net_541;
	wire new_net_1003;
	wire new_net_1395;
	wire new_net_6090;
	wire new_net_6802;
	wire new_net_5454;
	wire new_net_6195;
	wire new_net_5621;
	wire new_net_1219;
	wire new_net_791;
	wire new_net_1360;
	wire new_net_1814;
	wire _0433_;
	wire _1147_;
	wire _0937_;
	wire new_net_3890;
	wire new_net_4138;
	wire new_net_5004;
	wire new_net_4975;
	wire new_net_8143;
	wire new_net_342;
	wire new_net_1114;
	wire new_net_4701;
	wire new_net_2353;
	wire new_net_1571;
	wire new_net_1815;
	wire new_net_2043;
	wire new_net_213;
	wire new_net_825;
	wire new_net_4522;
	wire new_net_4817;
	wire new_net_5227;
	wire new_net_5969;
	wire new_net_6687;
	wire new_net_38;
	wire new_net_5364;
	wire new_net_6551;
	wire new_net_8165;
	wire new_net_928;
	wire new_net_2149;
	wire new_net_475;
	wire new_net_2550;
	wire new_net_1110;
	wire new_net_2567;
	wire _0434_;
	wire _1148_;
	wire _0938_;
	wire new_net_1715;
	wire new_net_2079;
	wire new_net_2046;
	wire new_net_3520;
	wire new_net_248;
	wire new_net_542;
	wire new_net_686;
	wire new_net_1004;
	wire new_net_1396;
	wire new_net_1721;
	wire new_net_2034;
	wire new_net_3923;
	wire new_net_4304;
	wire new_net_1929;
	wire new_net_3242;
	wire _1186_;
	wire new_net_2866;
	wire new_net_1839;
	wire new_net_894;
	wire new_net_1220;
	wire new_net_1361;
	wire _0939_;
	wire _0435_;
	wire _1149_;
	wire new_net_920;
	wire new_net_5025;
	wire new_net_5147;
	wire _0206_;
	wire new_net_396;
	wire new_net_3122;
	wire new_net_1077;
	wire new_net_1572;
	wire new_net_2551;
	wire new_net_214;
	wire new_net_826;
	wire new_net_1727;
	wire new_net_664;
	wire new_net_3821;
	wire new_net_3906;
	wire new_net_8224;
	wire new_net_860;
	wire _1150_;
	wire new_net_146;
	wire new_net_929;
	wire new_net_1429;
	wire new_net_2118;
	wire new_net_968;
	wire new_net_2181;
	wire new_net_476;
	wire new_net_2244;
	wire _0174_;
	wire new_net_699;
	wire new_net_5241;
	wire new_net_7679;
	wire new_net_6721;
	wire new_net_5123;
	wire new_net_249;
	wire new_net_543;
	wire new_net_687;
	wire new_net_792;
	wire new_net_1005;
	wire new_net_1397;
	wire new_net_2087;
	wire new_net_3891;
	wire new_net_4139;
	wire new_net_5947;
	wire new_net_4647;
	wire new_net_7183;
	wire new_net_7768;
	wire new_net_7610;
	wire new_net_4360;
	wire new_net_6127;
	wire new_net_1884;
	wire new_net_1945;
	wire new_net_895;
	wire new_net_2603;
	wire new_net_1221;
	wire new_net_1362;
	wire new_net_1739;
	wire new_net_1992;
	wire _0437_;
	wire _1151_;
	wire new_net_7195;
	wire new_net_7200;
	wire new_net_5525;
	wire new_net_7004;
	wire new_net_7834;
	wire new_net_2568;
	wire new_net_1837;
	wire new_net_3123;
	wire new_net_2102;
	wire new_net_1078;
	wire new_net_1573;
	wire new_net_215;
	wire new_net_827;
	wire new_net_3897;
	wire new_net_5353;
	wire new_net_5857;
	wire new_net_7426;
	wire new_net_7522;
	wire new_net_7883;
	wire new_net_7520;
	wire new_net_4509;
	wire new_net_1112;
	wire new_net_3521;
	wire new_net_147;
	wire new_net_1907;
	wire new_net_930;
	wire new_net_1430;
	wire new_net_969;
	wire new_net_2150;
	wire new_net_3175;
	wire _0438_;
	wire new_net_6363;
	wire new_net_3659;
	wire new_net_5757;
	wire _0876_;
	wire new_net_1786;
	wire new_net_1111;
	wire new_net_1883;
	wire new_net_2045;
	wire new_net_2;
	wire new_net_250;
	wire new_net_544;
	wire new_net_688;
	wire new_net_793;
	wire new_net_1006;
	wire new_net_1398;
	wire new_net_4095;
	wire new_net_8072;
	wire new_net_1680;
	wire new_net_2992;
	wire new_net_3282;
	wire new_net_5130;
	wire new_net_852;
	wire new_net_896;
	wire new_net_1222;
	wire new_net_1801;
	wire new_net_2387;
	wire _0943_;
	wire _0439_;
	wire _1153_;
	wire new_net_3907;
	wire new_net_5005;
	wire new_net_5845;
	wire new_net_6235;
	wire new_net_6775;
	wire new_net_8094;
	wire new_net_5215;
	wire new_net_1746;
	wire new_net_4587;
	wire new_net_1079;
	wire new_net_1574;
	wire new_net_2103;
	wire new_net_477;
	wire new_net_828;
	wire new_net_861;
	wire new_net_4558;
	wire new_net_5228;
	wire new_net_6085;
	wire new_net_6092;
	wire new_net_217;
	wire new_net_5232;
	wire new_net_7748;
	wire _0730_;
	wire new_net_8033;
	wire new_net_7080;
	wire new_net_1759;
	wire new_net_5109;
	wire new_net_2245;
	wire new_net_1113;
	wire new_net_148;
	wire new_net_931;
	wire new_net_2119;
	wire new_net_2182;
	wire _0944_;
	wire _0440_;
	wire _1154_;
	wire new_net_3892;
	wire new_net_7908;
	wire _1080_;
	wire new_net_5254;
	wire new_net_1363;
	wire new_net_1399;
	wire new_net_1783;
	wire new_net_251;
	wire new_net_689;
	wire new_net_1007;
	wire new_net_1302;
	wire new_net_4819;
	wire new_net_5126;
	wire new_net_5478;
	wire new_net_6417;
	wire new_net_6707;
	wire new_net_6501;
	wire new_net_1812;
	wire new_net_1836;
	wire new_net_897;
	wire new_net_3124;
	wire new_net_1223;
	wire new_net_216;
	wire _0441_;
	wire _1155_;
	wire _0945_;
	wire new_net_1788;
	wire new_net_4626;
	wire new_net_2030;
	wire new_net_5164;
	wire new_net_5535;
	wire new_net_1575;
	wire new_net_3522;
	wire new_net_1726;
	wire new_net_1794;
	wire new_net_2735;
	wire new_net_1431;
	wire new_net_478;
	wire new_net_862;
	wire new_net_970;
	wire new_net_3925;
	wire new_net_5046;
	wire new_net_6523;
	wire new_net_7356;
	wire new_net_3151;
	wire new_net_6282;
	wire new_net_7702;
	wire new_net_8063;
	wire new_net_7624;
	wire new_net_8275;
	wire new_net_7622;
	wire new_net_6916;
	wire new_net_4946;
	wire new_net_5887;
	wire new_net_6465;
	wire _0190_;
	wire _0988_;
	wire _1198_;
	wire new_net_1772;
	wire new_net_1591;
	wire _0484_;
	wire _0694_;
	wire new_net_1243;
	wire new_net_1483;
	wire new_net_4278;
	wire new_net_7646;
	wire new_net_6560;
	wire new_net_7145;
	wire new_net_408;
	wire new_net_1824;
	wire new_net_3624;
	wire new_net_1920;
	wire new_net_2965;
	wire new_net_3281;
	wire new_net_4313;
	wire new_net_4619;
	wire new_net_5858;
	wire new_net_6576;
	wire new_net_6826;
	wire new_net_6042;
	wire new_net_7245;
	wire new_net_4372;
	wire new_net_5680;
	wire new_net_6221;
	wire new_net_7906;
	wire new_net_6214;
	wire new_net_7160;
	wire new_net_6671;
	wire _0191_;
	wire _0485_;
	wire _1199_;
	wire new_net_742;
	wire new_net_1889;
	wire _0989_;
	wire new_net_340;
	wire new_net_1662;
	wire _0045_;
	wire new_net_3266;
	wire new_net_6843;
	wire new_net_7968;
	wire new_net_5702;
	wire new_net_95;
	wire new_net_269;
	wire new_net_305;
	wire new_net_1132;
	wire new_net_1315;
	wire new_net_3247;
	wire new_net_2986;
	wire new_net_1699;
	wire new_net_5263;
	wire new_net_5390;
	wire new_net_6865;
	wire new_net_6787;
	wire new_net_4037;
	wire _0192_;
	wire new_net_1280;
	wire new_net_1484;
	wire new_net_2204;
	wire new_net_3206;
	wire _0990_;
	wire new_net_1592;
	wire _0486_;
	wire new_net_3664;
	wire _1200_;
	wire new_net_6173;
	wire new_net_4563;
	wire new_net_7497;
	wire new_net_4494;
	wire new_net_5934;
	wire new_net_409;
	wire new_net_3374;
	wire new_net_2013;
	wire new_net_4640;
	wire new_net_4933;
	wire new_net_5367;
	wire new_net_6554;
	wire new_net_7579;
	wire new_net_7677;
	wire new_net_7878;
	wire new_net_4681;
	wire new_net_4954;
	wire new_net_3570;
	wire _0697_;
	wire _0991_;
	wire _0193_;
	wire new_net_743;
	wire new_net_1891;
	wire _0487_;
	wire new_net_1915;
	wire new_net_341;
	wire new_net_1663;
	wire new_net_7114;
	wire new_net_7659;
	wire new_net_6991;
	wire new_net_7286;
	wire new_net_96;
	wire new_net_270;
	wire new_net_306;
	wire new_net_1133;
	wire new_net_2106;
	wire new_net_3223;
	wire new_net_1700;
	wire new_net_4279;
	wire new_net_4732;
	wire new_net_5162;
	wire new_net_7214;
	wire new_net_7131;
	wire _0194_;
	wire _0698_;
	wire new_net_1245;
	wire new_net_3293;
	wire new_net_1281;
	wire new_net_3625;
	wire new_net_2966;
	wire _0992_;
	wire new_net_1593;
	wire _0488_;
	wire new_net_7440;
	wire new_net_5464;
	wire new_net_7236;
	wire new_net_6296;
	wire new_net_410;
	wire new_net_3267;
	wire new_net_3705;
	wire new_net_4299;
	wire new_net_4641;
	wire new_net_4696;
	wire new_net_4966;
	wire new_net_5984;
	wire new_net_6008;
	wire new_net_7176;
	wire new_net_7870;
	wire new_net_7952;
	wire new_net_3669;
	wire _0489_;
	wire _1203_;
	wire _0195_;
	wire _0699_;
	wire new_net_744;
	wire new_net_1316;
	wire _0993_;
	wire new_net_1833;
	wire new_net_1938;
	wire new_net_6028;
	wire new_net_7318;
	wire new_net_7856;
	wire new_net_97;
	wire new_net_271;
	wire new_net_307;
	wire new_net_1134;
	wire new_net_1485;
	wire new_net_3762;
	wire new_net_3207;
	wire new_net_4019;
	wire new_net_4244;
	wire new_net_5492;
	wire new_net_5514;
	wire new_net_6333;
	wire new_net_4155;
	wire new_net_6583;
	wire new_net_3924;
	wire new_net_8114;
	wire new_net_4268;
	wire _0196_;
	wire _1204_;
	wire _0700_;
	wire new_net_1246;
	wire new_net_3294;
	wire new_net_2205;
	wire _0994_;
	wire new_net_3375;
	wire _0490_;
	wire new_net_3389;
	wire new_net_4783;
	wire new_net_3971;
	wire new_net_7333;
	wire new_net_6433;
	wire new_net_7566;
	wire new_net_411;
	wire new_net_3670;
	wire new_net_2029;
	wire new_net_3939;
	wire new_net_6444;
	wire new_net_7154;
	wire new_net_7779;
	wire new_net_7803;
	wire new_net_7901;
	wire new_net_7411;
	wire new_net_343;
	wire new_net_1665;
	wire _0701_;
	wire _0995_;
	wire _0197_;
	wire _1205_;
	wire new_net_1701;
	wire new_net_3560;
	wire new_net_1317;
	wire _0491_;
	wire new_net_4121;
	wire new_net_4737;
	wire new_net_7790;
	wire new_net_7122;
	wire new_net_7788;
	wire new_net_5151;
	wire new_net_98;
	wire new_net_272;
	wire new_net_308;
	wire new_net_3283;
	wire new_net_1282;
	wire new_net_1486;
	wire new_net_3626;
	wire new_net_1594;
	wire new_net_4333;
	wire new_net_5860;
	wire new_net_6803;
	wire new_net_6196;
	wire new_net_5622;
	wire new_net_4576;
	wire new_net_7689;
	wire new_net_1797;
	wire _0702_;
	wire _0996_;
	wire _0198_;
	wire _1206_;
	wire new_net_1247;
	wire _0492_;
	wire new_net_3390;
	wire new_net_4351;
	wire new_net_4697;
	wire new_net_8144;
	wire new_net_7370;
	wire new_net_5968;
	wire new_net_4702;
	wire new_net_4597;
	wire new_net_1876;
	wire new_net_2988;
	wire new_net_412;
	wire new_net_745;
	wire new_net_3561;
	wire new_net_3604;
	wire new_net_3225;
	wire new_net_3249;
	wire new_net_4314;
	wire new_net_5265;
	wire new_net_6552;
	wire new_net_5655;
	wire new_net_8166;
	wire new_net_4832;
	wire new_net_1135;
	wire _0493_;
	wire _1207_;
	wire _0199_;
	wire new_net_344;
	wire new_net_1702;
	wire _0703_;
	wire new_net_3603;
	wire new_net_3208;
	wire _0997_;
	wire new_net_7303;
	wire new_net_6574;
	wire new_net_4854;
	wire new_net_8105;
	wire new_net_99;
	wire new_net_273;
	wire new_net_309;
	wire new_net_1283;
	wire new_net_3003;
	wire new_net_1860;
	wire new_net_1595;
	wire new_net_3295;
	wire new_net_4935;
	wire new_net_5163;
	wire _1208_;
	wire _0494_;
	wire _0200_;
	wire new_net_3671;
	wire _0704_;
	wire new_net_1248;
	wire new_net_2069;
	wire new_net_2206;
	wire _0998_;
	wire new_net_3940;
	wire new_net_4221;
	wire new_net_6685;
	wire new_net_746;
	wire new_net_1318;
	wire new_net_1666;
	wire new_net_3957;
	wire new_net_4281;
	wire new_net_4734;
	wire new_net_5243;
	wire new_net_5736;
	wire new_net_6107;
	wire new_net_3840;
	wire new_net_6250;
	wire new_net_5397;
	wire new_net_6095;
	wire new_net_1136;
	wire _0705_;
	wire _0999_;
	wire _1209_;
	wire _0495_;
	wire _0201_;
	wire new_net_345;
	wire new_net_3284;
	wire new_net_1487;
	wire new_net_3627;
	wire new_net_5242;
	wire new_net_8043;
	wire new_net_7680;
	wire new_net_6722;
	wire new_net_6896;
	wire new_net_1596;
	wire new_net_100;
	wire new_net_274;
	wire new_net_310;
	wire new_net_1284;
	wire new_net_4352;
	wire new_net_4698;
	wire new_net_5615;
	wire new_net_5986;
	wire new_net_6010;
	wire new_net_7184;
	wire new_net_7611;
	wire new_net_5264;
	wire new_net_6128;
	wire new_net_19;
	wire new_net_3226;
	wire _0706_;
	wire _1000_;
	wire _0496_;
	wire new_net_5;
	wire new_net_3250;
	wire new_net_1770;
	wire new_net_2989;
	wire _1210_;
	wire new_net_5721;
	wire new_net_6918;
	wire new_net_6467;
	wire new_net_6889;
	wire new_net_1319;
	wire new_net_2841;
	wire new_net_1667;
	wire new_net_1771;
	wire new_net_1703;
	wire new_net_3209;
	wire new_net_4021;
	wire new_net_4589;
	wire new_net_5494;
	wire new_net_7658;
	wire new_net_7717;
	wire new_net_7523;
	wire new_net_7884;
	wire new_net_7521;
	wire new_net_6364;
	wire new_net_1937;
	wire _0707_;
	wire _1001_;
	wire _0497_;
	wire _1211_;
	wire new_net_3296;
	wire _0203_;
	wire new_net_1488;
	wire new_net_4620;
	wire new_net_4642;
	wire new_net_5051;
	wire new_net_5634;
	wire new_net_5797;
	wire new_net_4367;
	wire new_net_101;
	wire new_net_275;
	wire new_net_311;
	wire new_net_3672;
	wire new_net_3941;
	wire new_net_4301;
	wire new_net_4316;
	wire new_net_4671;
	wire new_net_7156;
	wire new_net_7781;
	wire new_net_8073;
	wire _0178_;
	wire new_net_5897;
	wire new_net_4387;
	wire _0498_;
	wire _1212_;
	wire _0204_;
	wire _1002_;
	wire new_net_3268;
	wire _0708_;
	wire new_net_414;
	wire new_net_1250;
	wire new_net_1755;
	wire new_net_2207;
	wire new_net_7061;
	wire new_net_4882;
	wire new_net_6776;
	wire new_net_8095;
	wire new_net_5093;
	wire new_net_3628;
	wire new_net_346;
	wire new_net_1137;
	wire new_net_1668;
	wire new_net_1704;
	wire new_net_3285;
	wire new_net_4621;
	wire new_net_4964;
	wire new_net_6580;
	wire new_net_6258;
	wire new_net_7083;
	wire new_net_5233;
	wire new_net_7749;
	wire new_net_4240;
	wire new_net_8034;
	wire new_net_7081;
	wire _0499_;
	wire _1213_;
	wire _0205_;
	wire _1003_;
	wire new_net_1597;
	wire _0709_;
	wire new_net_1285;
	wire new_net_4152;
	wire new_net_4643;
	wire new_net_4699;
	wire new_net_4202;
	wire new_net_4926;
	wire new_net_5255;
	wire new_net_102;
	wire new_net_276;
	wire new_net_312;
	wire new_net_3227;
	wire new_net_3251;
	wire new_net_2990;
	wire new_net_3959;
	wire new_net_5267;
	wire new_net_5344;
	wire new_net_5394;
	wire new_net_5788;
	wire new_net_6418;
	wire new_net_4814;
	wire new_net_6708;
	wire new_net_4443;
	wire new_net_6502;
	wire new_net_748;
	wire new_net_1320;
	wire new_net_3210;
	wire _0710_;
	wire _1004_;
	wire _0500_;
	wire _1214_;
	wire new_net_1853;
	wire new_net_3743;
	wire new_net_1251;
	wire new_net_7998;
	wire new_net_5165;
	wire new_net_347;
	wire new_net_1138;
	wire new_net_2019;
	wire new_net_3391;
	wire new_net_1669;
	wire new_net_1489;
	wire new_net_3297;
	wire new_net_4937;
	wire new_net_4292;
	wire new_net_5047;
	wire new_net_6524;
	wire new_net_7357;
	wire new_net_5955;
	wire new_net_6283;
	wire new_net_7536;
	wire new_net_4071;
	wire new_net_7703;
	wire _0711_;
	wire _1005_;
	wire new_net_1598;
	wire _0501_;
	wire new_net_1913;
	wire new_net_2017;
	wire _1215_;
	wire new_net_3673;
	wire new_net_1781;
	wire _0207_;
	wire new_net_5180;
	wire new_net_7625;
	wire new_net_7623;
	wire new_net_8276;
	wire new_net_6917;
	wire new_net_6055;
	wire new_net_103;
	wire new_net_277;
	wire new_net_1993;
	wire new_net_3004;
	wire new_net_4245;
	wire new_net_4259;
	wire new_net_4283;
	wire new_net_4736;
	wire new_net_5245;
	wire new_net_5884;
	wire new_net_8086;
	wire new_net_5202;
	wire new_net_6561;
	wire new_net_7146;
	wire _0208_;
	wire new_net_2065;
	wire new_net_25;
	wire new_net_1321;
	wire new_net_2208;
	wire new_net_3605;
	wire _0502_;
	wire _1216_;
	wire _0712_;
	wire _1006_;
	wire new_net_5876;
	wire new_net_6827;
	wire new_net_7740;
	wire new_net_7246;
	wire new_net_6215;
	wire new_net_4598;
	wire new_net_7161;
	wire new_net_348;
	wire new_net_1139;
	wire new_net_1490;
	wire new_net_1939;
	wire new_net_3392;
	wire new_net_3763;
	wire new_net_1670;
	wire new_net_4153;
	wire new_net_4644;
	wire new_net_4700;
	wire new_net_6016;
	wire new_net_6672;
	wire new_net_6851;
	wire _0209_;
	wire new_net_1287;
	wire _0503_;
	wire _1217_;
	wire _1007_;
	wire new_net_3228;
	wire new_net_313;
	wire new_net_3252;
	wire new_net_3653;
	wire new_net_2991;
	wire new_net_6694;
	wire new_net_6866;
	wire new_net_5837;
	wire new_net_3878;
	wire new_net_6788;
	wire new_net_6;
	wire new_net_20;
	wire new_net_416;
	wire new_net_749;
	wire new_net_3211;
	wire new_net_3757;
	wire new_net_4023;
	wire new_net_4591;
	wire new_net_5496;
	wire new_net_7660;
	wire new_net_7984;
	wire new_net_7500;
	wire new_net_7331;
	wire new_net_4010;
	wire new_net_5935;
	wire new_net_3298;
	wire new_net_1253;
	wire _0210_;
	wire _0714_;
	wire _1008_;
	wire _0504_;
	wire new_net_2842;
	wire new_net_1706;
	wire _1218_;
	wire new_net_3934;
	wire new_net_4985;
	wire new_net_3788;
	wire new_net_349;
	wire new_net_1140;
	wire new_net_1599;
	wire new_net_1671;
	wire new_net_3674;
	wire new_net_3654;
	wire new_net_3376;
	wire new_net_3943;
	wire new_net_5863;
	wire new_net_7158;
	wire new_net_4396;
	wire new_net_7115;
	wire new_net_6992;
	wire new_net_7287;
	wire new_net_5026;
	wire _0715_;
	wire _0211_;
	wire _1219_;
	wire new_net_3572;
	wire _1009_;
	wire _0505_;
	wire new_net_104;
	wire new_net_314;
	wire new_net_2967;
	wire new_net_3269;
	wire new_net_7132;
	wire new_net_7016;
	wire new_net_1805;
	wire new_net_417;
	wire new_net_750;
	wire new_net_3630;
	wire new_net_1322;
	wire new_net_3606;
	wire new_net_1798;
	wire new_net_3287;
	wire new_net_4247;
	wire new_net_4623;
	wire new_net_3377;
	wire _0716_;
	wire _0212_;
	wire _0506_;
	wire _1220_;
	wire new_net_1491;
	wire new_net_2209;
	wire _1010_;
	wire new_net_1748;
	wire new_net_2843;
	wire new_net_6297;
	wire new_net_7871;
	wire new_net_7953;
	wire new_net_5694;
	wire new_net_2091;
	wire new_net_1141;
	wire new_net_1288;
	wire new_net_1600;
	wire new_net_1672;
	wire new_net_3229;
	wire new_net_2968;
	wire new_net_5269;
	wire new_net_5396;
	wire new_net_6133;
	wire new_net_6029;
	wire new_net_5906;
	wire new_net_4612;
	wire new_net_7810;
	wire new_net_4321;
	wire _1221_;
	wire _0717_;
	wire _0213_;
	wire _1011_;
	wire _0507_;
	wire new_net_105;
	wire new_net_315;
	wire new_net_4024;
	wire new_net_5497;
	wire new_net_7319;
	wire new_net_4332;
	wire new_net_5515;
	wire new_net_6334;
	wire new_net_1707;
	wire new_net_1254;
	wire new_net_3299;
	wire new_net_418;
	wire new_net_751;
	wire new_net_1323;
	wire new_net_2027;
	wire new_net_4939;
	wire new_net_5167;
	wire new_net_5373;
	wire new_net_7462;
	wire new_net_7341;
	wire new_net_7334;
	wire new_net_6216;
	wire new_net_7763;
	wire new_net_7269;
	wire new_net_350;
	wire _1222_;
	wire new_net_3675;
	wire _0718_;
	wire _1012_;
	wire _0214_;
	wire new_net_1492;
	wire _0508_;
	wire new_net_3944;
	wire new_net_3960;
	wire new_net_7567;
	wire new_net_7769;
	wire new_net_1142;
	wire new_net_1289;
	wire new_net_1601;
	wire new_net_1673;
	wire new_net_4261;
	wire new_net_4285;
	wire new_net_4738;
	wire new_net_5886;
	wire new_net_6111;
	wire new_net_6858;
	wire new_net_8237;
	wire new_net_4404;
	wire new_net_7201;
	wire new_net_7791;
	wire new_net_7123;
	wire new_net_7789;
	wire new_net_5152;
	wire _1223_;
	wire new_net_3005;
	wire _0215_;
	wire _0719_;
	wire new_net_3607;
	wire new_net_3631;
	wire new_net_3562;
	wire _1013_;
	wire _0509_;
	wire new_net_106;
	wire new_net_6804;
	wire new_net_7427;
	wire new_net_5456;
	wire new_net_6116;
	wire new_net_5623;
	wire new_net_4766;
	wire new_net_1708;
	wire new_net_419;
	wire new_net_752;
	wire new_net_1255;
	wire new_net_1728;
	wire new_net_3378;
	wire new_net_2844;
	wire new_net_3394;
	wire new_net_4337;
	wire new_net_4646;
	wire new_net_7857;
	wire new_net_6538;
	wire new_net_8145;
	wire new_net_4703;
	wire new_net_2969;
	wire new_net_351;
	wire new_net_1849;
	wire _0510_;
	wire _1224_;
	wire _0216_;
	wire _0720_;
	wire new_net_2210;
	wire _1014_;
	wire new_net_3230;
	wire new_net_8169;
	wire new_net_5366;
	wire new_net_6553;
	wire new_net_8167;
	wire new_net_4833;
	wire new_net_7294;
	wire new_net_3563;
	wire new_net_1143;
	wire new_net_1674;
	wire new_net_3758;
	wire new_net_4025;
	wire new_net_4154;
	wire new_net_4960;
	wire new_net_5498;
	wire new_net_7159;
	wire new_net_7662;
	wire new_net_6575;
	wire new_net_4855;
	wire _0511_;
	wire _1225_;
	wire _0217_;
	wire _0721_;
	wire new_net_3300;
	wire new_net_1324;
	wire _1015_;
	wire new_net_4940;
	wire new_net_5168;
	wire new_net_5374;
	wire new_net_7255;
	wire new_net_753;
	wire new_net_1256;
	wire new_net_3676;
	wire new_net_1493;
	wire new_net_3945;
	wire new_net_4162;
	wire new_net_4319;
	wire new_net_5865;
	wire new_net_7785;
	wire new_net_7907;
	wire new_net_4058;
	wire new_net_6686;
	wire new_net_7809;
	wire new_net_1602;
	wire _0512_;
	wire _0722_;
	wire _1016_;
	wire _0218_;
	wire _1226_;
	wire new_net_3006;
	wire new_net_1290;
	wire new_net_4262;
	wire new_net_4286;
	wire new_net_6251;
	wire new_net_6878;
	wire new_net_1675;
	wire new_net_107;
	wire new_net_317;
	wire new_net_1144;
	wire new_net_3608;
	wire new_net_3632;
	wire new_net_4592;
	wire new_net_4625;
	wire new_net_6096;
	wire new_net_6584;
	wire new_net_6725;
	wire new_net_8044;
	wire new_net_7681;
	wire new_net_3379;
	wire _0513_;
	wire new_net_3395;
	wire _0723_;
	wire _1017_;
	wire _1227_;
	wire new_net_1709;
	wire new_net_420;
	wire _0219_;
	wire new_net_1325;
	wire new_net_4651;
	wire new_net_7187;
	wire new_net_4649;
	wire new_net_7185;
	wire new_net_6129;
	wire new_net_6747;
	wire new_net_3231;
	wire new_net_2970;
	wire new_net_3253;
	wire new_net_352;
	wire new_net_754;
	wire new_net_1257;
	wire new_net_1494;
	wire new_net_5247;
	wire new_net_5271;
	wire new_net_5398;
	wire new_net_6745;
	wire new_net_6919;
	wire new_net_6468;
	wire new_net_4711;
	wire _1018_;
	wire new_net_1603;
	wire _0514_;
	wire new_net_1747;
	wire new_net_3254;
	wire _0220_;
	wire _1228_;
	wire _0724_;
	wire new_net_1291;
	wire new_net_2211;
	wire new_net_6890;
	wire new_net_7836;
	wire new_net_7524;
	wire new_net_7885;
	wire new_net_7441;
	wire new_net_4846;
	wire new_net_4577;
	wire new_net_108;
	wire new_net_1779;
	wire new_net_318;
	wire new_net_1145;
	wire new_net_1676;
	wire new_net_3301;
	wire new_net_4593;
	wire new_net_4941;
	wire new_net_5169;
	wire new_net_5741;
	wire new_net_5798;
	wire new_net_5759;
	wire new_net_4373;
	wire new_net_26;
	wire _0515_;
	wire _0725_;
	wire _1019_;
	wire _0221_;
	wire _1229_;
	wire new_net_3677;
	wire new_net_1710;
	wire new_net_3946;
	wire new_net_3812;
	wire new_net_353;
	wire new_net_755;
	wire new_net_1861;
	wire new_net_1495;
	wire new_net_4263;
	wire new_net_4287;
	wire new_net_4320;
	wire new_net_4355;
	wire new_net_4740;
	wire new_net_5888;
	wire new_net_6237;
	wire new_net_4099;
	wire new_net_6777;
	wire new_net_8096;
	wire new_net_7137;
	wire new_net_5389;
	wire _1020_;
	wire new_net_1604;
	wire new_net_1862;
	wire _0516_;
	wire new_net_3633;
	wire new_net_1866;
	wire _1230_;
	wire _0726_;
	wire new_net_3609;
	wire _0222_;
	wire new_net_6087;
	wire new_net_7084;
	wire new_net_7750;
	wire new_net_8035;
	wire new_net_7082;
	wire new_net_1272;
	wire new_net_5111;
	wire new_net_3380;
	wire new_net_109;
	wire new_net_283;
	wire new_net_1146;
	wire new_net_1326;
	wire new_net_3396;
	wire new_net_1677;
	wire _1194_;
	wire new_net_4339;
	wire new_net_4648;
	wire new_net_8258;
	wire new_net_5256;
	wire new_net_3232;
	wire _0727_;
	wire _1021_;
	wire _0517_;
	wire new_net_2971;
	wire new_net_1846;
	wire _1231_;
	wire new_net_422;
	wire new_net_1258;
	wire _0223_;
	wire new_net_6709;
	wire new_net_4630;
	wire new_net_3212;
	wire new_net_2095;
	wire new_net_756;
	wire new_net_1496;
	wire new_net_4027;
	wire new_net_4248;
	wire new_net_5500;
	wire new_net_7664;
	wire new_net_4628;
	wire new_net_7707;
	wire new_net_5166;
	wire new_net_2212;
	wire new_net_3215;
	wire new_net_1605;
	wire _0728_;
	wire _1022_;
	wire _0518_;
	wire new_net_1799;
	wire _1232_;
	wire new_net_3302;
	wire _0224_;
	wire new_net_6525;
	wire new_net_5048;
	wire new_net_7358;
	wire new_net_110;
	wire new_net_284;
	wire new_net_1147;
	wire new_net_1327;
	wire new_net_1711;
	wire new_net_3678;
	wire new_net_2071;
	wire new_net_3947;
	wire new_net_3962;
	wire new_net_5867;
	wire new_net_8065;
	wire new_net_5181;
	wire new_net_7626;
	wire new_net_8277;
	wire new_net_4948;
	wire new_net_5889;
	wire _0519_;
	wire _0729_;
	wire _1023_;
	wire _0225_;
	wire new_net_2845;
	wire new_net_3255;
	wire new_net_354;
	wire _0916_;
	wire _1233_;
	wire new_net_423;
	wire new_net_4874;
	wire new_net_8087;
	wire new_net_6942;
	wire new_net_4424;
	wire new_net_5375;
	wire new_net_6562;
	wire new_net_7147;
	wire new_net_1497;
	wire new_net_2038;
	wire new_net_3610;
	wire new_net_3213;
	wire new_net_3634;
	wire new_net_757;
	wire new_net_3759;
	wire new_net_3007;
	wire new_net_4249;
	wire new_net_4627;
	wire new_net_6658;
	wire new_net_4468;
	wire new_net_6828;
	wire new_net_7247;
	wire new_net_5682;
	wire new_net_6223;
	wire _0520_;
	wire _0226_;
	wire _1024_;
	wire new_net_1606;
	wire new_net_3381;
	wire new_net_320;
	wire new_net_1749;
	wire new_net_3397;
	wire new_net_1678;
	wire _1234_;
	wire new_net_4368;
	wire new_net_4599;
	wire new_net_7162;
	wire new_net_6017;
	wire new_net_6673;
	wire new_net_6852;
	wire new_net_6845;
	wire new_net_6434;
	wire new_net_3573;
	wire new_net_111;
	wire new_net_285;
	wire new_net_1328;
	wire new_net_3233;
	wire new_net_2846;
	wire new_net_2972;
	wire new_net_1712;
	wire new_net_4156;
	wire new_net_4305;
	wire new_net_5704;
	wire new_net_4806;
	wire new_net_6874;
	wire new_net_6867;
	wire new_net_424;
	wire _0227_;
	wire _0731_;
	wire _1025_;
	wire _0521_;
	wire new_net_355;
	wire _1235_;
	wire new_net_4028;
	wire new_net_4659;
	wire new_net_5501;
	wire new_net_6789;
	wire new_net_4039;
	wire new_net_7985;
	wire new_net_4565;
	wire new_net_3303;
	wire new_net_1498;
	wire new_net_1894;
	wire new_net_758;
	wire new_net_1294;
	wire new_net_2092;
	wire new_net_4943;
	wire new_net_4958;
	wire new_net_5171;
	wire new_net_5743;
	wire new_net_5936;
	wire new_net_6516;
	wire new_net_3574;
	wire _0228_;
	wire new_net_27;
	wire new_net_2213;
	wire _0732_;
	wire _1026_;
	wire new_net_13;
	wire new_net_1607;
	wire _0522_;
	wire new_net_321;
	wire new_net_4934;
	wire new_net_7290;
	wire new_net_7661;
	wire new_net_6993;
	wire new_net_7288;
	wire new_net_1844;
	wire new_net_112;
	wire new_net_286;
	wire new_net_1260;
	wire new_net_1713;
	wire new_net_4265;
	wire new_net_4289;
	wire new_net_4742;
	wire new_net_5890;
	wire new_net_6115;
	wire new_net_7634;
	wire new_net_4132;
	wire new_net_7216;
	wire new_net_7133;
	wire new_net_5656;
	wire _1237_;
	wire _0229_;
	wire new_net_3611;
	wire _0523_;
	wire _0733_;
	wire _1027_;
	wire new_net_3214;
	wire new_net_3635;
	wire new_net_3270;
	wire new_net_4306;
	wire new_net_5868;
	wire new_net_7238;
	wire new_net_1499;
	wire new_net_759;
	wire new_net_1295;
	wire new_net_1892;
	wire new_net_3382;
	wire new_net_3398;
	wire new_net_1847;
	wire new_net_4362;
	wire new_net_4650;
	wire new_net_4706;
	wire new_net_6298;
	wire new_net_7383;
	wire new_net_4239;
	wire _1238_;
	wire new_net_3008;
	wire new_net_3564;
	wire new_net_1329;
	wire _0524_;
	wire _0734_;
	wire _1028_;
	wire _0230_;
	wire new_net_1608;
	wire new_net_2094;
	wire new_net_6030;
	wire new_net_6769;
	wire new_net_7811;
	wire new_net_1714;
	wire new_net_3565;
	wire new_net_1261;
	wire new_net_1901;
	wire new_net_113;
	wire new_net_356;
	wire new_net_425;
	wire new_net_5502;
	wire new_net_7666;
	wire new_net_8008;
	wire new_net_5516;
	wire new_net_6335;
	wire _1239_;
	wire new_net_3304;
	wire _0231_;
	wire _0735_;
	wire _1029_;
	wire _0525_;
	wire new_net_4944;
	wire new_net_4957;
	wire new_net_5744;
	wire new_net_6340;
	wire new_net_6585;
	wire new_net_7465;
	wire new_net_8116;
	wire new_net_4270;
	wire new_net_7463;
	wire new_net_4785;
	wire new_net_7335;
	wire new_net_3973;
	wire new_net_2993;
	wire new_net_3288;
	wire new_net_3680;
	wire new_net_3575;
	wire new_net_1500;
	wire new_net_3949;
	wire new_net_3964;
	wire new_net_4595;
	wire new_net_5869;
	wire new_net_7270;
	wire new_net_6446;
	wire new_net_7770;
	wire new_net_1238;
	wire new_net_4588;
	wire new_net_6495;
	wire new_net_7413;
	wire new_net_8238;
	wire new_net_4739;
	wire new_net_4123;
	wire new_net_7202;
	wire new_net_3578;
	wire new_net_7792;
	wire new_net_7124;
	wire new_net_2340;
	wire new_net_3029;
	wire _0274_;
	wire _0778_;
	wire new_net_2920;
	wire new_net_2277;
	wire new_net_3089;
	wire new_net_4035;
	wire new_net_4439;
	wire new_net_4755;
	wire new_net_7428;
	wire new_net_7647;
	wire new_net_7691;
	wire new_net_6284;
	wire new_net_1890;
	wire new_net_3409;
	wire new_net_1448;
	wire new_net_60;
	wire new_net_4055;
	wire new_net_5183;
	wire new_net_5286;
	wire new_net_6150;
	wire new_net_6478;
	wire new_net_6600;
	wire new_net_6746;
	wire new_net_6539;
	wire new_net_7858;
	wire new_net_5970;
	wire new_net_4704;
	wire new_net_3443;
	wire _0275_;
	wire _0779_;
	wire new_net_3481;
	wire new_net_4571;
	wire new_net_5308;
	wire new_net_7453;
	wire new_net_8074;
	wire new_net_8170;
	wire new_net_8168;
	wire new_net_4834;
	wire new_net_6645;
	wire new_net_7969;
	wire new_net_2853;
	wire new_net_12;
	wire new_net_1519;
	wire new_net_1627;
	wire new_net_2668;
	wire new_net_5536;
	wire new_net_5560;
	wire new_net_6953;
	wire new_net_7221;
	wire new_net_4856;
	wire new_net_8107;
	wire new_net_2309;
	wire new_net_3110;
	wire new_net_1965;
	wire new_net_2120;
	wire new_net_2870;
	wire _0276_;
	wire _0780_;
	wire new_net_2487;
	wire new_net_2905;
	wire new_net_2795;
	wire new_net_7256;
	wire new_net_4090;
	wire new_net_1449;
	wire new_net_3803;
	wire new_net_4400;
	wire new_net_4419;
	wire new_net_4715;
	wire new_net_4979;
	wire new_net_6231;
	wire new_net_6353;
	wire new_net_6724;
	wire new_net_7095;
	wire new_net_3640;
	wire new_net_167;
	wire new_net_374;
	wire _0277_;
	wire _0781_;
	wire new_net_3693;
	wire new_net_3462;
	wire new_net_3588;
	wire new_net_3977;
	wire new_net_4178;
	wire new_net_4398;
	wire new_net_6252;
	wire new_net_4379;
	wire new_net_5399;
	wire new_net_3090;
	wire new_net_23;
	wire new_net_1520;
	wire new_net_3030;
	wire new_net_2921;
	wire new_net_3051;
	wire new_net_4036;
	wire new_net_4075;
	wire new_net_4440;
	wire new_net_4756;
	wire new_net_5244;
	wire new_net_8045;
	wire new_net_7682;
	wire new_net_61;
	wire new_net_2278;
	wire new_net_2341;
	wire _0278_;
	wire _0782_;
	wire new_net_3315;
	wire new_net_4056;
	wire new_net_5184;
	wire new_net_5287;
	wire new_net_6151;
	wire new_net_7186;
	wire new_net_5956;
	wire new_net_413;
	wire new_net_5266;
	wire new_net_6130;
	wire new_net_3482;
	wire new_net_1450;
	wire new_net_3329;
	wire new_net_4364;
	wire new_net_4572;
	wire new_net_4971;
	wire new_net_5309;
	wire new_net_6994;
	wire new_net_5723;
	wire new_net_6920;
	wire new_net_6469;
	wire new_net_6058;
	wire new_net_6891;
	wire new_net_3641;
	wire new_net_1628;
	wire new_net_168;
	wire new_net_375;
	wire _0783_;
	wire _0279_;
	wire new_net_2617;
	wire new_net_2669;
	wire new_net_5537;
	wire new_net_5561;
	wire new_net_7721;
	wire new_net_7719;
	wire new_net_7888;
	wire new_net_4682;
	wire new_net_7886;
	wire new_net_4583;
	wire new_net_2570;
	wire new_net_3111;
	wire new_net_3545;
	wire new_net_1521;
	wire new_net_2056;
	wire new_net_3339;
	wire new_net_2796;
	wire new_net_2871;
	wire new_net_2906;
	wire new_net_4383;
	wire new_net_5053;
	wire new_net_5716;
	wire new_net_6624;
	wire new_net_5760;
	wire new_net_2247;
	wire new_net_62;
	wire new_net_2310;
	wire _0280_;
	wire _0784_;
	wire new_net_2121;
	wire new_net_3014;
	wire new_net_3316;
	wire new_net_3804;
	wire new_net_4211;
	wire new_net_5899;
	wire new_net_3410;
	wire new_net_1451;
	wire new_net_3694;
	wire new_net_3463;
	wire new_net_3589;
	wire new_net_3978;
	wire new_net_4179;
	wire new_net_5756;
	wire new_net_6601;
	wire new_net_7063;
	wire new_net_6778;
	wire new_net_8097;
	wire new_net_5137;
	wire new_net_2922;
	wire new_net_3196;
	wire new_net_3091;
	wire new_net_1629;
	wire new_net_3546;
	wire _0281_;
	wire _0785_;
	wire new_net_169;
	wire new_net_2618;
	wire new_net_3031;
	wire new_net_7085;
	wire new_net_8036;
	wire new_net_1522;
	wire new_net_2854;
	wire new_net_2519;
	wire new_net_4057;
	wire new_net_5185;
	wire new_net_5288;
	wire new_net_6152;
	wire new_net_6255;
	wire new_net_6480;
	wire new_net_6748;
	wire new_net_8259;
	wire new_net_4928;
	wire new_net_3483;
	wire new_net_63;
	wire new_net_2279;
	wire new_net_2342;
	wire _0282_;
	wire _0786_;
	wire new_net_2039;
	wire new_net_5310;
	wire new_net_6995;
	wire new_net_7455;
	wire new_net_5346;
	wire new_net_2216;
	wire new_net_4816;
	wire new_net_6710;
	wire new_net_4448;
	wire new_net_4631;
	wire new_net_6504;
	wire new_net_2670;
	wire new_net_3642;
	wire new_net_376;
	wire new_net_3426;
	wire new_net_1452;
	wire new_net_5538;
	wire new_net_5562;
	wire new_net_6955;
	wire new_net_7096;
	wire new_net_7223;
	wire new_net_2489;
	wire new_net_2907;
	wire new_net_1750;
	wire new_net_2797;
	wire new_net_2571;
	wire new_net_1630;
	wire _0787_;
	wire _0283_;
	wire new_net_3340;
	wire new_net_3197;
	wire new_net_6526;
	wire new_net_4294;
	wire new_net_7359;
	wire new_net_7538;
	wire new_net_3317;
	wire new_net_1523;
	wire new_net_1966;
	wire new_net_3444;
	wire new_net_3805;
	wire new_net_4421;
	wire new_net_6233;
	wire new_net_6355;
	wire new_net_5182;
	wire new_net_6726;
	wire new_net_7627;
	wire new_net_8278;
	wire new_net_3464;
	wire new_net_3590;
	wire new_net_2248;
	wire new_net_64;
	wire new_net_2311;
	wire _0788_;
	wire _0284_;
	wire new_net_2122;
	wire new_net_3427;
	wire new_net_3695;
	wire new_net_8088;
	wire new_net_5204;
	wire new_net_6943;
	wire new_net_5376;
	wire new_net_1769;
	wire new_net_3594;
	wire new_net_4613;
	wire new_net_6563;
	wire new_net_7148;
	wire new_net_3032;
	wire new_net_2923;
	wire new_net_3092;
	wire new_net_377;
	wire new_net_4038;
	wire new_net_4077;
	wire new_net_4442;
	wire new_net_4717;
	wire new_net_4758;
	wire new_net_4857;
	wire new_net_5878;
	wire new_net_7742;
	wire new_net_6045;
	wire new_net_7248;
	wire new_net_5683;
	wire new_net_4369;
	wire new_net_6217;
	wire _0285_;
	wire _0789_;
	wire new_net_3411;
	wire new_net_3781;
	wire new_net_5186;
	wire new_net_5289;
	wire new_net_6153;
	wire new_net_6256;
	wire new_net_6481;
	wire new_net_6749;
	wire new_net_6308;
	wire new_net_1879;
	wire _0186_;
	wire new_net_6853;
	wire new_net_6435;
	wire new_net_3445;
	wire new_net_3484;
	wire new_net_1524;
	wire new_net_5125;
	wire new_net_5311;
	wire new_net_6996;
	wire new_net_7456;
	wire new_net_6696;
	wire new_net_6875;
	wire new_net_7821;
	wire new_net_5839;
	wire new_net_3880;
	wire new_net_1453;
	wire new_net_1855;
	wire _0790_;
	wire new_net_2671;
	wire new_net_2280;
	wire new_net_3643;
	wire _0286_;
	wire new_net_2343;
	wire new_net_2855;
	wire new_net_4402;
	wire new_net_7986;
	wire new_net_4405;
	wire new_net_7502;
	wire new_net_4907;
	wire new_net_4490;
	wire new_net_3938;
	wire new_net_2908;
	wire new_net_2798;
	wire new_net_3052;
	wire new_net_3198;
	wire new_net_3341;
	wire new_net_2552;
	wire new_net_2706;
	wire new_net_171;
	wire new_net_378;
	wire new_net_1631;
	wire new_net_3936;
	wire new_net_7704;
	wire new_net_4988;
	wire new_net_3318;
	wire new_net_2572;
	wire _0791_;
	wire _0287_;
	wire new_net_3782;
	wire new_net_3806;
	wire new_net_4212;
	wire new_net_4422;
	wire new_net_5430;
	wire new_net_6234;
	wire new_net_7289;
	wire new_net_3696;
	wire new_net_3465;
	wire new_net_65;
	wire new_net_1525;
	wire new_net_1735;
	wire new_net_3980;
	wire new_net_4181;
	wire new_net_5758;
	wire new_net_6603;
	wire new_net_4133;
	wire new_net_7217;
	wire new_net_2123;
	wire new_net_1454;
	wire new_net_2518;
	wire new_net_3033;
	wire new_net_2924;
	wire new_net_3053;
	wire new_net_2249;
	wire new_net_2553;
	wire _0792_;
	wire _0288_;
	wire new_net_2699;
	wire new_net_7239;
	wire new_net_172;
	wire new_net_379;
	wire new_net_2707;
	wire new_net_1632;
	wire new_net_3112;
	wire new_net_5187;
	wire new_net_5290;
	wire new_net_6154;
	wire new_net_6257;
	wire new_net_6377;
	wire new_net_4669;
	wire new_net_7873;
	wire new_net_7384;
	wire new_net_3015;
	wire new_net_3446;
	wire new_net_1753;
	wire new_net_3485;
	wire _0793_;
	wire _0289_;
	wire new_net_5312;
	wire new_net_6997;
	wire new_net_7457;
	wire new_net_6399;
	wire new_net_6031;
	wire new_net_7812;
	wire _0676_;
	wire new_net_2619;
	wire new_net_3018;
	wire new_net_66;
	wire new_net_2672;
	wire new_net_1526;
	wire new_net_2142;
	wire new_net_4573;
	wire new_net_5540;
	wire new_net_5564;
	wire new_net_6957;
	wire new_net_7321;
	wire new_net_5517;
	wire new_net_6336;
	wire new_net_6588;
	wire new_net_6586;
	wire new_net_2344;
	wire new_net_2909;
	wire new_net_2874;
	wire new_net_3428;
	wire new_net_1455;
	wire new_net_2491;
	wire new_net_2799;
	wire new_net_3342;
	wire _0794_;
	wire _0290_;
	wire new_net_7464;
	wire new_net_8117;
	wire new_net_2173;
	wire new_net_7343;
	wire _0187_;
	wire new_net_5539;
	wire new_net_7765;
	wire new_net_1873;
	wire new_net_3319;
	wire new_net_380;
	wire new_net_3113;
	wire new_net_3783;
	wire new_net_3807;
	wire new_net_4060;
	wire new_net_4386;
	wire new_net_4403;
	wire new_net_4423;
	wire new_net_7271;
	wire new_net_7771;
	wire new_net_3412;
	wire new_net_2620;
	wire new_net_3466;
	wire new_net_3016;
	wire new_net_3697;
	wire _0795_;
	wire _0291_;
	wire new_net_3981;
	wire new_net_4182;
	wire new_net_4213;
	wire new_net_7414;
	wire new_net_5438;
	wire new_net_8239;
	wire new_net_7203;
	wire new_net_7793;
	wire new_net_7125;
	wire new_net_3034;
	wire new_net_1527;
	wire new_net_2925;
	wire new_net_67;
	wire new_net_2554;
	wire new_net_3094;
	wire new_net_4040;
	wire new_net_4079;
	wire new_net_4444;
	wire new_net_4760;
	wire new_net_6118;
	wire new_net_1652;
	wire new_net_1633;
	wire new_net_2313;
	wire new_net_173;
	wire new_net_1986;
	wire new_net_2124;
	wire _0796_;
	wire _0292_;
	wire new_net_2250;
	wire new_net_2708;
	wire new_net_4059;
	wire new_net_6285;
	wire new_net_7859;
	wire new_net_7910;
	wire new_net_5971;
	wire new_net_4705;
	wire new_net_3413;
	wire new_net_3447;
	wire new_net_3486;
	wire new_net_381;
	wire new_net_5313;
	wire new_net_6998;
	wire new_net_7077;
	wire new_net_7458;
	wire new_net_2357;
	wire new_net_8075;
	wire new_net_5733;
	wire new_net_6930;
	wire new_net_8171;
	wire new_net_6479;
	wire new_net_4835;
	wire _0366_;
	wire _0797_;
	wire _0293_;
	wire new_net_2673;
	wire new_net_5541;
	wire new_net_5565;
	wire new_net_7099;
	wire new_net_7970;
	wire new_net_6160;
	wire new_net_6248;
	wire new_net_4093;
	wire new_net_2875;
	wire new_net_2517;
	wire new_net_2910;
	wire new_net_1456;
	wire new_net_1528;
	wire new_net_2800;
	wire new_net_3343;
	wire new_net_4837;
	wire new_net_5211;
	wire new_net_5417;
	wire new_net_8108;
	wire new_net_4673;
	wire new_net_7751;
	wire new_net_7257;
	wire new_net_2282;
	wire new_net_1634;
	wire new_net_2345;
	wire new_net_174;
	wire new_net_3320;
	wire _0798_;
	wire _0294_;
	wire new_net_3114;
	wire new_net_3784;
	wire new_net_3808;
	wire new_net_3591;
	wire new_net_3547;
	wire new_net_3467;
	wire new_net_2621;
	wire new_net_3429;
	wire new_net_3017;
	wire new_net_3698;
	wire new_net_382;
	wire new_net_3982;
	wire new_net_4183;
	wire new_net_8225;
	wire new_net_4334;
	wire new_net_6422;
	wire new_net_6420;
	wire new_net_68;
	wire new_net_3095;
	wire new_net_3644;
	wire new_net_2856;
	wire new_net_3035;
	wire _0295_;
	wire _0799_;
	wire new_net_1751;
	wire new_net_2926;
	wire new_net_2555;
	wire new_net_6727;
	wire new_net_8046;
	wire new_net_3177;
	wire new_net_1972;
	wire new_net_1457;
	wire new_net_1529;
	wire new_net_3199;
	wire new_net_5292;
	wire new_net_6156;
	wire new_net_6259;
	wire new_net_6484;
	wire new_net_6752;
	wire new_net_7226;
	wire new_net_7683;
	wire new_net_7189;
	wire new_net_2192;
	wire new_net_2251;
	wire new_net_1635;
	wire new_net_2314;
	wire new_net_3414;
	wire new_net_175;
	wire new_net_2125;
	wire new_net_3448;
	wire _0296_;
	wire _0800_;
	wire new_net_3487;
	wire new_net_5479;
	wire new_net_6921;
	wire new_net_6470;
	wire new_net_7005;
	wire _0003_;
	wire new_net_2573;
	wire new_net_3548;
	wire new_net_383;
	wire new_net_3592;
	wire new_net_2674;
	wire new_net_5542;
	wire new_net_7100;
	wire new_net_7845;
	wire new_net_7838;
	wire new_net_170;
	wire new_net_1365;
	wire new_net_7889;
	wire new_net_7526;
	wire new_net_7887;
	wire new_net_69;
	wire new_net_2857;
	wire new_net_2876;
	wire _0297_;
	wire _0801_;
	wire new_net_2493;
	wire new_net_2911;
	wire new_net_2801;
	wire new_net_3200;
	wire new_net_3344;
	wire new_net_4513;
	wire new_net_4848;
	wire new_net_4353;
	wire new_net_5761;
	wire new_net_3115;
	wire new_net_1530;
	wire new_net_1906;
	wire new_net_3321;
	wire new_net_3785;
	wire new_net_3809;
	wire new_net_4388;
	wire new_net_4425;
	wire new_net_4445;
	wire new_net_6224;
	wire new_net_6018;
	wire new_net_6674;
	wire _0058_;
	wire new_net_5900;
	wire new_net_3286;
	wire new_net_2283;
	wire new_net_1636;
	wire new_net_2346;
	wire new_net_176;
	wire new_net_3430;
	wire new_net_3699;
	wire _0298_;
	wire _0802_;
	wire new_net_3468;
	wire new_net_3983;
	wire new_net_6239;
	wire new_net_4101;
	wire new_net_7064;
	wire new_net_6779;
	wire new_net_8098;
	wire new_net_1387;
	wire new_net_2927;
	wire new_net_2556;
	wire new_net_2574;
	wire new_net_3096;
	wire new_net_384;
	wire new_net_3036;
	wire new_net_4081;
	wire new_net_4590;
	wire new_net_5520;
	wire new_net_6980;
	wire new_net_4310;
	wire new_net_7086;
	wire new_net_5236;
	wire new_net_8037;
	wire new_net_1756;
	wire _0299_;
	wire _0803_;
	wire new_net_1458;
	wire new_net_4446;
	wire new_net_5113;
	wire new_net_5293;
	wire new_net_5566;
	wire new_net_6260;
	wire new_net_6485;
	wire new_net_8260;
	wire new_net_3488;
	wire new_net_1531;
	wire _0678_;
	wire new_net_3449;
	wire new_net_4214;
	wire new_net_4575;
	wire new_net_4718;
	wire new_net_5258;
	wire new_net_5315;
	wire new_net_7000;
	wire new_net_2516;
	wire new_net_2675;
	wire new_net_2252;
	wire new_net_1637;
	wire new_net_2315;
	wire new_net_3549;
	wire new_net_177;
	wire new_net_2126;
	wire _0804_;
	wire _0300_;
	wire new_net_3615;
	wire new_net_4632;
	wire new_net_2802;
	wire new_net_3054;
	wire new_net_3201;
	wire new_net_3345;
	wire new_net_2709;
	wire new_net_2912;
	wire new_net_2877;
	wire new_net_70;
	wire new_net_385;
	wire new_net_4166;
	wire new_net_2803;
	wire new_net_3322;
	wire _0301_;
	wire _0805_;
	wire new_net_1459;
	wire new_net_3786;
	wire new_net_3810;
	wire new_net_4426;
	wire new_net_5563;
	wire new_net_6238;
	wire new_net_6360;
	wire new_net_2155;
	wire new_net_7628;
	wire new_net_8279;
	wire new_net_4950;
	wire new_net_3469;
	wire new_net_1903;
	wire new_net_1977;
	wire new_net_3431;
	wire new_net_3700;
	wire new_net_3984;
	wire new_net_4185;
	wire new_net_5762;
	wire new_net_6157;
	wire new_net_6607;
	wire new_net_6944;
	wire new_net_5377;
	wire new_net_6564;
	wire new_net_3037;
	wire new_net_2928;
	wire new_net_2557;
	wire new_net_2284;
	wire new_net_2575;
	wire new_net_3097;
	wire new_net_1638;
	wire new_net_2347;
	wire _0302_;
	wire _0806_;
	wire new_net_6660;
	wire new_net_6046;
	wire new_net_2710;
	wire new_net_71;
	wire new_net_386;
	wire new_net_4447;
	wire new_net_5294;
	wire new_net_5567;
	wire new_net_5684;
	wire new_net_6218;
	wire new_net_6261;
	wire new_net_6486;
	wire new_net_6309;
	wire _0059_;
	wire new_net_6854;
	wire new_net_6847;
	wire new_net_6436;
	wire new_net_1877;
	wire new_net_3450;
	wire new_net_1532;
	wire new_net_3489;
	wire _0303_;
	wire _0807_;
	wire new_net_5316;
	wire new_net_7001;
	wire new_net_7461;
	wire new_net_5706;
	wire new_net_2405;
	wire new_net_6876;
	wire new_net_7822;
	wire new_net_2676;
	wire new_net_1838;
	wire new_net_178;
	wire new_net_3550;
	wire new_net_4861;
	wire new_net_5544;
	wire new_net_6869;
	wire new_net_7102;
	wire new_net_4041;
	wire new_net_7987;
	wire new_net_4341;
	wire new_net_7503;
	wire new_net_223;
	wire new_net_2467;
	wire new_net_1973;
	wire new_net_2127;
	wire new_net_2878;
	wire new_net_1874;
	wire new_net_2495;
	wire new_net_3202;
	wire new_net_2253;
	wire new_net_2316;
	wire _0808_;
	wire _0304_;
	wire new_net_6518;
	wire new_net_7648;
	wire new_net_4684;
	wire new_net_2622;
	wire new_net_1460;
	wire new_net_3323;
	wire new_net_2804;
	wire new_net_3019;
	wire new_net_387;
	wire new_net_3787;
	wire new_net_3811;
	wire new_net_4406;
	wire new_net_4427;
	wire new_net_4936;
	wire new_net_6540;
	wire new_net_3774;
	wire new_net_7292;
	wire new_net_7663;
	wire new_net_6911;
	wire new_net_3470;
	wire new_net_1533;
	wire new_net_3701;
	wire _0809_;
	wire _0305_;
	wire new_net_3985;
	wire new_net_4186;
	wire new_net_5763;
	wire new_net_6158;
	wire new_net_6608;
	wire new_net_7636;
	wire new_net_8249;
	wire new_net_6267;
	wire new_net_7218;
	wire new_net_2751;
	wire new_net_7135;
	wire new_net_1982;
	wire new_net_3038;
	wire _0647_;
	wire new_net_2929;
	wire new_net_3098;
	wire new_net_2558;
	wire new_net_1639;
	wire new_net_179;
	wire new_net_3415;
	wire new_net_4083;
	wire _0956_;
	wire new_net_5468;
	wire new_net_2348;
	wire new_net_72;
	wire new_net_2285;
	wire new_net_2711;
	wire _0810_;
	wire _0306_;
	wire new_net_4763;
	wire new_net_5295;
	wire new_net_5568;
	wire new_net_6262;
	wire new_net_6378;
	wire new_net_6300;
	wire new_net_7385;
	wire new_net_2623;
	wire new_net_1461;
	wire new_net_3451;
	wire new_net_3490;
	wire new_net_388;
	wire new_net_2645;
	wire new_net_3116;
	wire new_net_4061;
	wire new_net_5317;
	wire new_net_6035;
	wire new_net_6400;
	wire new_net_5503;
	wire new_net_8009;
	wire new_net_6032;
	wire new_net_6688;
	wire new_net_1366;
	wire new_net_7813;
	wire new_net_3551;
	wire new_net_1534;
	wire new_net_2677;
	wire _0307_;
	wire _0811_;
	wire new_net_1761;
	wire new_net_5545;
	wire new_net_7103;
	wire new_net_7322;
	wire new_net_4399;
	wire new_net_6253;
	wire new_net_5518;
	wire new_net_6337;
	wire new_net_6589;
	wire new_net_3416;
	wire new_net_2879;
	wire new_net_3432;
	wire new_net_1856;
	wire new_net_3055;
	wire new_net_3203;
	wire new_net_1640;
	wire new_net_4720;
	wire new_net_4841;
	wire new_net_5191;
	wire new_net_6587;
	wire new_net_8118;
	wire new_net_2533;
	wire new_net_4272;
	wire new_net_7344;
	wire _0060_;
	wire new_net_3975;
	wire new_net_2128;
	wire _0812_;
	wire new_net_3324;
	wire new_net_2805;
	wire new_net_2254;
	wire new_net_73;
	wire _0369_;
	wire _0308_;
	wire new_net_2317;
	wire new_net_2882;
	wire new_net_7272;
	wire new_net_6899;
	wire new_net_5591;
	wire new_net_6448;
	wire new_net_7772;
	wire new_net_1782;
	wire new_net_1388;
	wire new_net_3702;
	wire new_net_3471;
	wire new_net_3986;
	wire new_net_4187;
	wire new_net_5764;
	wire new_net_6159;
	wire new_net_6609;
	wire new_net_7229;
	wire new_net_7854;
	wire new_net_6497;
	wire new_net_7415;
	wire new_net_7705;
	wire new_net_8240;
	wire new_net_4741;
	wire new_net_4125;
	wire new_net_7204;
	wire new_net_3580;
	wire new_net_7794;
	wire new_net_7126;
	wire new_net_2063;
	wire new_net_180;
	wire new_net_3039;
	wire new_net_2930;
	wire new_net_3056;
	wire new_net_2559;
	wire _0813_;
	wire _0309_;
	wire new_net_2112;
	wire new_net_3099;
	wire new_net_6097;
	wire _1096_;
	wire new_net_590;
	wire new_net_2712;
	wire new_net_4764;
	wire new_net_4862;
	wire new_net_5296;
	wire new_net_5569;
	wire new_net_6119;
	wire new_net_6263;
	wire _0680_;
	wire new_net_6756;
	wire new_net_7831;
	wire new_net_7693;
	wire new_net_6286;
	wire new_net_24;
	wire new_net_389;
	wire new_net_1462;
	wire new_net_3452;
	wire new_net_3346;
	wire new_net_3491;
	wire _0814_;
	wire _0310_;
	wire new_net_625;
	wire new_net_2286;
	wire new_net_4370;
	wire new_net_7909;
	wire new_net_5572;
	wire new_net_8076;
	wire new_net_2174;
	wire new_net_5734;
	wire new_net_6931;
	wire new_net_8172;
	wire new_net_1000;
	wire new_net_3552;
	wire new_net_2678;
	wire new_net_3433;
	wire new_net_1535;
	wire new_net_2576;
	wire new_net_4836;
	wire new_net_5546;
	wire new_net_7104;
	wire new_net_6647;
	wire new_net_8052;
	wire new_net_7971;
	wire _0957_;
	wire new_net_2419;
	wire new_net_3752;
	wire new_net_181;
	wire new_net_2880;
	wire new_net_2497;
	wire new_net_3204;
	wire _0815_;
	wire _0311_;
	wire new_net_4842;
	wire new_net_5192;
	wire new_net_5216;
	wire new_net_5422;
	wire new_net_4858;
	wire new_net_8109;
	wire new_net_4216;
	wire new_net_7752;
	wire new_net_2236;
	wire new_net_1642;
	wire new_net_2086;
	wire new_net_3325;
	wire new_net_2806;
	wire new_net_3347;
	wire new_net_74;
	wire new_net_3789;
	wire new_net_3813;
	wire new_net_4429;
	wire new_net_6241;
	wire new_net_7258;
	wire new_net_4092;
	wire new_net_316;
	wire new_net_2004;
	wire new_net_2318;
	wire new_net_390;
	wire new_net_2129;
	wire new_net_1463;
	wire new_net_3703;
	wire _0312_;
	wire _0816_;
	wire new_net_2255;
	wire new_net_3987;
	wire new_net_4188;
	wire new_net_7580;
	wire new_net_8226;
	wire new_net_4727;
	wire new_net_1823;
	wire new_net_6711;
	wire new_net_2560;
	wire new_net_3100;
	wire new_net_2068;
	wire new_net_2858;
	wire new_net_1875;
	wire new_net_3040;
	wire new_net_3593;
	wire new_net_1536;
	wire new_net_2931;
	wire new_net_4062;
	wire new_net_5403;
	wire new_net_5401;
	wire new_net_6099;
	wire _0061_;
	wire new_net_506;
	wire new_net_2713;
	wire new_net_2351;
	wire _0817_;
	wire _0313_;
	wire new_net_4043;
	wire new_net_4863;
	wire new_net_5246;
	wire _0370_;
	wire new_net_5570;
	wire new_net_6728;
	wire new_net_7018;
	wire new_net_7684;
	wire new_net_8047;
	wire _1236_;
	wire new_net_7190;
	wire new_net_1244;
	wire new_net_1643;
	wire new_net_1868;
	wire new_net_3453;
	wire new_net_3492;
	wire new_net_75;
	wire new_net_4449;
	wire new_net_4578;
	wire new_net_5319;
	wire new_net_5958;
	wire new_net_6487;
	wire new_net_2090;
	wire new_net_5268;
	wire new_net_6132;
	wire new_net_6750;
	wire new_net_5725;
	wire new_net_6922;
	wire _0754_;
	wire new_net_6471;
	wire new_net_2287;
	wire new_net_391;
	wire new_net_1464;
	wire new_net_1865;
	wire new_net_2679;
	wire _0818_;
	wire _0314_;
	wire new_net_4408;
	wire new_net_5547;
	wire new_net_7105;
	wire new_net_7846;
	wire new_net_7839;
	wire new_net_7723;
	wire new_net_7890;
	wire new_net_5669;
	wire new_net_3205;
	wire new_net_2859;
	wire new_net_2881;
	wire new_net_4044;
	wire new_net_4371;
	wire new_net_4843;
	wire new_net_5193;
	wire new_net_5217;
	wire new_net_5423;
	wire new_net_6220;
	wire new_net_5055;
	wire new_net_2807;
	wire new_net_3348;
	wire new_net_3645;
	wire new_net_3326;
	wire _0819_;
	wire _0315_;
	wire new_net_3790;
	wire new_net_3814;
	wire new_net_4430;
	wire new_net_6242;
	wire new_net_6225;
	wire new_net_7544;
	wire new_net_7466;
	wire new_net_6675;
	wire new_net_5901;
	wire new_net_2624;
	wire new_net_3704;
	wire new_net_2515;
	wire new_net_3988;
	wire new_net_4189;
	wire new_net_4765;
	wire new_net_5766;
	wire new_net_6161;
	wire new_net_6264;
	wire new_net_6611;
	wire _0958_;
	wire new_net_4389;
	wire new_net_6240;
	wire new_net_7065;
	wire new_net_4886;
	wire new_net_6780;
	wire new_net_7087;
	wire new_net_8038;
	wire _0064_;
	wire _0358_;
	wire _0862_;
	wire new_net_2214;
	wire new_net_3731;
	wire new_net_794;
	wire _1072_;
	wire new_net_3529;
	wire _0568_;
	wire new_net_614;
	wire new_net_4223;
	wire new_net_8261;
	wire new_net_444;
	wire new_net_2050;
	wire new_net_2815;
	wire new_net_2062;
	wire new_net_2587;
	wire new_net_3188;
	wire new_net_3823;
	wire new_net_3847;
	wire new_net_5657;
	wire new_net_6770;
	wire new_net_5348;
	wire new_net_4820;
	wire new_net_4818;
	wire _0065_;
	wire _0359_;
	wire new_net_724;
	wire new_net_2957;
	wire _0863_;
	wire new_net_1080;
	wire new_net_829;
	wire _1073_;
	wire _0569_;
	wire new_net_3765;
	wire new_net_6506;
	wire new_net_6771;
	wire new_net_3235;
	wire new_net_4118;
	wire new_net_4233;
	wire new_net_4774;
	wire new_net_6048;
	wire new_net_6273;
	wire new_net_6376;
	wire new_net_6498;
	wire new_net_7348;
	wire new_net_8066;
	wire new_net_6528;
	wire new_net_4296;
	wire new_net_4076;
	wire new_net_7188;
	wire new_net_7540;
	wire new_net_2451;
	wire _0570_;
	wire _0864_;
	wire _0066_;
	wire _0360_;
	wire new_net_2653;
	wire new_net_2349;
	wire new_net_795;
	wire new_net_1927;
	wire _1074_;
	wire new_net_6963;
	wire new_net_8280;
	wire new_net_7874;
	wire new_net_5983;
	wire new_net_7302;
	wire new_net_445;
	wire new_net_2688;
	wire new_net_3355;
	wire new_net_2608;
	wire new_net_3125;
	wire new_net_4921;
	wire new_net_7325;
	wire new_net_7476;
	wire new_net_8213;
	wire new_net_6945;
	wire new_net_8181;
	wire new_net_5909;
	wire new_net_7150;
	wire _0067_;
	wire _0361_;
	wire _0571_;
	wire new_net_1997;
	wire _0865_;
	wire new_net_2025;
	wire new_net_1081;
	wire new_net_830;
	wire _1075_;
	wire new_net_2002;
	wire new_net_5880;
	wire new_net_7250;
	wire new_net_582;
	wire new_net_3732;
	wire new_net_3530;
	wire new_net_4234;
	wire new_net_5435;
	wire new_net_5904;
	wire new_net_6219;
	wire new_net_7017;
	wire new_net_7199;
	wire new_net_7989;
	wire new_net_6310;
	wire new_net_6855;
	wire new_net_6437;
	wire _0068_;
	wire _0362_;
	wire new_net_2152;
	wire _0866_;
	wire new_net_2215;
	wire new_net_2816;
	wire _1076_;
	wire new_net_2588;
	wire _0572_;
	wire new_net_616;
	wire new_net_5707;
	wire new_net_6698;
	wire new_net_6877;
	wire new_net_7823;
	wire new_net_5841;
	wire new_net_725;
	wire new_net_4664;
	wire new_net_5060;
	wire new_net_5084;
	wire new_net_5333;
	wire new_net_5637;
	wire new_net_6792;
	wire new_net_7722;
	wire new_net_7868;
	wire new_net_8006;
	wire new_net_7504;
	wire new_net_4909;
	wire new_net_4492;
	wire _1077_;
	wire _0069_;
	wire _0363_;
	wire new_net_1729;
	wire _0867_;
	wire new_net_29;
	wire new_net_3236;
	wire _0573_;
	wire new_net_4119;
	wire new_net_4775;
	wire new_net_7649;
	wire new_net_796;
	wire new_net_2752;
	wire new_net_2654;
	wire new_net_3069;
	wire new_net_3766;
	wire new_net_5779;
	wire new_net_6198;
	wire new_net_6423;
	wire new_net_6521;
	wire new_net_7268;
	wire new_net_6541;
	wire _0070_;
	wire _0364_;
	wire new_net_446;
	wire _0868_;
	wire new_net_2689;
	wire new_net_3503;
	wire new_net_2064;
	wire _1078_;
	wire _0574_;
	wire new_net_617;
	wire new_net_7049;
	wire new_net_8250;
	wire new_net_4751;
	wire new_net_7136;
	wire new_net_6069;
	wire new_net_726;
	wire new_net_831;
	wire new_net_1082;
	wire new_net_2781;
	wire new_net_2088;
	wire new_net_4203;
	wire new_net_4798;
	wire new_net_4877;
	wire new_net_4901;
	wire new_net_6175;
	wire new_net_7241;
	wire _0575_;
	wire _0869_;
	wire _0071_;
	wire new_net_30;
	wire new_net_3733;
	wire _0365_;
	wire new_net_3216;
	wire _1079_;
	wire new_net_3531;
	wire new_net_5436;
	wire new_net_6379;
	wire new_net_4309;
	wire new_net_7386;
	wire new_net_4018;
	wire new_net_2606;
	wire new_net_797;
	wire new_net_2529;
	wire new_net_2817;
	wire new_net_3070;
	wire new_net_2589;
	wire new_net_3825;
	wire new_net_3849;
	wire new_net_5659;
	wire new_net_5698;
	wire new_net_6401;
	wire new_net_6318;
	wire new_net_6033;
	wire new_net_6689;
	wire new_net_4615;
	wire new_net_7814;
	wire _0072_;
	wire _0576_;
	wire new_net_618;
	wire new_net_3145;
	wire new_net_2153;
	wire new_net_2634;
	wire new_net_447;
	wire new_net_2005;
	wire new_net_2020;
	wire _0870_;
	wire new_net_7323;
	wire new_net_5519;
	wire new_net_6338;
	wire new_net_6590;
	wire new_net_727;
	wire new_net_832;
	wire new_net_1083;
	wire new_net_1734;
	wire new_net_1996;
	wire new_net_3237;
	wire new_net_4001;
	wire new_net_4120;
	wire new_net_4776;
	wire new_net_6275;
	wire new_net_8119;
	wire new_net_7345;
	wire new_net_7767;
	wire _1081_;
	wire _0073_;
	wire _0577_;
	wire new_net_3767;
	wire new_net_2753;
	wire new_net_2453;
	wire new_net_2655;
	wire new_net_3709;
	wire _0871_;
	wire _0367_;
	wire new_net_6900;
	wire new_net_7273;
	wire new_net_4390;
	wire new_net_798;
	wire new_net_3504;
	wire new_net_3127;
	wire new_net_2635;
	wire new_net_2940;
	wire new_net_2690;
	wire new_net_4460;
	wire new_net_4923;
	wire new_net_4956;
	wire new_net_5905;
	wire new_net_7416;
	wire new_net_7706;
	wire new_net_8241;
	wire new_net_4407;
	wire new_net_7205;
	wire new_net_7795;
	wire new_net_7127;
	wire _1082_;
	wire _0074_;
	wire _0578_;
	wire new_net_619;
	wire new_net_2085;
	wire _0872_;
	wire new_net_2089;
	wire _0368_;
	wire new_net_2833;
	wire new_net_4204;
	wire new_net_6893;
	wire _0928_;
	wire new_net_4224;
	wire new_net_6120;
	wire new_net_728;
	wire new_net_3710;
	wire new_net_3734;
	wire new_net_5437;
	wire new_net_7028;
	wire new_net_7991;
	wire new_net_6287;
	wire new_net_7861;
	wire new_net_7372;
	wire new_net_7912;
	wire new_net_2391;
	wire _0579_;
	wire _0873_;
	wire _1083_;
	wire new_net_2590;
	wire new_net_2607;
	wire _0075_;
	wire new_net_2818;
	wire new_net_2782;
	wire new_net_31;
	wire new_net_5573;
	wire new_net_6019;
	wire new_net_5735;
	wire new_net_6932;
	wire new_net_8173;
	wire new_net_3866;
	wire new_net_3523;
	wire new_net_448;
	wire new_net_799;
	wire new_net_2941;
	wire new_net_4666;
	wire new_net_5062;
	wire new_net_5086;
	wire new_net_5335;
	wire new_net_5639;
	wire new_net_7724;
	wire new_net_7972;
	wire new_net_833;
	wire new_net_3238;
	wire _0580_;
	wire _0874_;
	wire _0076_;
	wire _1084_;
	wire new_net_620;
	wire new_net_2154;
	wire new_net_1767;
	wire new_net_2217;
	wire new_net_4859;
	wire new_net_4215;
	wire new_net_7753;
	wire new_net_585;
	wire new_net_729;
	wire new_net_1085;
	wire new_net_3768;
	wire new_net_2754;
	wire new_net_3146;
	wire new_net_2656;
	wire new_net_5781;
	wire new_net_6200;
	wire new_net_6425;
	wire new_net_7259;
	wire new_net_5127;
	wire _0371_;
	wire new_net_2691;
	wire new_net_2958;
	wire _1085_;
	wire _0581_;
	wire _0875_;
	wire _0077_;
	wire new_net_3128;
	wire new_net_2636;
	wire new_net_4461;
	wire new_net_6007;
	wire new_net_7581;
	wire new_net_8227;
	wire new_net_6424;
	wire new_net_8205;
	wire new_net_449;
	wire new_net_800;
	wire new_net_4205;
	wire new_net_4800;
	wire new_net_4879;
	wire new_net_4903;
	wire new_net_6050;
	wire new_net_6177;
	wire new_net_6299;
	wire new_net_6402;
	wire new_net_6729;
	wire _0372_;
	wire _1086_;
	wire _0078_;
	wire new_net_834;
	wire new_net_3356;
	wire _0582_;
	wire new_net_621;
	wire new_net_3735;
	wire new_net_2528;
	wire new_net_3711;
	wire new_net_7685;
	wire new_net_4655;
	wire new_net_7191;
	wire new_net_5959;
	wire new_net_2819;
	wire new_net_586;
	wire new_net_730;
	wire new_net_1086;
	wire new_net_1928;
	wire new_net_2959;
	wire new_net_2591;
	wire new_net_2609;
	wire new_net_2011;
	wire new_net_2886;
	wire new_net_6751;
	wire new_net_5481;
	wire new_net_7629;
	wire new_net_5726;
	wire new_net_6923;
	wire new_net_4674;
	wire new_net_6472;
	wire new_net_7007;
	wire new_net_32;
	wire _0373_;
	wire _0583_;
	wire _0877_;
	wire _1087_;
	wire _0079_;
	wire new_net_2942;
	wire new_net_4667;
	wire new_net_5063;
	wire new_net_5336;
	wire new_net_7847;
	wire new_net_7840;
	wire new_net_7891;
	wire new_net_5007;
	wire new_net_7528;
	wire new_net_801;
	wire new_net_3239;
	wire new_net_4003;
	wire new_net_4098;
	wire new_net_4122;
	wire new_net_4778;
	wire new_net_6277;
	wire new_net_4850;
	wire new_net_6380;
	wire new_net_7019;
	wire new_net_5636;
	wire new_net_6047;
	wire new_net_2218;
	wire _0584_;
	wire _0878_;
	wire _0374_;
	wire new_net_2084;
	wire new_net_3071;
	wire _1088_;
	wire new_net_622;
	wire new_net_3769;
	wire _0080_;
	wire new_net_6226;
	wire new_net_7467;
	wire new_net_4532;
	wire new_net_6676;
	wire new_net_5902;
	wire new_net_3217;
	wire new_net_587;
	wire new_net_731;
	wire new_net_2692;
	wire new_net_3129;
	wire new_net_2637;
	wire new_net_2887;
	wire new_net_4925;
	wire new_net_4955;
	wire new_net_5907;
	wire new_net_4103;
	wire new_net_5218;
	wire new_net_7066;
	wire new_net_6781;
	wire new_net_450;
	wire _1089_;
	wire _0585_;
	wire _0879_;
	wire _0375_;
	wire new_net_2834;
	wire _0081_;
	wire new_net_4206;
	wire new_net_4801;
	wire new_net_4880;
	wire new_net_6091;
	wire new_net_7088;
	wire new_net_5238;
	wire new_net_8039;
	wire new_net_3712;
	wire new_net_3736;
	wire new_net_802;
	wire new_net_835;
	wire new_net_4235;
	wire new_net_7993;
	wire new_net_5115;
	wire new_net_8262;
	wire _1090_;
	wire _0586_;
	wire _0880_;
	wire _0376_;
	wire new_net_1087;
	wire new_net_2820;
	wire new_net_2592;
	wire new_net_623;
	wire _0082_;
	wire new_net_2393;
	wire new_net_2016;
	wire new_net_588;
	wire new_net_732;
	wire new_net_4668;
	wire new_net_5064;
	wire new_net_5337;
	wire new_net_7726;
	wire new_net_7872;
	wire new_net_4634;
	wire new_net_6507;
	wire new_net_2014;
	wire new_net_2640;
	wire new_net_451;
	wire _0587_;
	wire _0881_;
	wire _1091_;
	wire _0377_;
	wire new_net_3505;
	wire new_net_3240;
	wire _0083_;
	wire new_net_5170;
	wire new_net_6529;
	wire new_net_6790;
	wire new_net_2527;
	wire new_net_803;
	wire new_net_3358;
	wire new_net_836;
	wire new_net_3524;
	wire new_net_3532;
	wire new_net_3770;
	wire new_net_2756;
	wire new_net_4236;
	wire new_net_4683;
	wire new_net_6964;
	wire new_net_5071;
	wire new_net_2156;
	wire _0882_;
	wire _0588_;
	wire _1092_;
	wire new_net_33;
	wire _0378_;
	wire new_net_1088;
	wire new_net_2693;
	wire new_net_2219;
	wire new_net_624;
	wire new_net_4713;
	wire new_net_3824;
	wire new_net_6946;
	wire new_net_4688;
	wire new_net_4428;
	wire new_net_5910;
	wire new_net_2638;
	wire new_net_733;
	wire new_net_4802;
	wire new_net_4881;
	wire new_net_4905;
	wire new_net_5662;
	wire new_net_6052;
	wire new_net_6179;
	wire new_net_6301;
	wire new_net_6404;
	wire new_net_7151;
	wire new_net_6662;
	wire new_net_3713;
	wire _0085_;
	wire _0379_;
	wire _0883_;
	wire new_net_3737;
	wire _1093_;
	wire _0589_;
	wire new_net_5641;
	wire new_net_4377;
	wire new_net_5686;
	wire new_net_4048;
	wire new_net_6311;
	wire new_net_6856;
	wire new_net_6849;
	wire new_net_7396;
	wire new_net_804;
	wire new_net_837;
	wire new_net_2010;
	wire new_net_2821;
	wire new_net_2066;
	wire new_net_3829;
	wire new_net_3853;
	wire new_net_4462;
	wire new_net_6438;
	wire new_net_6503;
	wire new_net_7568;
	wire new_net_5708;
	wire new_net_5340;
	wire new_net_2421;
	wire _0086_;
	wire _0380_;
	wire _0884_;
	wire new_net_34;
	wire new_net_1784;
	wire new_net_1089;
	wire new_net_3508;
	wire _1094_;
	wire new_net_589;
	wire new_net_5842;
	wire new_net_6871;
	wire new_net_7824;
	wire new_net_7505;
	wire new_net_4569;
	wire new_net_452;
	wire new_net_734;
	wire new_net_2657;
	wire new_net_3241;
	wire new_net_4005;
	wire new_net_4100;
	wire new_net_4124;
	wire new_net_4780;
	wire new_net_5439;
	wire new_net_5908;
	wire new_net_2757;
	wire new_net_2457;
	wire _0087_;
	wire _0381_;
	wire new_net_1765;
	wire new_net_2658;
	wire _0885_;
	wire new_net_3072;
	wire new_net_3359;
	wire _1095_;
	wire new_net_4967;
	wire new_net_4969;
	wire new_net_4335;
	wire new_net_4938;
	wire new_net_7667;
	wire new_net_3131;
	wire new_net_1998;
	wire new_net_805;
	wire new_net_838;
	wire new_net_2694;
	wire new_net_2943;
	wire new_net_3506;
	wire new_net_1804;
	wire new_net_4463;
	wire new_net_4927;
	wire new_net_5028;
	wire new_net_7665;
	wire new_net_7050;
	wire new_net_7638;
	wire new_net_7222;
	wire new_net_6269;
	wire new_net_7220;
	wire _0592_;
	wire new_net_626;
	wire _0088_;
	wire _0382_;
	wire new_net_2157;
	wire new_net_2639;
	wire new_net_2009;
	wire _0886_;
	wire new_net_35;
	wire new_net_2220;
	wire new_net_6648;
	wire new_net_453;
	wire new_net_1974;
	wire new_net_2660;
	wire new_net_3714;
	wire new_net_3738;
	wire new_net_5338;
	wire new_net_5642;
	wire new_net_7242;
	wire new_net_7995;
	wire new_net_6302;
	wire _0593_;
	wire new_net_2395;
	wire _0089_;
	wire _0383_;
	wire new_net_2888;
	wire _0887_;
	wire new_net_2822;
	wire new_net_3073;
	wire _1097_;
	wire new_net_3830;
	wire new_net_5505;
	wire new_net_8011;
	wire new_net_6319;
	wire new_net_6034;
	wire new_net_839;
	wire new_net_1090;
	wire new_net_2890;
	wire new_net_2022;
	wire new_net_4670;
	wire new_net_5066;
	wire new_net_7630;
	wire new_net_7728;
	wire new_net_7815;
	wire new_net_6174;
	wire new_net_591;
	wire _0594_;
	wire new_net_627;
	wire _1098_;
	wire _0090_;
	wire new_net_2526;
	wire new_net_735;
	wire new_net_1760;
	wire _0888_;
	wire new_net_36;
	wire new_net_6339;
	wire new_net_6591;
	wire new_net_8120;
	wire new_net_4274;
	wire new_net_6100;
	wire new_net_7999;
	wire new_net_7346;
	wire new_net_454;
	wire new_net_2758;
	wire new_net_3772;
	wire new_net_3360;
	wire new_net_4906;
	wire new_net_5785;
	wire new_net_6204;
	wire new_net_6429;
	wire new_net_6527;
	wire new_net_7274;
	wire new_net_6901;
	wire new_net_6450;
	wire _1099_;
	wire new_net_1803;
	wire new_net_3533;
	wire _0595_;
	wire _0091_;
	wire new_net_2889;
	wire _0889_;
	wire _0385_;
	wire new_net_806;
	wire new_net_2695;
	wire new_net_7417;
	wire new_net_7591;
	wire new_net_8242;
	wire new_net_4127;
	wire new_net_7206;
	wire new_net_7796;
	wire new_net_7128;
	wire new_net_840;
	wire new_net_1091;
	wire new_net_4804;
	wire new_net_4883;
	wire new_net_5664;
	wire new_net_6054;
	wire new_net_6061;
	wire new_net_5157;
	wire new_net_6181;
	wire new_net_6303;
	wire new_net_5045;
	wire _1100_;
	wire new_net_592;
	wire new_net_2593;
	wire new_net_628;
	wire _0596_;
	wire _0890_;
	wire _0092_;
	wire new_net_2158;
	wire new_net_736;
	wire new_net_2659;
	wire new_net_7029;
	wire new_net_7695;
	wire new_net_6288;
	wire new_net_7373;
	wire new_net_3534;
	wire new_net_455;
	wire new_net_2823;
	wire new_net_3831;
	wire new_net_3855;
	wire new_net_6280;
	wire new_net_6505;
	wire new_net_8200;
	wire new_net_5574;
	wire new_net_5491;
	wire new_net_6933;
	wire new_net_8174;
	wire new_net_6482;
	wire new_net_2067;
	wire _1101_;
	wire _0597_;
	wire _0891_;
	wire _0093_;
	wire _0387_;
	wire new_net_807;
	wire new_net_5067;
	wire new_net_4838;
	wire new_net_7729;
	wire new_net_7973;
	wire new_net_3243;
	wire new_net_2594;
	wire new_net_841;
	wire new_net_1092;
	wire new_net_2001;
	wire new_net_3148;
	wire new_net_3220;
	wire new_net_4007;
	wire new_net_4102;
	wire new_net_4126;
	wire new_net_4860;
	wire _0388_;
	wire _1102_;
	wire _0094_;
	wire _0598_;
	wire new_net_629;
	wire new_net_3773;
	wire new_net_2759;
	wire new_net_2459;
	wire new_net_737;
	wire _0892_;
	wire new_net_7754;
	wire new_net_7260;
	wire new_net_7477;
	wire new_net_5128;
	wire new_net_2015;
	wire new_net_2696;
	wire new_net_2944;
	wire new_net_2107;
	wire new_net_2035;
	wire new_net_4465;
	wire new_net_4929;
	wire new_net_5090;
	wire new_net_5339;
	wire new_net_5643;
	wire new_net_7582;
	wire new_net_8228;
	wire new_net_4729;
	wire new_net_3848;
	wire new_net_3846;
	wire _0389_;
	wire new_net_1763;
	wire _0095_;
	wire _1103_;
	wire _0599_;
	wire new_net_3149;
	wire new_net_2641;
	wire _0893_;
	wire new_net_4805;
	wire new_net_4884;
	wire new_net_5405;
	wire new_net_6197;
	wire new_net_3716;
	wire new_net_593;
	wire new_net_1093;
	wire new_net_2003;
	wire new_net_2012;
	wire new_net_3740;
	wire new_net_7631;
	wire new_net_7875;
	wire new_net_7997;
	wire new_net_6730;
	wire new_net_8049;
	wire new_net_7020;
	wire new_net_7686;
	wire new_net_4168;
	wire new_net_7192;
	wire new_net_2222;
	wire _0390_;
	wire new_net_2824;
	wire _0600_;
	wire _0894_;
	wire _0096_;
	wire _1104_;
	wire new_net_2610;
	wire new_net_2397;
	wire _1136_;
	wire new_net_5270;
	wire new_net_6134;
	wire new_net_7512;
	wire new_net_5482;
	wire new_net_5727;
	wire new_net_6924;
	wire new_net_6473;
	wire new_net_2945;
	wire new_net_808;
	wire new_net_4685;
	wire new_net_5068;
	wire new_net_7008;
	wire new_net_7921;
	wire new_net_7848;
	wire new_net_7841;
	wire new_net_7725;
	wire new_net_7892;
	wire _0391_;
	wire new_net_3221;
	wire new_net_842;
	wire new_net_3244;
	wire _0601_;
	wire _0895_;
	wire _1105_;
	wire new_net_2595;
	wire _0097_;
	wire new_net_4008;
	wire new_net_7529;
	wire new_net_5800;
	wire new_net_4336;
	wire new_net_3074;
	wire new_net_39;
	wire new_net_594;
	wire new_net_630;
	wire new_net_2611;
	wire new_net_2760;
	wire new_net_4237;
	wire new_net_4908;
	wire new_net_5787;
	wire new_net_6206;
	wire new_net_6628;
	wire new_net_7546;
	wire new_net_7251;
	wire new_net_6227;
	wire new_net_7468;
	wire new_net_6677;
	wire new_net_457;
	wire _0392_;
	wire new_net_2697;
	wire _1106_;
	wire _0602_;
	wire _0896_;
	wire _0098_;
	wire new_net_4238;
	wire new_net_4466;
	wire new_net_4930;
	wire new_net_4890;
	wire new_net_7067;
	wire new_net_5141;
	wire new_net_3509;
	wire new_net_809;
	wire new_net_3150;
	wire new_net_2642;
	wire new_net_4885;
	wire new_net_5666;
	wire new_net_6056;
	wire new_net_6183;
	wire new_net_6281;
	wire new_net_6305;
	wire new_net_8192;
	wire new_net_5440;
	wire new_net_3717;
	wire _0897_;
	wire new_net_3741;
	wire _0393_;
	wire new_net_1094;
	wire new_net_3075;
	wire _1107_;
	wire new_net_843;
	wire _0603_;
	wire _0099_;
	wire new_net_7089;
	wire new_net_8040;
	wire new_net_2825;
	wire new_net_3361;
	wire new_net_40;
	wire new_net_631;
	wire new_net_739;
	wire new_net_3536;
	wire new_net_3403;
	wire new_net_2891;
	wire new_net_3833;
	wire new_net_3857;
	wire new_net_4932;
	wire new_net_4517;
	wire new_net_1872;
	wire new_net_3190;
	wire new_net_5433;
	wire new_net_4822;
	wire new_net_2160;
	wire new_net_458;
	wire new_net_2223;
	wire _0394_;
	wire _0604_;
	wire _0898_;
	wire _1108_;
	wire new_net_2023;
	wire _0100_;
	wire new_net_5069;
	wire new_net_6508;
	wire new_net_7643;
	wire new_net_8251;
	wire new_net_4136;
	wire new_net_2596;
	wire new_net_3222;
	wire new_net_1930;
	wire new_net_3245;
	wire new_net_4009;
	wire new_net_4104;
	wire new_net_4128;
	wire new_net_4784;
	wire new_net_5443;
	wire new_net_5912;
	wire new_net_6530;
	wire new_net_2461;
	wire new_net_1885;
	wire _0395_;
	wire new_net_1095;
	wire _0605_;
	wire _0899_;
	wire new_net_844;
	wire _1109_;
	wire new_net_595;
	wire _0101_;
	wire new_net_4078;
	wire new_net_7542;
	wire new_net_6965;
	wire new_net_7692;
	wire new_net_7876;
	wire new_net_632;
	wire new_net_740;
	wire new_net_2698;
	wire new_net_2612;
	wire new_net_3775;
	wire new_net_4467;
	wire new_net_4672;
	wire new_net_4931;
	wire new_net_5092;
	wire new_net_5341;
	wire new_net_5985;
	wire new_net_7304;
	wire new_net_7933;
	wire new_net_459;
	wire _0606_;
	wire _0900_;
	wire _0396_;
	wire new_net_810;
	wire new_net_3510;
	wire new_net_3525;
	wire _1110_;
	wire new_net_2108;
	wire _0102_;
	wire new_net_5911;
	wire new_net_8183;
	wire new_net_7152;
	wire new_net_7324;
	wire new_net_3718;
	wire new_net_3742;
	wire new_net_3076;
	wire new_net_7633;
	wire new_net_7731;
	wire new_net_7877;
	wire new_net_4604;
	wire _0103_;
	wire new_net_2399;
	wire new_net_2785;
	wire new_net_41;
	wire _1111_;
	wire _0607_;
	wire _0901_;
	wire _0397_;
	wire new_net_1096;
	wire new_net_2826;
	wire new_net_6857;
	wire new_net_6439;
	wire new_net_7397;
	wire new_net_7774;
	wire new_net_8021;
	wire new_net_633;
	wire new_net_2960;
	wire new_net_5070;
	wire new_net_6700;
	wire new_net_6879;
	wire new_net_7825;
	wire new_net_5843;
	wire _0104_;
	wire new_net_2161;
	wire new_net_460;
	wire _1112_;
	wire _0902_;
	wire new_net_2224;
	wire _0398_;
	wire new_net_811;
	wire new_net_1832;
	wire new_net_3246;
	wire new_net_3942;
	wire new_net_6612;
	wire new_net_2762;
	wire new_net_2892;
	wire new_net_845;
	wire new_net_2597;
	wire new_net_4687;
	wire new_net_4807;
	wire new_net_4910;
	wire new_net_5789;
	wire new_net_6057;
	wire new_net_6208;
	wire new_net_6121;
	wire new_net_5603;
	wire new_net_2613;
	wire new_net_3776;
	wire _0105_;
	wire new_net_1999;
	wire new_net_741;
	wire _0609_;
	wire _0903_;
	wire _1113_;
	wire new_net_42;
	wire _0399_;
	wire new_net_7295;
	wire new_net_7668;
	wire new_net_7913;
	wire new_net_7051;
	wire new_net_6973;
	wire new_net_7639;
	wire new_net_4753;
	wire new_net_5658;
	wire new_net_3152;
	wire new_net_2525;
	wire new_net_1730;
	wire new_net_1887;
	wire new_net_634;
	wire new_net_2036;
	wire new_net_3511;
	wire new_net_2835;
	wire new_net_4887;
	wire new_net_5668;
	wire new_net_7138;
	wire new_net_6071;
	wire new_net_6649;
	wire new_net_2415;
	wire _1138_;
	wire new_net_7243;
	wire new_net_7039;
	wire new_net_6381;
	wire new_net_7388;
	wire new_net_4020;
	wire new_net_1186;
	wire new_net_1150;
	wire new_net_2319;
	wire new_net_149;
	wire new_net_392;
	wire new_net_932;
	wire _0148_;
	wire _0652_;
	wire _1156_;
	wire new_net_2736;
	wire new_net_5700;
	wire new_net_6403;
	wire new_net_8012;
	wire new_net_6320;
	wire new_net_7816;
	wire new_net_114;
	wire new_net_1008;
	wire new_net_1044;
	wire new_net_3176;
	wire new_net_5846;
	wire _0690_;
	wire new_net_5925;
	wire new_net_7371;
	wire new_net_4965;
	wire new_net_7395;
	wire new_net_6342;
	wire new_net_5521;
	wire new_net_6592;
	wire new_net_1911;
	wire new_net_2042;
	wire new_net_3020;
	wire _0149_;
	wire _0653_;
	wire _1157_;
	wire new_net_760;
	wire new_net_4559;
	wire new_net_5229;
	wire new_net_5581;
	wire new_net_8123;
	wire new_net_8121;
	wire new_net_6101;
	wire new_net_8000;
	wire new_net_7347;
	wire new_net_2257;
	wire new_net_1956;
	wire new_net_3271;
	wire new_net_1808;
	wire new_net_3289;
	wire new_net_479;
	wire new_net_971;
	wire new_net_4141;
	wire new_net_5251;
	wire new_net_5378;
	wire new_net_5457;
	wire new_net_5543;
	wire new_net_7275;
	wire new_net_6902;
	wire new_net_5594;
	wire new_net_6451;
	wire new_net_546;
	wire new_net_1115;
	wire new_net_2288;
	wire new_net_1151;
	wire new_net_150;
	wire new_net_1187;
	wire new_net_1400;
	wire new_net_393;
	wire new_net_933;
	wire new_net_690;
	wire new_net_288;
	wire new_net_7708;
	wire new_net_7592;
	wire new_net_8243;
	wire new_net_7207;
	wire new_net_7797;
	wire new_net_43;
	wire new_net_115;
	wire new_net_511;
	wire new_net_1009;
	wire new_net_3305;
	wire new_net_3327;
	wire new_net_1045;
	wire new_net_4481;
	wire new_net_4504;
	wire new_net_4945;
	wire new_net_863;
	wire new_net_2724;
	wire new_net_1850;
	wire new_net_653;
	wire _0151_;
	wire _1159_;
	wire _0655_;
	wire new_net_3163;
	wire new_net_761;
	wire new_net_4596;
	wire new_net_7030;
	wire new_net_7696;
	wire new_net_7863;
	wire new_net_7374;
	wire new_net_5972;
	wire new_net_7954;
	wire new_net_14;
	wire new_net_972;
	wire new_net_1800;
	wire new_net_4250;
	wire new_net_4579;
	wire new_net_5703;
	wire new_net_5722;
	wire new_net_5801;
	wire new_net_6543;
	wire new_net_6646;
	wire new_net_2361;
	wire new_net_6021;
	wire new_net_5737;
	wire new_net_6934;
	wire new_net_8175;
	wire new_net_6483;
	wire new_net_1116;
	wire new_net_1152;
	wire new_net_151;
	wire new_net_1401;
	wire new_net_2320;
	wire new_net_934;
	wire _0656_;
	wire _0152_;
	wire _1160_;
	wire new_net_691;
	wire new_net_4839;
	wire new_net_7974;
	wire new_net_1249;
	wire new_net_44;
	wire new_net_116;
	wire new_net_512;
	wire new_net_1010;
	wire new_net_1046;
	wire new_net_4560;
	wire new_net_5230;
	wire new_net_6070;
	wire new_net_7164;
	wire new_net_7291;
	wire new_net_7755;
	wire new_net_864;
	wire new_net_2737;
	wire new_net_3272;
	wire _0153_;
	wire _0657_;
	wire _1161_;
	wire new_net_654;
	wire new_net_2725;
	wire new_net_480;
	wire new_net_762;
	wire new_net_5413;
	wire new_net_7261;
	wire new_net_7478;
	wire new_net_7650;
	wire new_net_394;
	wire new_net_547;
	wire new_net_1188;
	wire new_net_4821;
	wire new_net_5480;
	wire new_net_5504;
	wire new_net_5681;
	wire new_net_6222;
	wire new_net_6897;
	wire new_net_8010;
	wire new_net_6009;
	wire new_net_7583;
	wire new_net_8229;
	wire new_net_6426;
	wire new_net_2052;
	wire new_net_2057;
	wire new_net_1117;
	wire new_net_2289;
	wire new_net_7;
	wire new_net_1153;
	wire new_net_152;
	wire _1162_;
	wire _0154_;
	wire _0658_;
	wire new_net_6805;
	wire new_net_45;
	wire new_net_117;
	wire new_net_513;
	wire new_net_1011;
	wire new_net_1047;
	wire new_net_3164;
	wire new_net_6625;
	wire new_net_6731;
	wire new_net_7021;
	wire new_net_7499;
	wire new_net_8050;
	wire new_net_7687;
	wire new_net_8146;
	wire new_net_4657;
	wire new_net_7193;
	wire new_net_481;
	wire new_net_763;
	wire new_net_1905;
	wire new_net_865;
	wire new_net_2860;
	wire _1163_;
	wire _0155_;
	wire _0659_;
	wire new_net_973;
	wire new_net_5582;
	wire new_net_6135;
	wire new_net_6753;
	wire new_net_5483;
	wire new_net_5728;
	wire new_net_6925;
	wire new_net_6474;
	wire new_net_395;
	wire new_net_548;
	wire new_net_692;
	wire new_net_1189;
	wire new_net_1402;
	wire new_net_2514;
	wire new_net_4157;
	wire new_net_5848;
	wire new_net_5927;
	wire new_net_7009;
	wire new_net_7922;
	wire _0936_;
	wire new_net_7842;
	wire new_net_6947;
	wire new_net_4689;
	wire new_net_7893;
	wire new_net_1941;
	wire new_net_1118;
	wire new_net_1154;
	wire new_net_2321;
	wire _0156_;
	wire _1164_;
	wire _0660_;
	wire new_net_153;
	wire new_net_936;
	wire new_net_1806;
	wire new_net_7447;
	wire new_net_1658;
	wire new_net_4852;
	wire new_net_3958;
	wire new_net_5638;
	wire new_net_5767;
	wire new_net_6636;
	wire new_net_1012;
	wire new_net_1048;
	wire new_net_2726;
	wire new_net_118;
	wire new_net_514;
	wire new_net_655;
	wire new_net_1970;
	wire new_net_2738;
	wire new_net_3273;
	wire new_net_4143;
	wire new_net_4451;
	wire new_net_5765;
	wire new_net_7252;
	wire new_net_7469;
	wire new_net_4791;
	wire new_net_6312;
	wire new_net_6678;
	wire new_net_2501;
	wire new_net_482;
	wire new_net_764;
	wire new_net_866;
	wire _0661_;
	wire _0157_;
	wire _1165_;
	wire new_net_2861;
	wire new_net_974;
	wire new_net_4158;
	wire new_net_5995;
	wire new_net_7569;
	wire new_net_4105;
	wire new_net_5220;
	wire new_net_7068;
	wire new_net_5142;
	wire new_net_8193;
	wire new_net_693;
	wire new_net_1403;
	wire new_net_1740;
	wire new_net_1952;
	wire new_net_3307;
	wire new_net_4483;
	wire new_net_4506;
	wire new_net_4947;
	wire new_net_5357;
	wire new_net_5826;
	wire new_net_5441;
	wire _0765_;
	wire new_net_228;
	wire new_net_7090;
	wire new_net_1155;
	wire new_net_46;
	wire new_net_1940;
	wire new_net_2290;
	wire _0662_;
	wire _0158_;
	wire _1166_;
	wire new_net_154;
	wire new_net_2185;
	wire new_net_937;
	wire new_net_6894;
	wire new_net_935;
	wire new_net_8264;
	wire new_net_1922;
	wire new_net_119;
	wire new_net_515;
	wire new_net_656;
	wire new_net_1013;
	wire new_net_1049;
	wire new_net_5231;
	wire new_net_5583;
	wire new_net_5705;
	wire new_net_5724;
	wire new_net_4518;
	wire new_net_4823;
	wire new_net_975;
	wire new_net_483;
	wire new_net_765;
	wire new_net_15;
	wire new_net_549;
	wire _1167_;
	wire _0159_;
	wire _0663_;
	wire new_net_1190;
	wire new_net_1957;
	wire new_net_3619;
	wire new_net_4636;
	wire new_net_6270;
	wire new_net_2499;
	wire new_net_1845;
	wire new_net_1119;
	wire new_net_4562;
	wire new_net_4581;
	wire new_net_6072;
	wire new_net_254;
	wire new_net_6366;
	wire new_net_6898;
	wire new_net_7166;
	wire new_net_7293;
	wire _0969_;
	wire new_net_6531;
	wire new_net_3224;
	wire new_net_2037;
	wire new_net_47;
	wire _1168_;
	wire _0160_;
	wire new_net_1156;
	wire new_net_2322;
	wire new_net_155;
	wire new_net_2739;
	wire new_net_3274;
	wire _0664_;
	wire _0446_;
	wire new_net_4676;
	wire new_net_1014;
	wire new_net_1050;
	wire new_net_120;
	wire new_net_516;
	wire new_net_657;
	wire new_net_867;
	wire new_net_3665;
	wire new_net_4374;
	wire new_net_4600;
	wire new_net_4716;
	wire new_net_7305;
	wire new_net_3826;
	wire new_net_5746;
	wire new_net_7934;
	wire new_net_5914;
	wire new_net_397;
	wire new_net_694;
	wire new_net_976;
	wire new_net_3308;
	wire new_net_766;
	wire _0665_;
	wire _0161_;
	wire _1169_;
	wire new_net_550;
	wire new_net_1191;
	wire new_net_4586;
	wire new_net_6954;
	wire new_net_6664;
	wire new_net_1810;
	wire new_net_2513;
	wire new_net_8;
	wire new_net_1120;
	wire new_net_6627;
	wire new_net_7501;
	wire new_net_7525;
	wire new_net_4050;
	wire new_net_5824;
	wire new_net_939;
	wire new_net_1809;
	wire new_net_2186;
	wire new_net_1848;
	wire new_net_48;
	wire _0666_;
	wire _0162_;
	wire _1170_;
	wire new_net_2291;
	wire new_net_4251;
	wire new_net_5248;
	wire new_net_6440;
	wire new_net_7398;
	wire new_net_5342;
	wire new_net_4553;
	wire new_net_195;
	wire new_net_2409;
	wire new_net_8022;
	wire new_net_6701;
	wire new_net_3330;
	wire new_net_1921;
	wire new_net_484;
	wire new_net_517;
	wire new_net_868;
	wire new_net_1015;
	wire new_net_5850;
	wire new_net_5929;
	wire new_net_6880;
	wire new_net_7375;
	wire new_net_7826;
	wire new_net_6873;
	wire new_net_5844;
	wire _0766_;
	wire new_net_4311;
	wire new_net_1405;
	wire new_net_1976;
	wire new_net_695;
	wire new_net_977;
	wire new_net_767;
	wire new_net_1051;
	wire _1171_;
	wire _0667_;
	wire _0163_;
	wire new_net_551;
	wire new_net_6613;
	wire new_net_1985;
	wire new_net_2740;
	wire new_net_3275;
	wire new_net_3165;
	wire new_net_156;
	wire new_net_1121;
	wire new_net_1157;
	wire new_net_4145;
	wire new_net_4686;
	wire new_net_4983;
	wire new_net_6122;
	wire new_net_5059;
	wire new_net_3093;
	wire new_net_5057;
	wire new_net_5720;
	wire new_net_5604;
	wire new_net_7669;
	wire new_net_658;
	wire new_net_940;
	wire new_net_2503;
	wire new_net_3021;
	wire _1172_;
	wire _0164_;
	wire _0668_;
	wire new_net_49;
	wire new_net_2323;
	wire new_net_4375;
	wire new_net_7296;
	wire new_net_7914;
	wire new_net_7052;
	wire new_net_6974;
	wire new_net_7640;
	wire new_net_7224;
	wire new_net_1192;
	wire new_net_122;
	wire new_net_398;
	wire new_net_485;
	wire new_net_518;
	wire new_net_1016;
	wire new_net_2755;
	wire new_net_4485;
	wire new_net_4508;
	wire new_net_4949;
	wire new_net_7139;
	wire new_net_6650;
	wire new_net_6829;
	wire new_net_2727;
	wire new_net_3666;
	wire new_net_1;
	wire new_net_3178;
	wire new_net_768;
	wire new_net_1052;
	wire _0669_;
	wire _1173_;
	wire _0165_;
	wire new_net_552;
	wire new_net_5101;
	wire new_net_7163;
	wire new_net_6389;
	wire new_net_6382;
	wire new_net_6304;
	wire new_net_1158;
	wire new_net_2862;
	wire new_net_1831;
	wire new_net_3022;
	wire new_net_2007;
	wire new_net_157;
	wire new_net_3166;
	wire new_net_4159;
	wire _0019_;
	wire new_net_4582;
	wire new_net_2649;
	wire new_net_8013;
	wire new_net_6321;
	wire new_net_869;
	wire new_net_659;
	wire new_net_941;
	wire new_net_2187;
	wire new_net_1895;
	wire _0670_;
	wire _1174_;
	wire _0166_;
	wire new_net_2292;
	wire new_net_5851;
	wire new_net_7817;
	wire new_net_1659;
	wire new_net_4771;
	wire new_net_6176;
	wire new_net_6343;
	wire new_net_1193;
	wire new_net_1406;
	wire new_net_3290;
	wire new_net_978;
	wire new_net_123;
	wire new_net_399;
	wire new_net_486;
	wire new_net_519;
	wire new_net_696;
	wire new_net_4564;
	wire new_net_5522;
	wire new_net_6593;
	wire new_net_6104;
	wire new_net_8122;
	wire new_net_4276;
	wire new_net_6102;
	wire new_net_1724;
	wire new_net_1854;
	wire new_net_2741;
	wire new_net_3276;
	wire _1175_;
	wire _0671_;
	wire _0167_;
	wire new_net_769;
	wire new_net_4146;
	wire new_net_4989;
	wire new_net_7276;
	wire new_net_7488;
	wire new_net_5595;
	wire new_net_6452;
	wire new_net_1958;
	wire new_net_2863;
	wire new_net_3331;
	wire new_net_50;
	wire new_net_4376;
	wire new_net_4825;
	wire new_net_5484;
	wire new_net_5685;
	wire new_net_8014;
	wire new_net_8263;
	wire new_net_7593;
	wire new_net_8244;
	wire new_net_4129;
	wire new_net_7208;
	wire new_net_870;
	wire new_net_2324;
	wire new_net_660;
	wire new_net_942;
	wire new_net_1017;
	wire _1176_;
	wire _0767_;
	wire _0672_;
	wire _0168_;
	wire new_net_4486;
	wire new_net_6063;
	wire new_net_5159;
	wire new_net_7849;
	wire _0244_;
	wire new_net_2054;
	wire new_net_1407;
	wire new_net_3667;
	wire new_net_124;
	wire new_net_400;
	wire new_net_520;
	wire new_net_553;
	wire new_net_697;
	wire new_net_979;
	wire new_net_1053;
	wire new_net_7031;
	wire new_net_7697;
	wire new_net_2604;
	wire new_net_6290;
	wire new_net_7864;
	wire new_net_3167;
	wire new_net_1123;
	wire new_net_1159;
	wire new_net_158;
	wire new_net_3023;
	wire _0169_;
	wire _0673_;
	wire _1177_;
	wire new_net_5234;
	wire new_net_5507;
	wire new_net_6140;
	wire new_net_5493;
	wire new_net_6935;
	wire new_net_6548;
	wire new_net_1949;
	wire new_net_3309;
	wire new_net_51;
	wire new_net_3179;
	wire new_net_5852;
	wire new_net_5931;
	wire new_net_7377;
	wire new_net_8176;
	wire new_net_4840;
	wire new_net_7975;
	wire new_net_6162;
	wire new_net_2443;
	wire new_net_2293;
	wire new_net_1194;
	wire new_net_661;
	wire new_net_943;
	wire _0170_;
	wire _0674_;
	wire _1178_;
	wire new_net_1018;
	wire new_net_2188;
	wire new_net_487;
	wire new_net_2159;
	wire new_net_125;
	wire new_net_554;
	wire new_net_770;
	wire new_net_980;
	wire new_net_1054;
	wire new_net_3248;
	wire new_net_4147;
	wire new_net_4243;
	wire new_net_5257;
	wire new_net_5384;
	wire new_net_4242;
	wire new_net_2872;
	wire new_net_5414;
	wire new_net_7262;
	wire new_net_3393;
	wire new_net_7479;
	wire new_net_4543;
	wire new_net_7651;
	wire new_net_1124;
	wire new_net_1160;
	wire new_net_159;
	wire new_net_2864;
	wire new_net_3291;
	wire _1179_;
	wire _0171_;
	wire _0675_;
	wire new_net_2505;
	wire new_net_3332;
	wire _0416_;
	wire new_net_7584;
	wire new_net_8230;
	wire new_net_3850;
	wire new_net_6427;
	wire new_net_52;
	wire new_net_871;
	wire new_net_1776;
	wire new_net_3310;
	wire new_net_4160;
	wire new_net_4487;
	wire new_net_4510;
	wire new_net_2221;
	wire new_net_4951;
	wire new_net_5361;
	wire new_net_5407;
	wire new_net_7429;
	wire new_net_7601;
	wire new_net_8252;
	wire new_net_6407;
	wire new_net_6199;
	wire new_net_488;
	wire new_net_521;
	wire new_net_2325;
	wire new_net_1195;
	wire new_net_1408;
	wire new_net_3668;
	wire new_net_401;
	wire new_net_662;
	wire new_net_944;
	wire _0172_;
	wire new_net_4252;
	wire new_net_6732;
	wire new_net_8051;
	wire _0384_;
	wire new_net_7022;
	wire new_net_4170;
	wire new_net_8147;
	wire new_net_4658;
	wire new_net_7194;
	wire new_net_16;
	wire new_net_126;
	wire new_net_555;
	wire new_net_771;
	wire new_net_981;
	wire new_net_1055;
	wire new_net_3024;
	wire new_net_5235;
	wire new_net_5508;
	wire new_net_5709;
	wire new_net_5272;
	wire new_net_6136;
	wire new_net_6754;
	wire new_net_5729;
	wire new_net_6926;
	wire new_net_1125;
	wire new_net_160;
	wire _0173_;
	wire _1181_;
	wire _0677_;
	wire new_net_3180;
	wire new_net_5829;
	wire new_net_5853;
	wire new_net_5932;
	wire new_net_6475;
	wire new_net_7923;
	wire new_net_7843;
	wire new_net_7727;
	wire new_net_5506;
	wire _0245_;
	wire new_net_1813;
	wire new_net_1867;
	wire new_net_2028;
	wire new_net_53;
	wire new_net_872;
	wire new_net_4566;
	wire new_net_4584;
	wire new_net_6076;
	wire new_net_596;
	wire new_net_2599;
	wire new_net_6948;
	wire new_net_7448;
	wire new_net_682;
	wire new_net_5802;
	wire new_net_4338;
	wire new_net_1020;
	wire new_net_2189;
	wire new_net_1864;
	wire new_net_522;
	wire new_net_2294;
	wire new_net_1863;
	wire new_net_1196;
	wire new_net_1409;
	wire new_net_402;
	wire new_net_663;
	wire new_net_5768;
	wire new_net_6630;
	wire new_net_6637;
	wire new_net_7253;
	wire new_net_3816;
	wire new_net_7470;
	wire new_net_5083;
	wire new_net_6313;
	wire new_net_3292;
	wire new_net_3333;
	wire new_net_2080;
	wire new_net_1161;
	wire new_net_1963;
	wire new_net_2865;
	wire new_net_556;
	wire new_net_772;
	wire new_net_982;
	wire new_net_4378;
	wire new_net_7570;
	wire new_net_463;
	wire new_net_4892;
	wire new_net_7775;
	wire new_net_7069;
	wire new_net_1126;
	wire _1183_;
	wire new_net_1787;
	wire _0175_;
	wire _0679_;
	wire new_net_3311;
	wire new_net_4488;
	wire new_net_4511;
	wire new_net_5143;
	wire new_net_5362;
	wire new_net_6094;
	wire new_net_8194;
	wire new_net_5442;
	wire new_net_1816;
	wire new_net_54;
	wire new_net_489;
	wire new_net_873;
	wire new_net_1802;
	wire new_net_4601;
	wire new_net_6631;
	wire new_net_3779;
	wire new_net_7091;
	wire new_net_7402;
	wire new_net_8042;
	wire new_net_4164;
	wire new_net_6602;
	wire new_net_6895;
	wire _0940_;
	wire new_net_322;
	wire new_net_2973;
	wire new_net_700;
	wire new_net_3025;
	wire new_net_1021;
	wire new_net_1056;
	wire new_net_2081;
	wire new_net_127;
	wire new_net_2326;
	wire new_net_1197;
	wire _1184_;
	wire _0176_;
	wire new_net_1374;
	wire new_net_8265;
	wire new_net_1660;
	wire new_net_3192;
	wire new_net_8085;
	wire new_net_5352;
	wire new_net_3181;
	wire new_net_1785;
	wire new_net_1162;
	wire new_net_161;
	wire new_net_557;
	wire new_net_983;
	wire new_net_4824;
	wire new_net_5830;
	wire new_net_5854;
	wire new_net_5933;
	wire _0177_;
	wire _1185_;
	wire new_net_2742;
	wire _0681_;
	wire new_net_4567;
	wire new_net_5687;
	wire new_net_6077;
	wire new_net_6228;
	wire new_net_6903;
	wire new_net_7171;
	wire new_net_6367;
	wire new_net_3507;
	wire new_net_2413;
	wire new_net_3168;
	wire new_net_403;
	wire new_net_490;
	wire new_net_523;
	wire new_net_874;
	wire new_net_1410;
	wire new_net_4991;
	wire new_net_5259;
	wire new_net_5386;
	wire new_net_5465;
	wire new_net_4080;
	wire new_net_7040;
	wire new_net_2897;
	wire new_net_6967;
	wire new_net_4953;
	wire new_net_665;
	wire new_net_947;
	wire new_net_2190;
	wire new_net_2507;
	wire new_net_3334;
	wire new_net_773;
	wire new_net_1057;
	wire new_net_2295;
	wire new_net_128;
	wire _0682_;
	wire new_net_230;
	wire new_net_2246;
	wire new_net_5987;
	wire new_net_7306;
	wire new_net_8214;
	wire new_net_2783;
	wire new_net_3827;
	wire new_net_6036;
	wire new_net_3312;
	wire new_net_1127;
	wire new_net_162;
	wire new_net_984;
	wire new_net_3277;
	wire new_net_4489;
	wire new_net_4512;
	wire new_net_5363;
	wire new_net_5808;
	wire new_net_6550;
	wire new_net_8185;
	wire new_net_5913;
	wire new_net_2605;
	wire new_net_3169;
	wire _0683_;
	wire new_net_55;
	wire _1187_;
	wire _0179_;
	wire new_net_4602;
	wire new_net_6632;
	wire new_net_7403;
	wire new_net_7506;
	wire new_net_7530;
	wire new_net_8001;
	wire new_net_3144;
	wire new_net_2178;
	wire new_net_3026;
	wire new_net_404;
	wire new_net_524;
	wire new_net_701;
	wire new_net_875;
	wire new_net_1022;
	wire new_net_1198;
	wire new_net_1411;
	wire new_net_5237;
	wire new_net_5510;
	wire new_net_5825;
	wire new_net_6859;
	wire new_net_7399;
	wire new_net_5249;
	wire new_net_6441;
	wire new_net_8023;
	wire new_net_3278;
	wire new_net_948;
	wire new_net_666;
	wire new_net_774;
	wire new_net_558;
	wire _1188_;
	wire _0180_;
	wire _0684_;
	wire new_net_2327;
	wire new_net_5831;
	wire new_net_5847;
	wire new_net_6881;
	wire new_net_7827;
	wire new_net_6186;
	wire new_net_7510;
	wire new_net_1896;
	wire new_net_985;
	wire new_net_1128;
	wire new_net_2479;
	wire new_net_4161;
	wire new_net_4381;
	wire new_net_4568;
	wire new_net_6078;
	wire new_net_6229;
	wire new_net_6904;
	wire new_net_7508;
	wire new_net_2240;
	wire _0941_;
	wire new_net_491;
	wire new_net_17;
	wire _1189_;
	wire _0181_;
	wire _0685_;
	wire new_net_738;
	wire new_net_4992;
	wire new_net_5260;
	wire new_net_5387;
	wire new_net_5466;
	wire new_net_6614;
	wire new_net_1664;
	wire new_net_2987;
	wire new_net_545;
	wire new_net_6542;
	wire new_net_5605;
	wire new_net_2867;
	wire new_net_3335;
	wire new_net_129;
	wire new_net_702;
	wire new_net_876;
	wire new_net_1023;
	wire new_net_1058;
	wire new_net_1199;
	wire new_net_4227;
	wire new_net_4829;
	wire new_net_7297;
	wire new_net_7915;
	wire new_net_4380;
	wire new_net_7053;
	wire new_net_4757;
	wire new_net_6975;
	wire new_net_5738;
	wire new_net_1164;
	wire new_net_163;
	wire new_net_667;
	wire new_net_3313;
	wire new_net_2191;
	wire new_net_559;
	wire new_net_2296;
	wire _0686_;
	wire _1190_;
	wire _0182_;
	wire new_net_5660;
	wire new_net_7140;
	wire new_net_6073;
	wire _0386_;
	wire new_net_6651;
	wire _0695_;
	wire new_net_197;
	wire new_net_2728;
	wire new_net_3170;
	wire new_net_986;
	wire new_net_4585;
	wire new_net_6633;
	wire new_net_7404;
	wire new_net_7507;
	wire new_net_7531;
	wire new_net_7943;
	wire new_net_1252;
	wire new_net_5102;
	wire new_net_5314;
	wire new_net_1871;
	wire new_net_6383;
	wire new_net_1412;
	wire new_net_405;
	wire new_net_3027;
	wire new_net_492;
	wire new_net_57;
	wire new_net_525;
	wire _0687_;
	wire _0183_;
	wire _1191_;
	wire new_net_4149;
	wire new_net_7390;
	wire new_net_4022;
	wire new_net_6405;
	wire new_net_1200;
	wire new_net_1964;
	wire new_net_3279;
	wire new_net_1775;
	wire new_net_1059;
	wire _0247_;
	wire new_net_130;
	wire new_net_775;
	wire new_net_877;
	wire new_net_949;
	wire new_net_7818;
	wire new_net_560;
	wire new_net_1129;
	wire new_net_1165;
	wire new_net_2328;
	wire new_net_2729;
	wire new_net_164;
	wire new_net_668;
	wire _1192_;
	wire _0688_;
	wire _0184_;
	wire _0590_;
	wire new_net_1542;
	wire new_net_5523;
	wire new_net_6344;
	wire new_net_5938;
	wire new_net_6594;
	wire new_net_8125;
	wire new_net_6105;
	wire new_net_6103;
	wire new_net_2743;
	wire new_net_987;
	wire new_net_4993;
	wire new_net_5261;
	wire new_net_5388;
	wire new_net_5467;
	wire new_net_5589;
	wire new_net_6951;
	wire new_net_7612;
	wire new_net_7277;
	wire new_net_464;
	wire new_net_7489;
	wire _0974_;
	wire new_net_6455;
	wire new_net_5596;
	wire new_net_1413;
	wire new_net_2868;
	wire _0689_;
	wire new_net_406;
	wire new_net_703;
	wire new_net_1024;
	wire new_net_2509;
	wire new_net_3336;
	wire _1193_;
	wire _0185_;
	wire new_net_2633;
	wire new_net_7594;
	wire new_net_7632;
	wire new_net_8245;
	wire new_net_2051;
	wire new_net_1201;
	wire new_net_3314;
	wire new_net_776;
	wire new_net_878;
	wire new_net_950;
	wire new_net_4491;
	wire new_net_4514;
	wire new_net_5365;
	wire new_net_5810;
	wire new_net_6131;
	wire new_net_7799;
	wire new_net_7850;
	wire _0942_;
	wire new_net_2059;
	wire new_net_561;
	wire new_net_1130;
	wire new_net_2297;
	wire new_net_1166;
	wire new_net_1757;
	wire new_net_2744;
	wire new_net_669;
	wire new_net_2040;
	wire new_net_3171;
	wire new_net_1375;
	wire new_net_3408;
	wire new_net_7894;
	wire new_net_526;
	wire new_net_7032;
	wire new_net_7698;
	wire new_net_4180;
	wire new_net_6291;
	wire new_net_7865;
	wire new_net_3028;
	wire new_net_3182;
	wire new_net_58;
	wire new_net_493;
	wire new_net_988;
	wire new_net_5239;
	wire new_net_5512;
	wire new_net_5689;
	wire new_net_5732;
	wire new_net_6230;
	wire new_net_7376;
	wire new_net_7956;
	wire new_net_5688;
	wire new_net_6141;
	wire new_net_2363;
	wire new_net_6023;
	wire new_net_131;
	wire new_net_1414;
	wire new_net_2033;
	wire new_net_3280;
	wire new_net_407;
	wire new_net_704;
	wire new_net_1025;
	wire new_net_1060;
	wire _0691_;
	wire _1195_;
	wire new_net_8003;
	wire new_net_1439;
	wire _0696_;
	wire new_net_1202;
	wire new_net_1870;
	wire new_net_18;
	wire new_net_165;
	wire new_net_879;
	wire new_net_4570;
	wire new_net_6080;
	wire new_net_6906;
	wire new_net_7174;
	wire new_net_7301;
	wire _1146_;
	wire new_net_2072;
	wire new_net_2962;
	wire new_net_2166;
	wire new_net_1167;
	wire new_net_2329;
	wire new_net_670;
	wire _1196_;
	wire _0692_;
	wire _0188_;
	wire new_net_4603;
	wire new_net_4768;
	wire new_net_4994;
	wire new_net_5262;
	wire _0771_;
	wire new_net_231;
	wire new_net_1286;
	wire new_net_2873;
	wire new_net_5415;
	wire new_net_7263;
	wire new_net_7480;
	wire new_net_938;
	wire new_net_3337;
	wire new_net_2869;
	wire new_net_3183;
	wire new_net_59;
	wire _0248_;
	wire new_net_494;
	wire new_net_527;
	wire new_net_989;
	wire new_net_4163;
	wire new_net_4217;
	wire new_net_7652;
	wire new_net_1731;
	wire new_net_3600;
	wire new_net_3126;
	wire new_net_7585;
	wire new_net_8231;
	wire new_net_3851;
	wire new_net_777;
	wire new_net_1061;
	wire new_net_132;
	wire new_net_1415;
	wire new_net_951;
	wire _1197_;
	wire _0693_;
	wire _0189_;
	wire _0591_;
	wire new_net_3771;
	wire new_net_6428;
	wire new_net_6807;
	wire new_net_7430;
	wire new_net_7602;
	wire new_net_166;
	wire new_net_562;
	wire new_net_880;
	wire new_net_1131;
	wire new_net_5711;
	wire new_net_6635;
	wire new_net_7406;
	wire new_net_7509;
	wire new_net_8253;
	wire new_net_2259;
	wire new_net_6733;
	wire new_net_7023;
	wire new_net_8148;
	wire _0975_;
	input G1;
	input G10;
	input G100;
	input G101;
	input G102;
	input G103;
	input G104;
	input G105;
	input G106;
	input G107;
	input G108;
	input G109;
	input G11;
	input G110;
	input G111;
	input G112;
	input G113;
	input G114;
	input G115;
	input G116;
	input G117;
	input G118;
	input G119;
	input G12;
	input G120;
	input G121;
	input G122;
	input G123;
	input G124;
	input G125;
	input G126;
	input G127;
	input G128;
	input G129;
	input G13;
	input G130;
	input G131;
	input G132;
	input G133;
	input G134;
	input G135;
	input G136;
	input G137;
	input G138;
	input G139;
	input G14;
	input G140;
	input G141;
	input G142;
	input G143;
	input G144;
	input G145;
	input G146;
	input G147;
	input G148;
	input G149;
	input G15;
	input G150;
	input G151;
	input G152;
	input G153;
	input G154;
	input G155;
	input G156;
	input G157;
	input G158;
	input G159;
	input G16;
	input G160;
	input G161;
	input G162;
	input G163;
	input G164;
	input G165;
	input G166;
	input G167;
	input G168;
	input G169;
	input G17;
	input G170;
	input G171;
	input G172;
	input G173;
	input G174;
	input G175;
	input G176;
	input G177;
	input G178;
	input G18;
	input G19;
	input G2;
	input G20;
	input G21;
	input G22;
	input G23;
	input G24;
	input G25;
	input G26;
	input G27;
	input G28;
	input G29;
	input G3;
	input G30;
	input G31;
	input G32;
	input G33;
	input G34;
	input G35;
	input G36;
	input G37;
	input G38;
	input G39;
	input G4;
	input G40;
	input G41;
	input G42;
	input G43;
	input G44;
	input G45;
	input G46;
	input G47;
	input G48;
	input G49;
	input G5;
	input G50;
	input G51;
	input G52;
	input G53;
	input G54;
	input G55;
	input G56;
	input G57;
	input G58;
	input G59;
	input G6;
	input G60;
	input G61;
	input G62;
	input G63;
	input G64;
	input G65;
	input G66;
	input G67;
	input G68;
	input G69;
	input G7;
	input G70;
	input G71;
	input G72;
	input G73;
	input G74;
	input G75;
	input G76;
	input G77;
	input G78;
	input G79;
	input G8;
	input G80;
	input G81;
	input G82;
	input G83;
	input G84;
	input G85;
	input G86;
	input G87;
	input G88;
	input G89;
	input G9;
	input G90;
	input G91;
	input G92;
	input G93;
	input G94;
	input G95;
	input G96;
	input G97;
	input G98;
	input G99;
	output G5193;
	output G5194;
	output G5195;
	output G5196;
	output G5197;
	output G5198;
	output G5199;
	output G5200;
	output G5201;
	output G5202;
	output G5203;
	output G5204;
	output G5205;
	output G5206;
	output G5207;
	output G5208;
	output G5209;
	output G5210;
	output G5211;
	output G5212;
	output G5213;
	output G5214;
	output G5215;
	output G5216;
	output G5217;
	output G5218;
	output G5219;
	output G5220;
	output G5221;
	output G5222;
	output G5223;
	output G5224;
	output G5225;
	output G5226;
	output G5227;
	output G5228;
	output G5229;
	output G5230;
	output G5231;
	output G5232;
	output G5233;
	output G5234;
	output G5235;
	output G5236;
	output G5237;
	output G5238;
	output G5239;
	output G5240;
	output G5241;
	output G5242;
	output G5243;
	output G5244;
	output G5245;
	output G5246;
	output G5247;
	output G5248;
	output G5249;
	output G5250;
	output G5251;
	output G5252;
	output G5253;
	output G5254;
	output G5255;
	output G5256;
	output G5257;
	output G5258;
	output G5259;
	output G5260;
	output G5261;
	output G5262;
	output G5263;
	output G5264;
	output G5265;
	output G5266;
	output G5267;
	output G5268;
	output G5269;
	output G5270;
	output G5271;
	output G5272;
	output G5273;
	output G5274;
	output G5275;
	output G5276;
	output G5277;
	output G5278;
	output G5279;
	output G5280;
	output G5281;
	output G5282;
	output G5283;
	output G5284;
	output G5285;
	output G5286;
	output G5287;
	output G5288;
	output G5289;
	output G5290;
	output G5291;
	output G5292;
	output G5293;
	output G5294;
	output G5295;
	output G5296;
	output G5297;
	output G5298;
	output G5299;
	output G5300;
	output G5301;
	output G5302;
	output G5303;
	output G5304;
	output G5305;
	output G5306;
	output G5307;
	output G5308;
	output G5309;
	output G5310;
	output G5311;
	output G5312;
	output G5313;
	output G5314;
	output G5315;

	and_bb _1248_ (
		.a(new_net_1633),
		.b(new_net_1523),
		.c(_0578_)
	);

	and_bi _1249_ (
		.a(new_net_1337),
		.b(new_net_1530),
		.c(_0579_)
	);

	and_ii _1250_ (
		.a(_0579_),
		.b(_0578_),
		.c(_0580_)
	);

	and_bb _1251_ (
		.a(new_net_175),
		.b(new_net_1518),
		.c(_0581_)
	);

	and_bi _1252_ (
		.a(new_net_2107),
		.b(new_net_1524),
		.c(_0582_)
	);

	and_ii _1253_ (
		.a(_0582_),
		.b(_0581_),
		.c(_0583_)
	);

	or_ii _1254_ (
		.a(new_net_305),
		.b(new_net_243),
		.c(_0584_)
	);

	and_ii _1255_ (
		.a(new_net_309),
		.b(new_net_249),
		.c(_0585_)
	);

	and_bi _1256_ (
		.a(new_net_329),
		.b(new_net_2108),
		.c(new_net_1)
	);

	inv _1257_ (
		.din(new_net_1277),
		.dout(new_net_2379)
	);

	inv _1258_ (
		.din(new_net_1634),
		.dout(new_net_2487)
	);

	inv _1259_ (
		.din(new_net_1626),
		.dout(new_net_2415)
	);

	inv _1260_ (
		.din(G151),
		.dout(new_net_24)
	);

	inv _1261_ (
		.din(new_net_1624),
		.dout(new_net_2359)
	);

	inv _1262_ (
		.din(new_net_847),
		.dout(new_net_2463)
	);

	inv _1263_ (
		.din(new_net_1340),
		.dout(new_net_2429)
	);

	inv _1264_ (
		.din(new_net_1260),
		.dout(new_net_2)
	);

	inv _1265_ (
		.din(new_net_1707),
		.dout(new_net_2465)
	);

	inv _1266_ (
		.din(new_net_1439),
		.dout(new_net_2441)
	);

	inv _1267_ (
		.din(new_net_208),
		.dout(new_net_2403)
	);

	inv _1268_ (
		.din(new_net_1404),
		.dout(new_net_2419)
	);

	inv _1269_ (
		.din(new_net_1400),
		.dout(new_net_2375)
	);

	or_bi _1270_ (
		.a(new_net_2109),
		.b(new_net_1271),
		.c(new_net_2389)
	);

	or_ii _1271_ (
		.a(G154),
		.b(G136),
		.c(new_net_13)
	);

	or_ii _1272_ (
		.a(new_net_1272),
		.b(new_net_2110),
		.c(new_net_0)
	);

	or_bi _1273_ (
		.a(new_net_914),
		.b(new_net_2111),
		.c(new_net_2351)
	);

	inv _1274_ (
		.din(new_net_55),
		.dout(new_net_25)
	);

	inv _1275_ (
		.din(new_net_1338),
		.dout(new_net_26)
	);

	or_ii _1276_ (
		.a(new_net_2112),
		.b(new_net_1304),
		.c(_0586_)
	);

	and_bi _1277_ (
		.a(new_net_2113),
		.b(new_net_1310),
		.c(_0587_)
	);

	and_bi _1278_ (
		.a(_0586_),
		.b(_0587_),
		.c(_0588_)
	);

	or_bb _1279_ (
		.a(new_net_2114),
		.b(new_net_913),
		.c(new_net_2507)
	);

	or_ii _1280_ (
		.a(new_net_2115),
		.b(new_net_1305),
		.c(_0589_)
	);

	and_bi _1281_ (
		.a(new_net_2116),
		.b(new_net_1311),
		.c(_0590_)
	);

	and_bi _1282_ (
		.a(_0589_),
		.b(_0590_),
		.c(_0591_)
	);

	or_bb _1283_ (
		.a(new_net_2117),
		.b(new_net_912),
		.c(new_net_27)
	);

	or_bi _1284_ (
		.a(new_net_908),
		.b(new_net_2118),
		.c(new_net_2495)
	);

	or_bi _1285_ (
		.a(new_net_220),
		.b(new_net_1230),
		.c(_0592_)
	);

	and_bi _1286_ (
		.a(new_net_2119),
		.b(new_net_93),
		.c(_0593_)
	);

	and_bb _1287_ (
		.a(new_net_1032),
		.b(new_net_1529),
		.c(_0594_)
	);

	and_bi _1288_ (
		.a(new_net_848),
		.b(new_net_1515),
		.c(_0595_)
	);

	and_ii _1289_ (
		.a(_0595_),
		.b(_0594_),
		.c(_0596_)
	);

	or_bb _1290_ (
		.a(new_net_553),
		.b(new_net_331),
		.c(_0597_)
	);

	and_bb _1291_ (
		.a(new_net_556),
		.b(new_net_332),
		.c(_0598_)
	);

	and_bi _1292_ (
		.a(_0597_),
		.b(_0598_),
		.c(_0599_)
	);

	or_bb _1293_ (
		.a(new_net_718),
		.b(new_net_1231),
		.c(_0600_)
	);

	inv _1294_ (
		.din(new_net_221),
		.dout(_0601_)
	);

	and_ii _1295_ (
		.a(new_net_1033),
		.b(new_net_982),
		.c(_0602_)
	);

	and_bi _1296_ (
		.a(new_net_1031),
		.b(new_net_1007),
		.c(_0603_)
	);

	and_ii _1297_ (
		.a(_0603_),
		.b(_0602_),
		.c(_0604_)
	);

	and_bi _1298_ (
		.a(new_net_1233),
		.b(new_net_686),
		.c(_0605_)
	);

	or_bb _1299_ (
		.a(_0605_),
		.b(new_net_614),
		.c(_0606_)
	);

	and_bi _1300_ (
		.a(_0600_),
		.b(new_net_2120),
		.c(_0607_)
	);

	and_ii _1301_ (
		.a(_0607_),
		.b(new_net_2121),
		.c(new_net_4)
	);

	and_bi _1302_ (
		.a(new_net_2122),
		.b(new_net_84),
		.c(_0608_)
	);

	inv _1303_ (
		.din(new_net_557),
		.dout(_0609_)
	);

	or_ii _1304_ (
		.a(new_net_1655),
		.b(new_net_1516),
		.c(_0610_)
	);

	and_bi _1305_ (
		.a(new_net_1708),
		.b(new_net_1519),
		.c(_0611_)
	);

	and_bi _1306_ (
		.a(_0610_),
		.b(new_net_2123),
		.c(_0612_)
	);

	and_bi _1307_ (
		.a(new_net_1591),
		.b(new_net_61),
		.c(_0613_)
	);

	inv _1308_ (
		.din(new_net_1592),
		.dout(_0614_)
	);

	or_ii _1309_ (
		.a(new_net_63),
		.b(new_net_131),
		.c(_0615_)
	);

	and_bi _1310_ (
		.a(new_net_1711),
		.b(new_net_1431),
		.c(_0616_)
	);

	and_bi _1311_ (
		.a(new_net_104),
		.b(_0616_),
		.c(_0617_)
	);

	and_bi _1312_ (
		.a(new_net_554),
		.b(new_net_1434),
		.c(_0618_)
	);

	and_bb _1313_ (
		.a(new_net_191),
		.b(new_net_1713),
		.c(_0619_)
	);

	or_bb _1314_ (
		.a(new_net_398),
		.b(new_net_2124),
		.c(_0620_)
	);

	or_bb _1315_ (
		.a(new_net_216),
		.b(new_net_1213),
		.c(_0621_)
	);

	or_bb _1316_ (
		.a(new_net_1657),
		.b(new_net_456),
		.c(_0622_)
	);

	and_bi _1317_ (
		.a(new_net_1662),
		.b(new_net_342),
		.c(_0623_)
	);

	and_bi _1318_ (
		.a(_0622_),
		.b(_0623_),
		.c(_0624_)
	);

	or_bb _1319_ (
		.a(_0624_),
		.b(new_net_134),
		.c(_0625_)
	);

	or_ii _1320_ (
		.a(new_net_1688),
		.b(new_net_1656),
		.c(_0626_)
	);

	and_bi _1321_ (
		.a(new_net_1674),
		.b(new_net_1661),
		.c(_0627_)
	);

	and_bi _1322_ (
		.a(_0626_),
		.b(_0627_),
		.c(_0628_)
	);

	and_bi _1323_ (
		.a(new_net_133),
		.b(_0628_),
		.c(_0629_)
	);

	and_bi _1324_ (
		.a(_0625_),
		.b(_0629_),
		.c(_0630_)
	);

	and_bi _1325_ (
		.a(new_net_1214),
		.b(new_net_442),
		.c(_0631_)
	);

	or_bb _1326_ (
		.a(_0631_),
		.b(new_net_610),
		.c(_0632_)
	);

	and_bi _1327_ (
		.a(_0621_),
		.b(new_net_2125),
		.c(_0633_)
	);

	and_ii _1328_ (
		.a(_0633_),
		.b(new_net_2126),
		.c(new_net_12)
	);

	and_bi _1329_ (
		.a(new_net_2127),
		.b(new_net_101),
		.c(_0634_)
	);

	or_ii _1330_ (
		.a(new_net_1555),
		.b(new_net_1243),
		.c(_0635_)
	);

	and_bi _1331_ (
		.a(new_net_2128),
		.b(new_net_1553),
		.c(_0636_)
	);

	and_bi _1332_ (
		.a(_0635_),
		.b(new_net_2129),
		.c(_0637_)
	);

	and_bi _1333_ (
		.a(new_net_898),
		.b(new_net_536),
		.c(_0638_)
	);

	and_bi _1334_ (
		.a(new_net_539),
		.b(new_net_899),
		.c(_0639_)
	);

	or_bb _1335_ (
		.a(new_net_640),
		.b(new_net_558),
		.c(_0640_)
	);

	and_bi _1336_ (
		.a(new_net_50),
		.b(new_net_720),
		.c(_0641_)
	);

	and_bi _1337_ (
		.a(new_net_724),
		.b(new_net_53),
		.c(_0642_)
	);

	and_ii _1338_ (
		.a(new_net_2130),
		.b(new_net_818),
		.c(_0643_)
	);

	or_bb _1339_ (
		.a(new_net_1026),
		.b(new_net_1215),
		.c(_0644_)
	);

	inv _1340_ (
		.din(new_net_900),
		.dout(_0645_)
	);

	or_bb _1341_ (
		.a(new_net_1250),
		.b(new_net_462),
		.c(_0646_)
	);

	and_bi _1342_ (
		.a(new_net_1245),
		.b(new_net_335),
		.c(_0647_)
	);

	and_bi _1343_ (
		.a(_0646_),
		.b(_0647_),
		.c(_0648_)
	);

	or_bb _1344_ (
		.a(_0648_),
		.b(new_net_1290),
		.c(_0649_)
	);

	or_ii _1345_ (
		.a(new_net_1694),
		.b(new_net_1249),
		.c(_0650_)
	);

	and_bi _1346_ (
		.a(new_net_1667),
		.b(new_net_1244),
		.c(_0651_)
	);

	and_bi _1347_ (
		.a(_0650_),
		.b(_0651_),
		.c(_0652_)
	);

	and_bi _1348_ (
		.a(new_net_1293),
		.b(_0652_),
		.c(_0653_)
	);

	and_bi _1349_ (
		.a(_0649_),
		.b(_0653_),
		.c(_0654_)
	);

	and_bi _1350_ (
		.a(new_net_1203),
		.b(new_net_845),
		.c(_0655_)
	);

	or_bb _1351_ (
		.a(_0655_),
		.b(new_net_623),
		.c(_0656_)
	);

	and_bi _1352_ (
		.a(_0644_),
		.b(new_net_2131),
		.c(_0657_)
	);

	and_ii _1353_ (
		.a(_0657_),
		.b(new_net_2132),
		.c(new_net_3)
	);

	and_bi _1354_ (
		.a(new_net_2133),
		.b(new_net_94),
		.c(_0658_)
	);

	and_ii _1355_ (
		.a(new_net_1261),
		.b(new_net_1531),
		.c(_0659_)
	);

	and_bi _1356_ (
		.a(new_net_1265),
		.b(new_net_1119),
		.c(_0660_)
	);

	and_bi _1357_ (
		.a(new_net_1121),
		.b(new_net_1268),
		.c(_0661_)
	);

	and_ii _1358_ (
		.a(new_net_1345),
		.b(new_net_923),
		.c(_0662_)
	);

	inv _1359_ (
		.din(new_net_1288),
		.dout(_0663_)
	);

	and_bb _1360_ (
		.a(new_net_1602),
		.b(new_net_1525),
		.c(_0664_)
	);

	and_bi _1361_ (
		.a(new_net_1625),
		.b(new_net_1527),
		.c(_0665_)
	);

	or_bb _1362_ (
		.a(_0665_),
		.b(_0664_),
		.c(_0666_)
	);

	and_bi _1363_ (
		.a(new_net_1090),
		.b(new_net_1020),
		.c(_0667_)
	);

	and_bi _1364_ (
		.a(new_net_1019),
		.b(new_net_1091),
		.c(_0668_)
	);

	and_ii _1365_ (
		.a(new_net_370),
		.b(new_net_1103),
		.c(_0669_)
	);

	inv _1366_ (
		.din(new_net_1180),
		.dout(_0670_)
	);

	or_bi _1367_ (
		.a(new_net_1192),
		.b(new_net_400),
		.c(_0671_)
	);

	and_bi _1368_ (
		.a(new_net_973),
		.b(new_net_608),
		.c(_0672_)
	);

	inv _1369_ (
		.din(new_net_924),
		.dout(_0673_)
	);

	and_bi _1370_ (
		.a(new_net_1432),
		.b(new_net_371),
		.c(_0674_)
	);

	or_bb _1371_ (
		.a(_0674_),
		.b(new_net_1104),
		.c(_0675_)
	);

	or_bi _1372_ (
		.a(new_net_1320),
		.b(new_net_814),
		.c(_0676_)
	);

	and_bi _1373_ (
		.a(_0676_),
		.b(new_net_1346),
		.c(_0677_)
	);

	or_bb _1374_ (
		.a(new_net_2134),
		.b(new_net_1262),
		.c(_0678_)
	);

	or_bb _1375_ (
		.a(new_net_2135),
		.b(new_net_1520),
		.c(_0679_)
	);

	and_bi _1376_ (
		.a(new_net_1513),
		.b(new_net_1465),
		.c(_0680_)
	);

	or_bi _1377_ (
		.a(_0680_),
		.b(new_net_1387),
		.c(_0681_)
	);

	and_bi _1378_ (
		.a(new_net_1254),
		.b(new_net_1685),
		.c(_0682_)
	);

	and_bi _1379_ (
		.a(new_net_1687),
		.b(new_net_1256),
		.c(_0683_)
	);

	or_bb _1380_ (
		.a(new_net_1429),
		.b(new_net_1410),
		.c(_0684_)
	);

	and_bi _1381_ (
		.a(new_net_1451),
		.b(new_net_1360),
		.c(_0685_)
	);

	and_bi _1382_ (
		.a(new_net_1361),
		.b(new_net_1450),
		.c(_0686_)
	);

	or_bb _1383_ (
		.a(_0686_),
		.b(_0685_),
		.c(_0687_)
	);

	or_bb _1384_ (
		.a(new_net_562),
		.b(new_net_1220),
		.c(_0688_)
	);

	inv _1385_ (
		.din(new_net_1255),
		.dout(_0689_)
	);

	or_bb _1386_ (
		.a(new_net_1466),
		.b(new_net_457),
		.c(_0690_)
	);

	and_bi _1387_ (
		.a(new_net_1472),
		.b(new_net_343),
		.c(_0691_)
	);

	and_bi _1388_ (
		.a(_0690_),
		.b(_0691_),
		.c(_0692_)
	);

	or_bb _1389_ (
		.a(_0692_),
		.b(new_net_1594),
		.c(_0693_)
	);

	or_ii _1390_ (
		.a(new_net_1467),
		.b(new_net_1689),
		.c(_0694_)
	);

	and_bi _1391_ (
		.a(new_net_1675),
		.b(new_net_1471),
		.c(_0695_)
	);

	and_bi _1392_ (
		.a(_0694_),
		.b(_0695_),
		.c(_0696_)
	);

	and_bi _1393_ (
		.a(new_net_1595),
		.b(_0696_),
		.c(_0697_)
	);

	and_bi _1394_ (
		.a(_0693_),
		.b(_0697_),
		.c(_0698_)
	);

	and_bi _1395_ (
		.a(new_net_1216),
		.b(new_net_171),
		.c(_0699_)
	);

	or_bb _1396_ (
		.a(_0699_),
		.b(new_net_612),
		.c(_0700_)
	);

	and_bi _1397_ (
		.a(_0688_),
		.b(new_net_2136),
		.c(_0701_)
	);

	and_ii _1398_ (
		.a(_0701_),
		.b(new_net_2137),
		.c(new_net_6)
	);

	and_bi _1399_ (
		.a(new_net_2138),
		.b(new_net_102),
		.c(_0702_)
	);

	and_bi _1400_ (
		.a(new_net_609),
		.b(new_net_1321),
		.c(_0703_)
	);

	or_bb _1401_ (
		.a(new_net_597),
		.b(new_net_975),
		.c(_0704_)
	);

	and_bb _1402_ (
		.a(new_net_600),
		.b(new_net_977),
		.c(_0705_)
	);

	and_bi _1403_ (
		.a(_0704_),
		.b(_0705_),
		.c(_0706_)
	);

	or_bb _1404_ (
		.a(new_net_234),
		.b(new_net_1236),
		.c(_0707_)
	);

	or_bi _1405_ (
		.a(new_net_1266),
		.b(new_net_1666),
		.c(_0708_)
	);

	and_bi _1406_ (
		.a(new_net_1270),
		.b(new_net_461),
		.c(_0709_)
	);

	and_bi _1407_ (
		.a(_0708_),
		.b(_0709_),
		.c(_0710_)
	);

	and_bi _1408_ (
		.a(new_net_1217),
		.b(new_net_1335),
		.c(_0711_)
	);

	or_bb _1409_ (
		.a(_0711_),
		.b(new_net_611),
		.c(_0712_)
	);

	and_bi _1410_ (
		.a(_0707_),
		.b(new_net_2139),
		.c(_0713_)
	);

	and_ii _1411_ (
		.a(_0713_),
		.b(new_net_2140),
		.c(new_net_8)
	);

	and_bi _1412_ (
		.a(new_net_2141),
		.b(new_net_103),
		.c(_0714_)
	);

	and_ii _1413_ (
		.a(new_net_399),
		.b(new_net_1433),
		.c(_0715_)
	);

	and_bi _1414_ (
		.a(new_net_178),
		.b(new_net_1183),
		.c(_0716_)
	);

	and_bi _1415_ (
		.a(new_net_1181),
		.b(new_net_179),
		.c(_0717_)
	);

	or_bb _1416_ (
		.a(_0717_),
		.b(_0716_),
		.c(_0718_)
	);

	or_bb _1417_ (
		.a(new_net_491),
		.b(new_net_1204),
		.c(_0719_)
	);

	or_bb _1418_ (
		.a(new_net_1608),
		.b(new_net_460),
		.c(_0720_)
	);

	and_bi _1419_ (
		.a(new_net_1603),
		.b(new_net_337),
		.c(_0721_)
	);

	and_bi _1420_ (
		.a(_0720_),
		.b(_0721_),
		.c(_0722_)
	);

	or_bb _1421_ (
		.a(_0722_),
		.b(new_net_1018),
		.c(_0723_)
	);

	or_ii _1422_ (
		.a(new_net_1693),
		.b(new_net_1609),
		.c(_0724_)
	);

	and_bi _1423_ (
		.a(new_net_1668),
		.b(new_net_1604),
		.c(_0725_)
	);

	and_bi _1424_ (
		.a(_0724_),
		.b(_0725_),
		.c(_0726_)
	);

	and_bi _1425_ (
		.a(new_net_1017),
		.b(_0726_),
		.c(_0727_)
	);

	and_bi _1426_ (
		.a(_0723_),
		.b(_0727_),
		.c(_0728_)
	);

	and_bi _1427_ (
		.a(new_net_1226),
		.b(new_net_653),
		.c(_0729_)
	);

	or_bb _1428_ (
		.a(_0729_),
		.b(new_net_627),
		.c(_0730_)
	);

	and_bi _1429_ (
		.a(_0719_),
		.b(new_net_2142),
		.c(_0731_)
	);

	and_ii _1430_ (
		.a(_0731_),
		.b(new_net_2143),
		.c(new_net_10)
	);

	and_bi _1431_ (
		.a(new_net_2144),
		.b(new_net_95),
		.c(_0732_)
	);

	or_ii _1432_ (
		.a(new_net_1548),
		.b(new_net_1142),
		.c(_0733_)
	);

	and_bi _1433_ (
		.a(new_net_2145),
		.b(new_net_1544),
		.c(_0734_)
	);

	and_bi _1434_ (
		.a(_0733_),
		.b(new_net_2146),
		.c(_0735_)
	);

	and_bi _1435_ (
		.a(new_net_1077),
		.b(new_net_784),
		.c(_0736_)
	);

	and_bi _1436_ (
		.a(new_net_787),
		.b(new_net_1078),
		.c(_0737_)
	);

	or_bb _1437_ (
		.a(new_net_1644),
		.b(new_net_1509),
		.c(_0738_)
	);

	inv _1438_ (
		.din(new_net_65),
		.dout(_0739_)
	);

	inv _1439_ (
		.din(new_net_995),
		.dout(_0740_)
	);

	or_ii _1440_ (
		.a(new_net_1552),
		.b(new_net_1174),
		.c(_0741_)
	);

	and_bi _1441_ (
		.a(new_net_2147),
		.b(new_net_1545),
		.c(_0742_)
	);

	or_bi _1442_ (
		.a(new_net_156),
		.b(new_net_362),
		.c(_0743_)
	);

	and_bi _1443_ (
		.a(new_net_257),
		.b(_0743_),
		.c(_0744_)
	);

	and_bi _1444_ (
		.a(new_net_363),
		.b(new_net_157),
		.c(_0745_)
	);

	and_bi _1445_ (
		.a(new_net_996),
		.b(new_net_202),
		.c(_0746_)
	);

	and_ii _1446_ (
		.a(new_net_212),
		.b(new_net_603),
		.c(_0747_)
	);

	or_bi _1447_ (
		.a(new_net_722),
		.b(new_net_863),
		.c(_0748_)
	);

	or_ii _1448_ (
		.a(new_net_1549),
		.b(new_net_1113),
		.c(_0749_)
	);

	and_bi _1449_ (
		.a(new_net_2148),
		.b(new_net_1546),
		.c(_0750_)
	);

	and_bi _1450_ (
		.a(_0749_),
		.b(new_net_2149),
		.c(_0751_)
	);

	and_bi _1451_ (
		.a(new_net_962),
		.b(new_net_313),
		.c(_0752_)
	);

	and_bi _1452_ (
		.a(new_net_314),
		.b(new_net_964),
		.c(_0753_)
	);

	or_bb _1453_ (
		.a(new_net_1511),
		.b(new_net_333),
		.c(_0754_)
	);

	or_ii _1454_ (
		.a(new_net_1561),
		.b(new_net_1071),
		.c(_0755_)
	);

	and_bi _1455_ (
		.a(new_net_2150),
		.b(new_net_1557),
		.c(_0756_)
	);

	and_bi _1456_ (
		.a(_0755_),
		.b(new_net_2151),
		.c(_0757_)
	);

	and_bi _1457_ (
		.a(new_net_262),
		.b(new_net_917),
		.c(_0758_)
	);

	and_bi _1458_ (
		.a(new_net_919),
		.b(new_net_265),
		.c(_0759_)
	);

	or_bb _1459_ (
		.a(new_net_477),
		.b(new_net_364),
		.c(_0760_)
	);

	or_bb _1460_ (
		.a(new_net_542),
		.b(new_net_1649),
		.c(_0761_)
	);

	or_bb _1461_ (
		.a(new_net_606),
		.b(new_net_970),
		.c(_0762_)
	);

	or_bi _1462_ (
		.a(new_net_698),
		.b(new_net_76),
		.c(_0763_)
	);

	and_bi _1463_ (
		.a(new_net_51),
		.b(new_net_529),
		.c(_0764_)
	);

	or_bi _1464_ (
		.a(new_net_699),
		.b(new_net_52),
		.c(_0765_)
	);

	and_bi _1465_ (
		.a(new_net_561),
		.b(new_net_604),
		.c(_0766_)
	);

	and_ii _1466_ (
		.a(new_net_334),
		.b(new_net_213),
		.c(_0767_)
	);

	and_bi _1467_ (
		.a(_0767_),
		.b(new_net_1099),
		.c(_0768_)
	);

	or_bb _1468_ (
		.a(_0768_),
		.b(new_net_1512),
		.c(_0769_)
	);

	and_ii _1469_ (
		.a(new_net_630),
		.b(new_net_365),
		.c(_0770_)
	);

	or_bb _1470_ (
		.a(_0770_),
		.b(new_net_479),
		.c(_0771_)
	);

	and_bi _1471_ (
		.a(new_net_1678),
		.b(new_net_78),
		.c(_0772_)
	);

	and_bi _1472_ (
		.a(new_net_77),
		.b(new_net_1679),
		.c(_0773_)
	);

	or_bb _1473_ (
		.a(_0773_),
		.b(_0772_),
		.c(_0774_)
	);

	and_bi _1474_ (
		.a(new_net_2152),
		.b(new_net_705),
		.c(_0775_)
	);

	or_bb _1475_ (
		.a(_0775_),
		.b(new_net_867),
		.c(_0776_)
	);

	or_bb _1476_ (
		.a(new_net_773),
		.b(new_net_1225),
		.c(_0777_)
	);

	inv _1477_ (
		.din(new_net_1079),
		.dout(_0778_)
	);

	or_bb _1478_ (
		.a(new_net_1144),
		.b(new_net_463),
		.c(_0779_)
	);

	and_bi _1479_ (
		.a(new_net_1137),
		.b(new_net_336),
		.c(_0780_)
	);

	and_bi _1480_ (
		.a(_0779_),
		.b(_0780_),
		.c(_0781_)
	);

	or_bb _1481_ (
		.a(_0781_),
		.b(new_net_810),
		.c(_0782_)
	);

	or_ii _1482_ (
		.a(new_net_1692),
		.b(new_net_1143),
		.c(_0783_)
	);

	and_bi _1483_ (
		.a(new_net_1669),
		.b(new_net_1138),
		.c(_0784_)
	);

	and_bi _1484_ (
		.a(new_net_2153),
		.b(_0784_),
		.c(_0785_)
	);

	and_bi _1485_ (
		.a(new_net_811),
		.b(_0785_),
		.c(_0786_)
	);

	and_bi _1486_ (
		.a(_0782_),
		.b(_0786_),
		.c(_0787_)
	);

	and_bi _1487_ (
		.a(new_net_1221),
		.b(new_net_949),
		.c(_0788_)
	);

	or_bb _1488_ (
		.a(_0788_),
		.b(new_net_616),
		.c(_0789_)
	);

	and_bi _1489_ (
		.a(_0777_),
		.b(new_net_2154),
		.c(_0790_)
	);

	and_ii _1490_ (
		.a(_0790_),
		.b(new_net_2155),
		.c(new_net_5)
	);

	and_bi _1491_ (
		.a(new_net_2156),
		.b(new_net_85),
		.c(_0791_)
	);

	or_bb _1492_ (
		.a(new_net_1651),
		.b(new_net_972),
		.c(_0792_)
	);

	and_bb _1493_ (
		.a(new_net_631),
		.b(_0792_),
		.c(_0793_)
	);

	or_bi _1494_ (
		.a(new_net_54),
		.b(new_net_634),
		.c(_0794_)
	);

	and_bi _1495_ (
		.a(new_net_2157),
		.b(new_net_1105),
		.c(_0795_)
	);

	or_ii _1496_ (
		.a(new_net_792),
		.b(new_net_543),
		.c(_0796_)
	);

	and_ii _1497_ (
		.a(new_net_793),
		.b(new_net_541),
		.c(_0797_)
	);

	and_bi _1498_ (
		.a(_0796_),
		.b(_0797_),
		.c(_0798_)
	);

	or_bb _1499_ (
		.a(new_net_1280),
		.b(new_net_1205),
		.c(_0799_)
	);

	inv _1500_ (
		.din(new_net_918),
		.dout(_0800_)
	);

	or_bb _1501_ (
		.a(new_net_1066),
		.b(new_net_458),
		.c(_0801_)
	);

	and_bi _1502_ (
		.a(new_net_1072),
		.b(new_net_344),
		.c(_0802_)
	);

	and_bi _1503_ (
		.a(_0801_),
		.b(_0802_),
		.c(_0803_)
	);

	or_bb _1504_ (
		.a(_0803_),
		.b(new_net_1299),
		.c(_0804_)
	);

	or_ii _1505_ (
		.a(new_net_1690),
		.b(new_net_1067),
		.c(_0805_)
	);

	and_bi _1506_ (
		.a(new_net_1676),
		.b(new_net_1073),
		.c(_0806_)
	);

	and_bi _1507_ (
		.a(_0805_),
		.b(_0806_),
		.c(_0807_)
	);

	and_bi _1508_ (
		.a(new_net_1300),
		.b(_0807_),
		.c(_0808_)
	);

	and_bi _1509_ (
		.a(_0804_),
		.b(_0808_),
		.c(_0809_)
	);

	and_bi _1510_ (
		.a(new_net_1237),
		.b(new_net_1427),
		.c(_0810_)
	);

	or_bb _1511_ (
		.a(_0810_),
		.b(new_net_618),
		.c(_0811_)
	);

	and_bi _1512_ (
		.a(_0799_),
		.b(new_net_2158),
		.c(_0812_)
	);

	and_ii _1513_ (
		.a(_0812_),
		.b(new_net_2159),
		.c(new_net_7)
	);

	and_bi _1514_ (
		.a(new_net_2160),
		.b(new_net_92),
		.c(_0813_)
	);

	and_ii _1515_ (
		.a(new_net_819),
		.b(new_net_560),
		.c(_0814_)
	);

	and_bi _1516_ (
		.a(new_net_864),
		.b(new_net_1540),
		.c(_0815_)
	);

	and_ii _1517_ (
		.a(new_net_1581),
		.b(new_net_211),
		.c(_0816_)
	);

	or_ii _1518_ (
		.a(new_net_1258),
		.b(new_net_1650),
		.c(_0817_)
	);

	or_bb _1519_ (
		.a(new_net_1259),
		.b(new_net_1648),
		.c(_0818_)
	);

	or_ii _1520_ (
		.a(_0818_),
		.b(_0817_),
		.c(_0819_)
	);

	or_bb _1521_ (
		.a(new_net_1703),
		.b(new_net_1206),
		.c(_0820_)
	);

	inv _1522_ (
		.din(new_net_963),
		.dout(_0821_)
	);

	or_bb _1523_ (
		.a(new_net_1108),
		.b(new_net_459),
		.c(_0822_)
	);

	and_bi _1524_ (
		.a(new_net_1115),
		.b(new_net_345),
		.c(_0823_)
	);

	and_bi _1525_ (
		.a(_0822_),
		.b(_0823_),
		.c(_0824_)
	);

	or_bb _1526_ (
		.a(_0824_),
		.b(new_net_46),
		.c(_0825_)
	);

	or_ii _1527_ (
		.a(new_net_1691),
		.b(new_net_1109),
		.c(_0826_)
	);

	and_bi _1528_ (
		.a(new_net_1677),
		.b(new_net_1114),
		.c(_0827_)
	);

	and_bi _1529_ (
		.a(new_net_2161),
		.b(_0827_),
		.c(_0828_)
	);

	and_bi _1530_ (
		.a(new_net_47),
		.b(_0828_),
		.c(_0829_)
	);

	and_bi _1531_ (
		.a(_0825_),
		.b(_0829_),
		.c(_0830_)
	);

	and_bi _1532_ (
		.a(new_net_1238),
		.b(new_net_1080),
		.c(_0831_)
	);

	or_bb _1533_ (
		.a(_0831_),
		.b(new_net_619),
		.c(_0832_)
	);

	and_bi _1534_ (
		.a(_0820_),
		.b(new_net_2162),
		.c(_0833_)
	);

	and_ii _1535_ (
		.a(_0833_),
		.b(new_net_2163),
		.c(new_net_9)
	);

	and_bi _1536_ (
		.a(new_net_2164),
		.b(new_net_90),
		.c(_0834_)
	);

	and_bi _1537_ (
		.a(new_net_1541),
		.b(new_net_865),
		.c(_0835_)
	);

	or_bb _1538_ (
		.a(new_net_2165),
		.b(new_net_1582),
		.c(_0836_)
	);

	or_bb _1539_ (
		.a(new_net_41),
		.b(new_net_1227),
		.c(_0837_)
	);

	or_bb _1540_ (
		.a(new_net_1176),
		.b(new_net_464),
		.c(_0838_)
	);

	and_bi _1541_ (
		.a(new_net_1169),
		.b(new_net_338),
		.c(_0839_)
	);

	and_bi _1542_ (
		.a(_0838_),
		.b(_0839_),
		.c(_0840_)
	);

	or_bb _1543_ (
		.a(_0840_),
		.b(new_net_258),
		.c(_0841_)
	);

	or_ii _1544_ (
		.a(new_net_1695),
		.b(new_net_1175),
		.c(_0842_)
	);

	and_bi _1545_ (
		.a(new_net_1670),
		.b(new_net_1170),
		.c(_0843_)
	);

	and_bi _1546_ (
		.a(_0842_),
		.b(_0843_),
		.c(_0844_)
	);

	and_bi _1547_ (
		.a(new_net_259),
		.b(_0844_),
		.c(_0845_)
	);

	and_bi _1548_ (
		.a(_0841_),
		.b(_0845_),
		.c(_0846_)
	);

	and_bi _1549_ (
		.a(new_net_1207),
		.b(new_net_925),
		.c(_0847_)
	);

	or_bb _1550_ (
		.a(_0847_),
		.b(new_net_628),
		.c(_0848_)
	);

	and_bi _1551_ (
		.a(_0837_),
		.b(new_net_2166),
		.c(_0849_)
	);

	and_ii _1552_ (
		.a(_0849_),
		.b(new_net_2167),
		.c(new_net_11)
	);

	and_bi _1553_ (
		.a(new_net_906),
		.b(new_net_98),
		.c(_0850_)
	);

	inv _1554_ (
		.din(new_net_1232),
		.dout(_0851_)
	);

	or_ii _1555_ (
		.a(new_net_1165),
		.b(new_net_585),
		.c(_0852_)
	);

	or_bb _1556_ (
		.a(new_net_1637),
		.b(new_net_1377),
		.c(_0853_)
	);

	and_bi _1557_ (
		.a(new_net_1635),
		.b(new_net_1038),
		.c(_0854_)
	);

	and_bi _1558_ (
		.a(_0853_),
		.b(_0854_),
		.c(_0855_)
	);

	and_bi _1559_ (
		.a(new_net_1208),
		.b(new_net_224),
		.c(_0856_)
	);

	or_bb _1560_ (
		.a(_0856_),
		.b(new_net_624),
		.c(_0857_)
	);

	and_bi _1561_ (
		.a(_0852_),
		.b(new_net_2168),
		.c(_0858_)
	);

	and_ii _1562_ (
		.a(_0858_),
		.b(new_net_2169),
		.c(new_net_18)
	);

	and_bi _1563_ (
		.a(new_net_2170),
		.b(new_net_99),
		.c(_0859_)
	);

	and_bb _1564_ (
		.a(new_net_1396),
		.b(new_net_1528),
		.c(_0860_)
	);

	and_bi _1565_ (
		.a(new_net_2171),
		.b(new_net_1514),
		.c(_0861_)
	);

	and_ii _1566_ (
		.a(_0861_),
		.b(_0860_),
		.c(_0862_)
	);

	and_bi _1567_ (
		.a(new_net_903),
		.b(new_net_33),
		.c(_0863_)
	);

	and_bi _1568_ (
		.a(new_net_35),
		.b(new_net_904),
		.c(_0864_)
	);

	and_bb _1569_ (
		.a(new_net_1412),
		.b(new_net_1517),
		.c(_0865_)
	);

	and_bi _1570_ (
		.a(new_net_2172),
		.b(new_net_1521),
		.c(_0866_)
	);

	and_ii _1571_ (
		.a(_0866_),
		.b(_0865_),
		.c(_0867_)
	);

	and_bi _1572_ (
		.a(new_net_1194),
		.b(new_net_682),
		.c(_0868_)
	);

	or_bi _1573_ (
		.a(new_net_58),
		.b(new_net_779),
		.c(_0869_)
	);

	and_bi _1574_ (
		.a(_0869_),
		.b(new_net_324),
		.c(_0870_)
	);

	and_ii _1575_ (
		.a(new_net_59),
		.b(new_net_325),
		.c(_0871_)
	);

	and_bi _1576_ (
		.a(new_net_685),
		.b(new_net_1196),
		.c(_0872_)
	);

	and_ii _1577_ (
		.a(new_net_1198),
		.b(new_net_781),
		.c(_0873_)
	);

	and_bb _1578_ (
		.a(new_net_228),
		.b(new_net_205),
		.c(_0874_)
	);

	and_bi _1579_ (
		.a(new_net_1362),
		.b(new_net_1430),
		.c(_0875_)
	);

	and_ii _1580_ (
		.a(_0875_),
		.b(new_net_1411),
		.c(_0876_)
	);

	and_bi _1581_ (
		.a(new_net_253),
		.b(new_net_1613),
		.c(_0877_)
	);

	and_bi _1582_ (
		.a(new_net_2173),
		.b(_0877_),
		.c(_0878_)
	);

	or_ii _1583_ (
		.a(new_net_144),
		.b(new_net_306),
		.c(_0879_)
	);

	and_ii _1584_ (
		.a(new_net_145),
		.b(new_net_310),
		.c(_0880_)
	);

	and_bi _1585_ (
		.a(_0879_),
		.b(_0880_),
		.c(_0881_)
	);

	or_bb _1586_ (
		.a(new_net_401),
		.b(new_net_1218),
		.c(_0882_)
	);

	or_bb _1587_ (
		.a(new_net_173),
		.b(new_net_987),
		.c(_0883_)
	);

	and_bi _1588_ (
		.a(new_net_177),
		.b(new_net_1012),
		.c(_0884_)
	);

	and_bi _1589_ (
		.a(_0883_),
		.b(_0884_),
		.c(_0885_)
	);

	and_bi _1590_ (
		.a(new_net_1239),
		.b(new_net_484),
		.c(_0886_)
	);

	or_bb _1591_ (
		.a(_0886_),
		.b(new_net_620),
		.c(_0887_)
	);

	and_bi _1592_ (
		.a(_0882_),
		.b(new_net_2174),
		.c(_0888_)
	);

	and_ii _1593_ (
		.a(_0888_),
		.b(new_net_2175),
		.c(new_net_19)
	);

	and_bi _1594_ (
		.a(new_net_2176),
		.b(new_net_91),
		.c(_0889_)
	);

	and_ii _1595_ (
		.a(new_net_1614),
		.b(new_net_1200),
		.c(_0890_)
	);

	and_bi _1596_ (
		.a(new_net_1617),
		.b(new_net_783),
		.c(_0891_)
	);

	or_bb _1597_ (
		.a(_0891_),
		.b(_0890_),
		.c(_0892_)
	);

	or_bi _1598_ (
		.a(new_net_1485),
		.b(new_net_207),
		.c(_0893_)
	);

	and_bi _1599_ (
		.a(new_net_1486),
		.b(new_net_206),
		.c(_0894_)
	);

	and_bi _1600_ (
		.a(_0893_),
		.b(_0894_),
		.c(_0895_)
	);

	or_bb _1601_ (
		.a(new_net_163),
		.b(new_net_1209),
		.c(_0896_)
	);

	inv _1602_ (
		.din(new_net_905),
		.dout(_0897_)
	);

	or_bb _1603_ (
		.a(new_net_1394),
		.b(new_net_979),
		.c(_0898_)
	);

	and_bi _1604_ (
		.a(new_net_1398),
		.b(new_net_1005),
		.c(_0899_)
	);

	and_bi _1605_ (
		.a(_0898_),
		.b(_0899_),
		.c(_0900_)
	);

	or_bb _1606_ (
		.a(_0900_),
		.b(new_net_346),
		.c(_0901_)
	);

	or_ii _1607_ (
		.a(new_net_1393),
		.b(new_net_1039),
		.c(_0902_)
	);

	and_bi _1608_ (
		.a(new_net_1379),
		.b(new_net_1397),
		.c(_0903_)
	);

	and_bi _1609_ (
		.a(_0902_),
		.b(_0903_),
		.c(_0904_)
	);

	and_bi _1610_ (
		.a(new_net_349),
		.b(_0904_),
		.c(_0905_)
	);

	and_bi _1611_ (
		.a(_0901_),
		.b(_0905_),
		.c(_0906_)
	);

	and_bi _1612_ (
		.a(new_net_1240),
		.b(new_net_842),
		.c(_0907_)
	);

	or_bb _1613_ (
		.a(_0907_),
		.b(new_net_621),
		.c(_0908_)
	);

	and_bi _1614_ (
		.a(_0896_),
		.b(new_net_2177),
		.c(_0909_)
	);

	or_bb _1615_ (
		.a(_0909_),
		.b(new_net_2178),
		.c(_0910_)
	);

	inv _1616_ (
		.din(new_net_890),
		.dout(new_net_2455)
	);

	and_bi _1617_ (
		.a(new_net_2179),
		.b(new_net_86),
		.c(_0911_)
	);

	and_bi _1618_ (
		.a(new_net_231),
		.b(new_net_1618),
		.c(_0912_)
	);

	or_bi _1619_ (
		.a(new_net_229),
		.b(new_net_1615),
		.c(_0913_)
	);

	and_bi _1620_ (
		.a(_0913_),
		.b(_0912_),
		.c(_0914_)
	);

	or_bb _1621_ (
		.a(new_net_350),
		.b(new_net_1228),
		.c(_0915_)
	);

	or_bb _1622_ (
		.a(new_net_1416),
		.b(new_net_983),
		.c(_0916_)
	);

	and_bi _1623_ (
		.a(new_net_1414),
		.b(new_net_1008),
		.c(_0917_)
	);

	and_bi _1624_ (
		.a(_0916_),
		.b(_0917_),
		.c(_0918_)
	);

	and_bi _1625_ (
		.a(new_net_1197),
		.b(_0918_),
		.c(_0919_)
	);

	or_ii _1626_ (
		.a(new_net_1417),
		.b(new_net_1045),
		.c(_0920_)
	);

	and_bi _1627_ (
		.a(new_net_1365),
		.b(new_net_1413),
		.c(_0921_)
	);

	and_bi _1628_ (
		.a(_0920_),
		.b(_0921_),
		.c(_0922_)
	);

	or_bb _1629_ (
		.a(_0922_),
		.b(new_net_1195),
		.c(_0923_)
	);

	and_bi _1630_ (
		.a(_0923_),
		.b(_0919_),
		.c(_0924_)
	);

	and_bi _1631_ (
		.a(new_net_1229),
		.b(new_net_1462),
		.c(_0925_)
	);

	or_bb _1632_ (
		.a(_0925_),
		.b(new_net_629),
		.c(_0926_)
	);

	and_bi _1633_ (
		.a(_0915_),
		.b(new_net_2180),
		.c(_0927_)
	);

	and_ii _1634_ (
		.a(_0927_),
		.b(new_net_2181),
		.c(new_net_22)
	);

	and_bi _1635_ (
		.a(new_net_2182),
		.b(new_net_96),
		.c(_0928_)
	);

	or_ii _1636_ (
		.a(new_net_838),
		.b(new_net_1562),
		.c(_0929_)
	);

	and_bi _1637_ (
		.a(new_net_2183),
		.b(new_net_1547),
		.c(_0930_)
	);

	and_bi _1638_ (
		.a(new_net_1343),
		.b(new_net_448),
		.c(_0931_)
	);

	and_bi _1639_ (
		.a(new_net_1094),
		.b(new_net_1383),
		.c(_0932_)
	);

	inv _1640_ (
		.din(new_net_1095),
		.dout(_0933_)
	);

	or_bi _1641_ (
		.a(new_net_449),
		.b(new_net_1344),
		.c(_0934_)
	);

	and_bi _1642_ (
		.a(new_net_1406),
		.b(new_net_777),
		.c(_0935_)
	);

	and_ii _1643_ (
		.a(new_net_849),
		.b(new_net_1389),
		.c(_0936_)
	);

	inv _1644_ (
		.din(new_net_770),
		.dout(_0937_)
	);

	or_ii _1645_ (
		.a(new_net_1556),
		.b(new_net_871),
		.c(_0938_)
	);

	and_bi _1646_ (
		.a(new_net_2184),
		.b(new_net_1554),
		.c(_0939_)
	);

	and_bi _1647_ (
		.a(_0938_),
		.b(new_net_2185),
		.c(_0940_)
	);

	or_bb _1648_ (
		.a(new_net_1564),
		.b(new_net_1060),
		.c(_0941_)
	);

	and_bi _1649_ (
		.a(new_net_1566),
		.b(new_net_771),
		.c(_0942_)
	);

	inv _1650_ (
		.din(new_net_825),
		.dout(_0943_)
	);

	or_ii _1651_ (
		.a(new_net_1558),
		.b(new_net_749),
		.c(_0944_)
	);

	and_bi _1652_ (
		.a(new_net_2186),
		.b(new_net_1550),
		.c(_0945_)
	);

	and_bi _1653_ (
		.a(_0944_),
		.b(new_net_2187),
		.c(_0946_)
	);

	or_bb _1654_ (
		.a(new_net_499),
		.b(new_net_1628),
		.c(_0947_)
	);

	and_bi _1655_ (
		.a(new_net_500),
		.b(new_net_828),
		.c(_0948_)
	);

	inv _1656_ (
		.din(new_net_1053),
		.dout(_0949_)
	);

	or_ii _1657_ (
		.a(new_net_1559),
		.b(new_net_951),
		.c(_0950_)
	);

	and_bi _1658_ (
		.a(new_net_2188),
		.b(new_net_1551),
		.c(_0951_)
	);

	and_bi _1659_ (
		.a(new_net_127),
		.b(new_net_901),
		.c(_0952_)
	);

	or_bb _1660_ (
		.a(new_net_158),
		.b(new_net_741),
		.c(_0953_)
	);

	and_ii _1661_ (
		.a(new_net_1131),
		.b(new_net_655),
		.c(_0954_)
	);

	and_bi _1662_ (
		.a(new_net_43),
		.b(new_net_1294),
		.c(_0955_)
	);

	and_ii _1663_ (
		.a(new_net_198),
		.b(new_net_1599),
		.c(_0956_)
	);

	and_bi _1664_ (
		.a(new_net_1585),
		.b(new_net_1435),
		.c(_0957_)
	);

	or_bb _1665_ (
		.a(new_net_540),
		.b(new_net_67),
		.c(_0958_)
	);

	and_ii _1666_ (
		.a(new_net_633),
		.b(new_net_2189),
		.c(_0959_)
	);

	and_bi _1667_ (
		.a(new_net_478),
		.b(new_net_1645),
		.c(_0960_)
	);

	or_bb _1668_ (
		.a(_0960_),
		.b(new_net_1510),
		.c(_0961_)
	);

	or_bb _1669_ (
		.a(new_net_2190),
		.b(_0959_),
		.c(_0962_)
	);

	and_ii _1670_ (
		.a(new_net_409),
		.b(new_net_868),
		.c(_0963_)
	);

	and_bi _1671_ (
		.a(new_net_1588),
		.b(new_net_1601),
		.c(_0964_)
	);

	and_bi _1672_ (
		.a(new_net_45),
		.b(new_net_657),
		.c(_0965_)
	);

	or_bi _1673_ (
		.a(new_net_902),
		.b(new_net_128),
		.c(_0966_)
	);

	or_bb _1674_ (
		.a(_0966_),
		.b(new_net_1055),
		.c(_0967_)
	);

	or_ii _1675_ (
		.a(new_net_452),
		.b(new_net_1133),
		.c(_0968_)
	);

	and_bi _1676_ (
		.a(new_net_405),
		.b(new_net_472),
		.c(_0969_)
	);

	or_ii _1677_ (
		.a(new_net_1035),
		.b(new_net_389),
		.c(_0970_)
	);

	and_ii _1678_ (
		.a(new_net_1157),
		.b(new_net_358),
		.c(_0971_)
	);

	and_bi _1679_ (
		.a(new_net_1579),
		.b(_0971_),
		.c(_0972_)
	);

	and_bi _1680_ (
		.a(new_net_521),
		.b(new_net_1446),
		.c(_0973_)
	);

	and_bi _1681_ (
		.a(new_net_1444),
		.b(new_net_522),
		.c(_0974_)
	);

	and_ii _1682_ (
		.a(_0974_),
		.b(_0973_),
		.c(_0975_)
	);

	or_ii _1683_ (
		.a(new_net_1719),
		.b(new_net_587),
		.c(_0976_)
	);

	or_bb _1684_ (
		.a(new_net_839),
		.b(new_net_1013),
		.c(_0977_)
	);

	and_bi _1685_ (
		.a(new_net_835),
		.b(new_net_978),
		.c(_0978_)
	);

	and_bi _1686_ (
		.a(_0977_),
		.b(_0978_),
		.c(_0979_)
	);

	and_bi _1687_ (
		.a(new_net_1096),
		.b(_0979_),
		.c(_0980_)
	);

	or_ii _1688_ (
		.a(new_net_840),
		.b(new_net_1378),
		.c(_0981_)
	);

	and_bi _1689_ (
		.a(new_net_1040),
		.b(new_net_836),
		.c(_0982_)
	);

	and_bi _1690_ (
		.a(_0981_),
		.b(_0982_),
		.c(_0983_)
	);

	and_bi _1691_ (
		.a(new_net_1407),
		.b(_0983_),
		.c(_0984_)
	);

	and_ii _1692_ (
		.a(_0984_),
		.b(_0980_),
		.c(_0985_)
	);

	and_bi _1693_ (
		.a(new_net_1234),
		.b(new_net_735),
		.c(_0986_)
	);

	or_bb _1694_ (
		.a(_0986_),
		.b(new_net_615),
		.c(_0987_)
	);

	and_bi _1695_ (
		.a(_0976_),
		.b(new_net_2191),
		.c(_0988_)
	);

	and_ii _1696_ (
		.a(_0988_),
		.b(new_net_2192),
		.c(new_net_17)
	);

	and_bi _1697_ (
		.a(new_net_2193),
		.b(new_net_88),
		.c(_0989_)
	);

	and_bi _1698_ (
		.a(new_net_1036),
		.b(new_net_361),
		.c(_0990_)
	);

	and_bi _1699_ (
		.a(new_net_199),
		.b(_0990_),
		.c(_0991_)
	);

	or_bb _1700_ (
		.a(new_net_72),
		.b(new_net_392),
		.c(_0992_)
	);

	and_bb _1701_ (
		.a(new_net_73),
		.b(new_net_390),
		.c(_0993_)
	);

	and_bi _1702_ (
		.a(_0992_),
		.b(_0993_),
		.c(_0994_)
	);

	or_bb _1703_ (
		.a(new_net_1161),
		.b(new_net_1222),
		.c(_0995_)
	);

	or_bb _1704_ (
		.a(new_net_877),
		.b(new_net_465),
		.c(_0996_)
	);

	and_bi _1705_ (
		.a(new_net_872),
		.b(new_net_339),
		.c(_0997_)
	);

	and_bi _1706_ (
		.a(_0996_),
		.b(_0997_),
		.c(_0998_)
	);

	or_bb _1707_ (
		.a(_0998_),
		.b(new_net_1063),
		.c(_0999_)
	);

	or_ii _1708_ (
		.a(new_net_1696),
		.b(new_net_878),
		.c(_1000_)
	);

	and_bi _1709_ (
		.a(new_net_1671),
		.b(new_net_873),
		.c(_1001_)
	);

	and_bi _1710_ (
		.a(_1000_),
		.b(_1001_),
		.c(_1002_)
	);

	and_bi _1711_ (
		.a(new_net_1062),
		.b(_1002_),
		.c(_1003_)
	);

	and_bi _1712_ (
		.a(_0999_),
		.b(_1003_),
		.c(_1004_)
	);

	and_bi _1713_ (
		.a(new_net_1223),
		.b(new_net_503),
		.c(_1005_)
	);

	or_bb _1714_ (
		.a(_1005_),
		.b(new_net_617),
		.c(_1006_)
	);

	and_bi _1715_ (
		.a(_0995_),
		.b(new_net_2194),
		.c(_1007_)
	);

	and_ii _1716_ (
		.a(_1007_),
		.b(new_net_2195),
		.c(new_net_20)
	);

	and_bi _1717_ (
		.a(new_net_2196),
		.b(new_net_89),
		.c(_1008_)
	);

	and_bi _1718_ (
		.a(new_net_455),
		.b(new_net_359),
		.c(_1009_)
	);

	and_bb _1719_ (
		.a(new_net_356),
		.b(new_net_1134),
		.c(_1010_)
	);

	and_ii _1720_ (
		.a(_1010_),
		.b(_1009_),
		.c(_1011_)
	);

	or_bb _1721_ (
		.a(new_net_1186),
		.b(new_net_406),
		.c(_1012_)
	);

	or_bi _1722_ (
		.a(new_net_656),
		.b(new_net_44),
		.c(_1013_)
	);

	and_bi _1723_ (
		.a(new_net_1187),
		.b(new_net_507),
		.c(_1014_)
	);

	and_bi _1724_ (
		.a(_1012_),
		.b(_1014_),
		.c(_1015_)
	);

	or_bb _1725_ (
		.a(new_net_1597),
		.b(new_net_1210),
		.c(_1016_)
	);

	or_bb _1726_ (
		.a(new_net_756),
		.b(new_net_466),
		.c(_1017_)
	);

	and_bi _1727_ (
		.a(new_net_751),
		.b(new_net_340),
		.c(_1018_)
	);

	and_bi _1728_ (
		.a(_1017_),
		.b(_1018_),
		.c(_1019_)
	);

	and_bi _1729_ (
		.a(new_net_827),
		.b(_1019_),
		.c(_1020_)
	);

	or_ii _1730_ (
		.a(new_net_1697),
		.b(new_net_755),
		.c(_1021_)
	);

	and_bi _1731_ (
		.a(new_net_1672),
		.b(new_net_750),
		.c(_1022_)
	);

	and_bi _1732_ (
		.a(_1021_),
		.b(_1022_),
		.c(_1023_)
	);

	and_bi _1733_ (
		.a(new_net_1629),
		.b(_1023_),
		.c(_1024_)
	);

	and_ii _1734_ (
		.a(_1024_),
		.b(_1020_),
		.c(_1025_)
	);

	and_bi _1735_ (
		.a(new_net_1211),
		.b(new_net_694),
		.c(_1026_)
	);

	or_bb _1736_ (
		.a(_1026_),
		.b(new_net_625),
		.c(_1027_)
	);

	and_bi _1737_ (
		.a(_1016_),
		.b(new_net_2197),
		.c(_1028_)
	);

	and_ii _1738_ (
		.a(_1028_),
		.b(new_net_2198),
		.c(new_net_21)
	);

	and_bi _1739_ (
		.a(new_net_2199),
		.b(new_net_97),
		.c(_1029_)
	);

	or_ii _1740_ (
		.a(new_net_473),
		.b(new_net_360),
		.c(_1030_)
	);

	and_ii _1741_ (
		.a(new_net_474),
		.b(new_net_357),
		.c(_1031_)
	);

	and_bi _1742_ (
		.a(_1030_),
		.b(_1031_),
		.c(_1032_)
	);

	or_bb _1743_ (
		.a(new_net_82),
		.b(new_net_1224),
		.c(_1033_)
	);

	or_bb _1744_ (
		.a(new_net_958),
		.b(new_net_467),
		.c(_1034_)
	);

	and_bi _1745_ (
		.a(new_net_952),
		.b(new_net_341),
		.c(_1035_)
	);

	and_bi _1746_ (
		.a(_1034_),
		.b(_1035_),
		.c(_1036_)
	);

	or_bb _1747_ (
		.a(_1036_),
		.b(new_net_743),
		.c(_1037_)
	);

	or_ii _1748_ (
		.a(new_net_1698),
		.b(new_net_957),
		.c(_1038_)
	);

	and_bi _1749_ (
		.a(new_net_1673),
		.b(new_net_953),
		.c(_1039_)
	);

	and_bi _1750_ (
		.a(_1038_),
		.b(_1039_),
		.c(_1040_)
	);

	and_bi _1751_ (
		.a(new_net_744),
		.b(_1040_),
		.c(_1041_)
	);

	and_bi _1752_ (
		.a(_1037_),
		.b(_1041_),
		.c(_1042_)
	);

	and_bi _1753_ (
		.a(new_net_1235),
		.b(new_net_1056),
		.c(_1043_)
	);

	or_bb _1754_ (
		.a(_1043_),
		.b(new_net_613),
		.c(_1044_)
	);

	and_bi _1755_ (
		.a(_1033_),
		.b(new_net_2200),
		.c(_1045_)
	);

	and_ii _1756_ (
		.a(_1045_),
		.b(new_net_2201),
		.c(new_net_23)
	);

	inv _1757_ (
		.din(new_net_122),
		.dout(_1046_)
	);

	inv _1758_ (
		.din(new_net_662),
		.dout(_1047_)
	);

	and_bi _1759_ (
		.a(new_net_210),
		.b(new_net_721),
		.c(_1048_)
	);

	and_bi _1760_ (
		.a(new_net_723),
		.b(new_net_866),
		.c(_1049_)
	);

	and_bi _1761_ (
		.a(new_net_971),
		.b(new_net_2202),
		.c(_1050_)
	);

	or_bb _1762_ (
		.a(new_net_214),
		.b(new_net_559),
		.c(_1051_)
	);

	or_bi _1763_ (
		.a(new_net_1100),
		.b(_1051_),
		.c(_1052_)
	);

	and_bi _1764_ (
		.a(new_net_2203),
		.b(new_net_195),
		.c(_1053_)
	);

	or_bb _1765_ (
		.a(_1053_),
		.b(new_net_2204),
		.c(_1054_)
	);

	and_bi _1766_ (
		.a(new_net_1329),
		.b(new_net_635),
		.c(_1055_)
	);

	and_bi _1767_ (
		.a(new_net_632),
		.b(new_net_1330),
		.c(_1056_)
	);

	or_bb _1768_ (
		.a(_1056_),
		.b(_1055_),
		.c(_1057_)
	);

	or_bb _1769_ (
		.a(new_net_1381),
		.b(new_net_706),
		.c(_1058_)
	);

	and_bb _1770_ (
		.a(new_net_1382),
		.b(new_net_707),
		.c(_1059_)
	);

	or_bb _1771_ (
		.a(_1059_),
		.b(new_net_1419),
		.c(_1060_)
	);

	and_bi _1772_ (
		.a(new_net_2205),
		.b(_1060_),
		.c(_1061_)
	);

	and_ii _1773_ (
		.a(new_net_605),
		.b(new_net_642),
		.c(_1062_)
	);

	and_bi _1774_ (
		.a(new_net_641),
		.b(new_net_215),
		.c(_1063_)
	);

	and_ii _1775_ (
		.a(_1063_),
		.b(new_net_2206),
		.c(_1064_)
	);

	or_bb _1776_ (
		.a(new_net_1577),
		.b(new_net_1107),
		.c(_1065_)
	);

	and_bb _1777_ (
		.a(new_net_1578),
		.b(new_net_1106),
		.c(_1066_)
	);

	and_bi _1778_ (
		.a(_1065_),
		.b(_1066_),
		.c(_1067_)
	);

	or_bb _1779_ (
		.a(new_net_196),
		.b(new_net_79),
		.c(_1068_)
	);

	and_bi _1780_ (
		.a(new_net_197),
		.b(new_net_66),
		.c(_1069_)
	);

	or_bi _1781_ (
		.a(_1069_),
		.b(_1068_),
		.c(_1070_)
	);

	and_bi _1782_ (
		.a(new_net_700),
		.b(new_net_1680),
		.c(_1071_)
	);

	or_bi _1783_ (
		.a(new_net_487),
		.b(new_net_1701),
		.c(_1072_)
	);

	and_bi _1784_ (
		.a(new_net_488),
		.b(new_net_1702),
		.c(_1073_)
	);

	or_bi _1785_ (
		.a(_1073_),
		.b(_1072_),
		.c(_1074_)
	);

	or_bi _1786_ (
		.a(new_net_1589),
		.b(new_net_997),
		.c(_1075_)
	);

	inv _1787_ (
		.din(new_net_1420),
		.dout(_1076_)
	);

	and_bi _1788_ (
		.a(new_net_1590),
		.b(new_net_998),
		.c(_1077_)
	);

	or_bb _1789_ (
		.a(_1077_),
		.b(new_net_1282),
		.c(_1078_)
	);

	and_bi _1790_ (
		.a(new_net_2207),
		.b(_1078_),
		.c(_1079_)
	);

	or_bb _1791_ (
		.a(_1079_),
		.b(_1061_),
		.c(_1080_)
	);

	or_bi _1792_ (
		.a(new_net_1037),
		.b(new_net_201),
		.c(_1081_)
	);

	and_bb _1793_ (
		.a(new_net_68),
		.b(new_net_1587),
		.c(_1082_)
	);

	or_bb _1794_ (
		.a(_1082_),
		.b(new_net_1600),
		.c(_1083_)
	);

	or_bb _1795_ (
		.a(new_net_407),
		.b(new_net_1445),
		.c(_1084_)
	);

	and_bi _1796_ (
		.a(new_net_1447),
		.b(new_net_508),
		.c(_1085_)
	);

	or_bi _1797_ (
		.a(new_net_475),
		.b(new_net_368),
		.c(_1086_)
	);

	and_bi _1798_ (
		.a(new_net_1132),
		.b(new_net_69),
		.c(_1087_)
	);

	or_bb _1799_ (
		.a(_1087_),
		.b(new_net_1295),
		.c(_1088_)
	);

	or_bb _1800_ (
		.a(new_net_701),
		.b(new_net_547),
		.c(_1089_)
	);

	and_bi _1801_ (
		.a(new_net_369),
		.b(new_net_476),
		.c(_1090_)
	);

	and_bi _1802_ (
		.a(new_net_702),
		.b(new_net_884),
		.c(_1091_)
	);

	and_bi _1803_ (
		.a(_1089_),
		.b(_1091_),
		.c(_1092_)
	);

	and_bi _1804_ (
		.a(new_net_446),
		.b(new_net_266),
		.c(_1093_)
	);

	and_bi _1805_ (
		.a(new_net_267),
		.b(new_net_447),
		.c(_1094_)
	);

	or_bb _1806_ (
		.a(_1094_),
		.b(_1093_),
		.c(_1095_)
	);

	or_bi _1807_ (
		.a(new_net_1423),
		.b(new_net_408),
		.c(_1096_)
	);

	and_bb _1808_ (
		.a(new_net_200),
		.b(new_net_1586),
		.c(_1097_)
	);

	and_ii _1809_ (
		.a(new_net_2208),
		.b(new_net_1436),
		.c(_1098_)
	);

	or_bi _1810_ (
		.a(new_net_393),
		.b(new_net_454),
		.c(_1099_)
	);

	and_bi _1811_ (
		.a(new_net_391),
		.b(new_net_453),
		.c(_1100_)
	);

	or_bi _1812_ (
		.a(_1100_),
		.b(_1099_),
		.c(_1101_)
	);

	or_bb _1813_ (
		.a(new_net_372),
		.b(new_net_548),
		.c(_1102_)
	);

	and_bi _1814_ (
		.a(new_net_373),
		.b(new_net_885),
		.c(_1103_)
	);

	and_bi _1815_ (
		.a(_1102_),
		.b(_1103_),
		.c(_1104_)
	);

	or_bi _1816_ (
		.a(new_net_70),
		.b(new_net_638),
		.c(_1105_)
	);

	and_bi _1817_ (
		.a(new_net_71),
		.b(new_net_639),
		.c(_1106_)
	);

	or_bb _1818_ (
		.a(_1106_),
		.b(new_net_410),
		.c(_1107_)
	);

	or_bi _1819_ (
		.a(_1107_),
		.b(new_net_2209),
		.c(_1108_)
	);

	or_ii _1820_ (
		.a(new_net_690),
		.b(new_net_1283),
		.c(_1109_)
	);

	and_bi _1821_ (
		.a(_1096_),
		.b(new_net_2210),
		.c(_1110_)
	);

	and_bi _1822_ (
		.a(new_net_532),
		.b(new_net_412),
		.c(_1111_)
	);

	or_bb _1823_ (
		.a(new_net_2211),
		.b(new_net_1424),
		.c(_1112_)
	);

	and_bi _1824_ (
		.a(new_net_530),
		.b(new_net_691),
		.c(_1113_)
	);

	or_bb _1825_ (
		.a(_1113_),
		.b(new_net_1284),
		.c(_1114_)
	);

	and_bi _1826_ (
		.a(_1112_),
		.b(_1114_),
		.c(_1115_)
	);

	or_bb _1827_ (
		.a(_1115_),
		.b(_1110_),
		.c(_1116_)
	);

	and_bb _1828_ (
		.a(new_net_544),
		.b(new_net_1652),
		.c(_1117_)
	);

	and_bi _1829_ (
		.a(new_net_607),
		.b(new_net_2212),
		.c(_1118_)
	);

	or_bb _1830_ (
		.a(new_net_527),
		.b(new_net_833),
		.c(_1119_)
	);

	and_bb _1831_ (
		.a(new_net_528),
		.b(new_net_834),
		.c(_1120_)
	);

	and_bi _1832_ (
		.a(_1119_),
		.b(_1120_),
		.c(_1121_)
	);

	and_ii _1833_ (
		.a(new_net_806),
		.b(new_net_1683),
		.c(_1122_)
	);

	and_bb _1834_ (
		.a(new_net_807),
		.b(new_net_1684),
		.c(_1123_)
	);

	or_bb _1835_ (
		.a(_1123_),
		.b(new_net_1212),
		.c(_1124_)
	);

	or_bb _1836_ (
		.a(_1124_),
		.b(new_net_2213),
		.c(_1125_)
	);

	or_bb _1837_ (
		.a(new_net_874),
		.b(new_net_988),
		.c(_1126_)
	);

	and_bi _1838_ (
		.a(new_net_879),
		.b(new_net_1014),
		.c(_1127_)
	);

	and_bi _1839_ (
		.a(_1126_),
		.b(_1127_),
		.c(_1128_)
	);

	and_bi _1840_ (
		.a(new_net_772),
		.b(_1128_),
		.c(_1129_)
	);

	or_ii _1841_ (
		.a(new_net_875),
		.b(new_net_1041),
		.c(_1130_)
	);

	and_bi _1842_ (
		.a(new_net_1369),
		.b(new_net_880),
		.c(_1131_)
	);

	and_bi _1843_ (
		.a(_1130_),
		.b(_1131_),
		.c(_1132_)
	);

	and_bi _1844_ (
		.a(new_net_1061),
		.b(_1132_),
		.c(_1133_)
	);

	and_ii _1845_ (
		.a(_1133_),
		.b(_1129_),
		.c(_1134_)
	);

	or_bb _1846_ (
		.a(new_net_757),
		.b(new_net_991),
		.c(_1135_)
	);

	and_bi _1847_ (
		.a(new_net_752),
		.b(new_net_1001),
		.c(_1136_)
	);

	and_bi _1848_ (
		.a(_1135_),
		.b(_1136_),
		.c(_1137_)
	);

	and_bi _1849_ (
		.a(new_net_826),
		.b(_1137_),
		.c(_1138_)
	);

	or_ii _1850_ (
		.a(new_net_758),
		.b(new_net_1046),
		.c(_1139_)
	);

	and_bi _1851_ (
		.a(new_net_1373),
		.b(new_net_753),
		.c(_1140_)
	);

	and_bi _1852_ (
		.a(_1139_),
		.b(_1140_),
		.c(_1141_)
	);

	and_bi _1853_ (
		.a(new_net_1630),
		.b(_1141_),
		.c(_1142_)
	);

	and_ii _1854_ (
		.a(_1142_),
		.b(_1138_),
		.c(_1143_)
	);

	and_bi _1855_ (
		.a(new_net_1408),
		.b(new_net_470),
		.c(_1144_)
	);

	and_bi _1856_ (
		.a(new_net_471),
		.b(new_net_1409),
		.c(_1145_)
	);

	and_ii _1857_ (
		.a(_1145_),
		.b(_1144_),
		.c(_1146_)
	);

	or_bb _1858_ (
		.a(new_net_959),
		.b(new_net_992),
		.c(_1147_)
	);

	and_bi _1859_ (
		.a(new_net_954),
		.b(new_net_1002),
		.c(_1148_)
	);

	and_bi _1860_ (
		.a(_1147_),
		.b(_1148_),
		.c(_1149_)
	);

	and_bi _1861_ (
		.a(new_net_1054),
		.b(_1149_),
		.c(_1150_)
	);

	or_ii _1862_ (
		.a(new_net_960),
		.b(new_net_1047),
		.c(_1151_)
	);

	and_bi _1863_ (
		.a(new_net_1374),
		.b(new_net_955),
		.c(_1152_)
	);

	and_bi _1864_ (
		.a(_1151_),
		.b(_1152_),
		.c(_1153_)
	);

	and_bi _1865_ (
		.a(new_net_742),
		.b(_1153_),
		.c(_1154_)
	);

	and_ii _1866_ (
		.a(_1154_),
		.b(_1150_),
		.c(_1155_)
	);

	and_ii _1867_ (
		.a(new_net_1709),
		.b(new_net_738),
		.c(_1156_)
	);

	and_bb _1868_ (
		.a(new_net_1710),
		.b(new_net_736),
		.c(_1157_)
	);

	and_ii _1869_ (
		.a(_1157_),
		.b(_1156_),
		.c(_1158_)
	);

	and_bb _1870_ (
		.a(new_net_831),
		.b(new_net_1456),
		.c(_1159_)
	);

	and_ii _1871_ (
		.a(new_net_832),
		.b(new_net_1457),
		.c(_1160_)
	);

	or_bb _1872_ (
		.a(_1160_),
		.b(_1159_),
		.c(_1161_)
	);

	or_bb _1873_ (
		.a(new_net_1171),
		.b(new_net_989),
		.c(_1162_)
	);

	and_bi _1874_ (
		.a(new_net_1177),
		.b(new_net_1015),
		.c(_1163_)
	);

	and_bi _1875_ (
		.a(_1162_),
		.b(_1163_),
		.c(_1164_)
	);

	or_bb _1876_ (
		.a(_1164_),
		.b(new_net_261),
		.c(_1165_)
	);

	or_ii _1877_ (
		.a(new_net_1172),
		.b(new_net_1042),
		.c(_1166_)
	);

	and_bi _1878_ (
		.a(new_net_1370),
		.b(new_net_1178),
		.c(_1167_)
	);

	and_bi _1879_ (
		.a(_1166_),
		.b(_1167_),
		.c(_1168_)
	);

	and_bi _1880_ (
		.a(new_net_260),
		.b(_1168_),
		.c(_1169_)
	);

	and_bi _1881_ (
		.a(_1165_),
		.b(_1169_),
		.c(_1170_)
	);

	or_bb _1882_ (
		.a(new_net_1116),
		.b(new_net_993),
		.c(_1171_)
	);

	and_bi _1883_ (
		.a(new_net_1110),
		.b(new_net_1003),
		.c(_1172_)
	);

	and_bi _1884_ (
		.a(_1171_),
		.b(_1172_),
		.c(_1173_)
	);

	or_bb _1885_ (
		.a(_1173_),
		.b(new_net_48),
		.c(_1174_)
	);

	or_ii _1886_ (
		.a(new_net_1117),
		.b(new_net_1048),
		.c(_1175_)
	);

	and_bi _1887_ (
		.a(new_net_1375),
		.b(new_net_1111),
		.c(_1176_)
	);

	and_bi _1888_ (
		.a(_1175_),
		.b(_1176_),
		.c(_1177_)
	);

	and_bi _1889_ (
		.a(new_net_49),
		.b(_1177_),
		.c(_1178_)
	);

	and_bi _1890_ (
		.a(_1174_),
		.b(_1178_),
		.c(_1179_)
	);

	and_ii _1891_ (
		.a(new_net_1318),
		.b(new_net_1646),
		.c(_1180_)
	);

	and_bb _1892_ (
		.a(new_net_1319),
		.b(new_net_1647),
		.c(_1181_)
	);

	and_ii _1893_ (
		.a(_1181_),
		.b(_1180_),
		.c(_1182_)
	);

	or_bb _1894_ (
		.a(new_net_1145),
		.b(new_net_994),
		.c(_1183_)
	);

	and_bi _1895_ (
		.a(new_net_1139),
		.b(new_net_1004),
		.c(_1184_)
	);

	and_bi _1896_ (
		.a(_1183_),
		.b(_1184_),
		.c(_1185_)
	);

	or_bb _1897_ (
		.a(_1185_),
		.b(new_net_812),
		.c(_1186_)
	);

	or_ii _1898_ (
		.a(new_net_1146),
		.b(new_net_1049),
		.c(_1187_)
	);

	and_bi _1899_ (
		.a(new_net_1376),
		.b(new_net_1140),
		.c(_1188_)
	);

	and_bi _1900_ (
		.a(_1187_),
		.b(_1188_),
		.c(_1189_)
	);

	and_bi _1901_ (
		.a(new_net_813),
		.b(_1189_),
		.c(_1190_)
	);

	and_bi _1902_ (
		.a(_1186_),
		.b(_1190_),
		.c(_1191_)
	);

	or_bb _1903_ (
		.a(new_net_1246),
		.b(new_net_980),
		.c(_1192_)
	);

	and_bi _1904_ (
		.a(new_net_1251),
		.b(new_net_1006),
		.c(_1193_)
	);

	and_bi _1905_ (
		.a(_1192_),
		.b(_1193_),
		.c(_1194_)
	);

	or_bb _1906_ (
		.a(_1194_),
		.b(new_net_1292),
		.c(_1195_)
	);

	or_ii _1907_ (
		.a(new_net_1247),
		.b(new_net_1043),
		.c(_1196_)
	);

	and_bi _1908_ (
		.a(new_net_1380),
		.b(new_net_1252),
		.c(_1197_)
	);

	and_bi _1909_ (
		.a(_1196_),
		.b(_1197_),
		.c(_1198_)
	);

	and_bi _1910_ (
		.a(new_net_1291),
		.b(_1198_),
		.c(_1199_)
	);

	and_bi _1911_ (
		.a(_1195_),
		.b(_1199_),
		.c(_1200_)
	);

	or_bb _1912_ (
		.a(new_net_1074),
		.b(new_net_984),
		.c(_1201_)
	);

	and_bi _1913_ (
		.a(new_net_1068),
		.b(new_net_1009),
		.c(_1202_)
	);

	and_bi _1914_ (
		.a(_1201_),
		.b(_1202_),
		.c(_1203_)
	);

	and_bi _1915_ (
		.a(new_net_920),
		.b(_1203_),
		.c(_1204_)
	);

	or_ii _1916_ (
		.a(new_net_1075),
		.b(new_net_1050),
		.c(_1205_)
	);

	and_bi _1917_ (
		.a(new_net_1366),
		.b(new_net_1069),
		.c(_1206_)
	);

	and_bi _1918_ (
		.a(_1205_),
		.b(_1206_),
		.c(_1207_)
	);

	and_bi _1919_ (
		.a(new_net_1301),
		.b(_1207_),
		.c(_1208_)
	);

	and_ii _1920_ (
		.a(_1208_),
		.b(_1204_),
		.c(_1209_)
	);

	or_bb _1921_ (
		.a(new_net_595),
		.b(new_net_1402),
		.c(_1210_)
	);

	and_bb _1922_ (
		.a(new_net_596),
		.b(new_net_1403),
		.c(_1211_)
	);

	and_bi _1923_ (
		.a(_1210_),
		.b(_1211_),
		.c(_1212_)
	);

	and_ii _1924_ (
		.a(new_net_289),
		.b(new_net_366),
		.c(_1213_)
	);

	and_bb _1925_ (
		.a(new_net_290),
		.b(new_net_367),
		.c(_1214_)
	);

	and_ii _1926_ (
		.a(_1214_),
		.b(_1213_),
		.c(_1215_)
	);

	and_ii _1927_ (
		.a(new_net_1241),
		.b(new_net_1097),
		.c(_1216_)
	);

	and_bb _1928_ (
		.a(new_net_1242),
		.b(new_net_1098),
		.c(_1217_)
	);

	or_bb _1929_ (
		.a(_1217_),
		.b(_1216_),
		.c(_1218_)
	);

	or_bi _1930_ (
		.a(new_net_869),
		.b(new_net_1491),
		.c(_1219_)
	);

	and_bi _1931_ (
		.a(new_net_870),
		.b(new_net_1492),
		.c(_1220_)
	);

	or_bb _1932_ (
		.a(_1220_),
		.b(new_net_586),
		.c(_1221_)
	);

	and_bi _1933_ (
		.a(new_net_2214),
		.b(_1221_),
		.c(_1222_)
	);

	or_bb _1934_ (
		.a(_1222_),
		.b(new_net_626),
		.c(_1223_)
	);

	or_bi _1935_ (
		.a(new_net_2215),
		.b(_1125_),
		.c(_1224_)
	);

	or_bi _1936_ (
		.a(new_net_222),
		.b(new_net_2216),
		.c(_1225_)
	);

	or_ii _1937_ (
		.a(new_net_2217),
		.b(new_net_509),
		.c(_1226_)
	);

	and_bi _1938_ (
		.a(new_net_1574),
		.b(new_net_549),
		.c(_1227_)
	);

	inv _1939_ (
		.din(new_net_1453),
		.dout(_1228_)
	);

	and_bi _1940_ (
		.a(new_net_347),
		.b(new_net_36),
		.c(_1229_)
	);

	or_bi _1941_ (
		.a(new_net_861),
		.b(new_net_780),
		.c(_1230_)
	);

	and_bi _1942_ (
		.a(new_net_1202),
		.b(new_net_348),
		.c(_1231_)
	);

	or_bb _1943_ (
		.a(_1231_),
		.b(new_net_862),
		.c(_1232_)
	);

	and_ii _1944_ (
		.a(new_net_230),
		.b(new_net_37),
		.c(_1233_)
	);

	and_bi _1945_ (
		.a(new_net_2218),
		.b(_1233_),
		.c(_1234_)
	);

	and_bi _1946_ (
		.a(new_net_2219),
		.b(_1234_),
		.c(_1235_)
	);

	and_ii _1947_ (
		.a(new_net_34),
		.b(new_net_244),
		.c(_1236_)
	);

	and_bb _1948_ (
		.a(new_net_38),
		.b(new_net_248),
		.c(_1237_)
	);

	and_ii _1949_ (
		.a(_1237_),
		.b(_1236_),
		.c(_1238_)
	);

	or_bi _1950_ (
		.a(new_net_1507),
		.b(new_net_167),
		.c(_1239_)
	);

	and_bi _1951_ (
		.a(new_net_1508),
		.b(new_net_169),
		.c(_1240_)
	);

	and_bi _1952_ (
		.a(_1239_),
		.b(_1240_),
		.c(_1241_)
	);

	or_bb _1953_ (
		.a(new_net_2220),
		.b(new_net_1616),
		.c(_1242_)
	);

	and_bi _1954_ (
		.a(new_net_782),
		.b(new_net_326),
		.c(_1243_)
	);

	or_bb _1955_ (
		.a(_1243_),
		.b(new_net_60),
		.c(_1244_)
	);

	and_bi _1956_ (
		.a(new_net_1201),
		.b(new_net_247),
		.c(_1245_)
	);

	and_bi _1957_ (
		.a(new_net_245),
		.b(new_net_1199),
		.c(_1246_)
	);

	and_ii _1958_ (
		.a(_1246_),
		.b(_1245_),
		.c(_1247_)
	);

	or_bb _1959_ (
		.a(new_net_1631),
		.b(new_net_1331),
		.c(_0000_)
	);

	and_bb _1960_ (
		.a(new_net_1632),
		.b(new_net_1332),
		.c(_0001_)
	);

	and_bi _1961_ (
		.a(_0000_),
		.b(_0001_),
		.c(_0002_)
	);

	and_bi _1962_ (
		.a(new_net_1619),
		.b(new_net_2221),
		.c(_0003_)
	);

	and_bi _1963_ (
		.a(_1242_),
		.b(_0003_),
		.c(_0004_)
	);

	and_bi _1964_ (
		.a(new_net_599),
		.b(new_net_815),
		.c(_0005_)
	);

	and_bi _1965_ (
		.a(new_net_1347),
		.b(new_net_598),
		.c(_0006_)
	);

	and_ii _1966_ (
		.a(_0006_),
		.b(_0005_),
		.c(_0007_)
	);

	or_bi _1967_ (
		.a(new_net_555),
		.b(new_net_1190),
		.c(_0008_)
	);

	and_bi _1968_ (
		.a(new_net_1712),
		.b(new_net_2222),
		.c(_0009_)
	);

	and_ii _1969_ (
		.a(new_net_1714),
		.b(new_net_1191),
		.c(_0010_)
	);

	or_bb _1970_ (
		.a(new_net_2223),
		.b(new_net_192),
		.c(_0011_)
	);

	or_bb _1971_ (
		.a(_0011_),
		.b(new_net_2224),
		.c(_0012_)
	);

	or_bb _1972_ (
		.a(new_net_1452),
		.b(new_net_976),
		.c(_0013_)
	);

	and_bb _1973_ (
		.a(new_net_1449),
		.b(new_net_974),
		.c(_0014_)
	);

	and_bi _1974_ (
		.a(_0013_),
		.b(_0014_),
		.c(_0015_)
	);

	or_bb _1975_ (
		.a(new_net_775),
		.b(new_net_601),
		.c(_0016_)
	);

	and_bb _1976_ (
		.a(new_net_776),
		.b(new_net_602),
		.c(_0017_)
	);

	or_bi _1977_ (
		.a(_0017_),
		.b(_0016_),
		.c(_0018_)
	);

	or_bb _1978_ (
		.a(new_net_1058),
		.b(new_net_1182),
		.c(_0019_)
	);

	and_bi _1979_ (
		.a(new_net_1059),
		.b(new_net_1193),
		.c(_0020_)
	);

	and_bi _1980_ (
		.a(_0019_),
		.b(_0020_),
		.c(_0021_)
	);

	and_bi _1981_ (
		.a(new_net_788),
		.b(new_net_534),
		.c(_0022_)
	);

	and_bi _1982_ (
		.a(new_net_535),
		.b(new_net_789),
		.c(_0023_)
	);

	or_bb _1983_ (
		.a(_0023_),
		.b(_0022_),
		.c(_0024_)
	);

	and_ii _1984_ (
		.a(new_net_1324),
		.b(new_net_497),
		.c(_0025_)
	);

	and_bb _1985_ (
		.a(new_net_1325),
		.b(new_net_498),
		.c(_0026_)
	);

	or_bb _1986_ (
		.a(_0026_),
		.b(new_net_1219),
		.c(_0027_)
	);

	or_bb _1987_ (
		.a(_0027_),
		.b(new_net_2225),
		.c(_0028_)
	);

	and_bi _1988_ (
		.a(new_net_1371),
		.b(new_net_1269),
		.c(_0029_)
	);

	and_bi _1989_ (
		.a(new_net_1267),
		.b(new_net_981),
		.c(_0030_)
	);

	and_ii _1990_ (
		.a(_0030_),
		.b(_0029_),
		.c(_0031_)
	);

	and_ii _1991_ (
		.a(new_net_327),
		.b(new_net_688),
		.c(_0032_)
	);

	and_bb _1992_ (
		.a(new_net_328),
		.b(new_net_689),
		.c(_0033_)
	);

	or_bb _1993_ (
		.a(_0033_),
		.b(_0032_),
		.c(_0034_)
	);

	or_bb _1994_ (
		.a(new_net_1473),
		.b(new_net_985),
		.c(_0035_)
	);

	and_bi _1995_ (
		.a(new_net_1468),
		.b(new_net_1010),
		.c(_0036_)
	);

	and_bi _1996_ (
		.a(_0035_),
		.b(_0036_),
		.c(_0037_)
	);

	and_bi _1997_ (
		.a(new_net_1257),
		.b(_0037_),
		.c(_0038_)
	);

	or_ii _1998_ (
		.a(new_net_1474),
		.b(new_net_1051),
		.c(_0039_)
	);

	and_bi _1999_ (
		.a(new_net_1367),
		.b(new_net_1469),
		.c(_0040_)
	);

	and_bi _2000_ (
		.a(_0039_),
		.b(_0040_),
		.c(_0041_)
	);

	and_bi _2001_ (
		.a(new_net_1596),
		.b(_0041_),
		.c(_0042_)
	);

	and_ii _2002_ (
		.a(_0042_),
		.b(_0038_),
		.c(_0043_)
	);

	or_bi _2003_ (
		.a(new_net_241),
		.b(new_net_1487),
		.c(_0044_)
	);

	and_bi _2004_ (
		.a(new_net_242),
		.b(new_net_1488),
		.c(_0045_)
	);

	and_bi _2005_ (
		.a(_0044_),
		.b(_0045_),
		.c(_0046_)
	);

	or_bb _2006_ (
		.a(new_net_1663),
		.b(new_net_986),
		.c(_0047_)
	);

	and_bi _2007_ (
		.a(new_net_1658),
		.b(new_net_1011),
		.c(_0048_)
	);

	and_bi _2008_ (
		.a(_0047_),
		.b(_0048_),
		.c(_0049_)
	);

	and_bi _2009_ (
		.a(new_net_1593),
		.b(_0049_),
		.c(_0050_)
	);

	or_ii _2010_ (
		.a(new_net_1664),
		.b(new_net_1052),
		.c(_0051_)
	);

	and_bi _2011_ (
		.a(new_net_1368),
		.b(new_net_1659),
		.c(_0052_)
	);

	and_bi _2012_ (
		.a(_0051_),
		.b(_0052_),
		.c(_0053_)
	);

	and_bi _2013_ (
		.a(new_net_132),
		.b(_0053_),
		.c(_0054_)
	);

	or_bb _2014_ (
		.a(_0054_),
		.b(_0050_),
		.c(_0055_)
	);

	or_bb _2015_ (
		.a(new_net_1605),
		.b(new_net_990),
		.c(_0056_)
	);

	and_bi _2016_ (
		.a(new_net_1610),
		.b(new_net_1016),
		.c(_0057_)
	);

	and_bi _2017_ (
		.a(_0056_),
		.b(_0057_),
		.c(_0058_)
	);

	and_bi _2018_ (
		.a(new_net_1289),
		.b(_0058_),
		.c(_0059_)
	);

	or_ii _2019_ (
		.a(new_net_1606),
		.b(new_net_1044),
		.c(_0060_)
	);

	and_bi _2020_ (
		.a(new_net_1372),
		.b(new_net_1611),
		.c(_0061_)
	);

	and_bi _2021_ (
		.a(_0060_),
		.b(_0061_),
		.c(_0062_)
	);

	and_bi _2022_ (
		.a(new_net_1021),
		.b(_0062_),
		.c(_0063_)
	);

	or_bb _2023_ (
		.a(_0063_),
		.b(_0059_),
		.c(_0064_)
	);

	and_ii _2024_ (
		.a(new_net_39),
		.b(new_net_636),
		.c(_0065_)
	);

	and_bb _2025_ (
		.a(new_net_40),
		.b(new_net_637),
		.c(_0066_)
	);

	and_ii _2026_ (
		.a(_0066_),
		.b(_0065_),
		.c(_0067_)
	);

	or_bb _2027_ (
		.a(new_net_74),
		.b(new_net_495),
		.c(_0068_)
	);

	and_bb _2028_ (
		.a(new_net_75),
		.b(new_net_496),
		.c(_0069_)
	);

	and_bi _2029_ (
		.a(_0068_),
		.b(_0069_),
		.c(_0070_)
	);

	and_ii _2030_ (
		.a(new_net_1463),
		.b(new_net_844),
		.c(_0071_)
	);

	and_bb _2031_ (
		.a(new_net_1464),
		.b(new_net_843),
		.c(_0072_)
	);

	and_ii _2032_ (
		.a(new_net_2226),
		.b(new_net_287),
		.c(_0073_)
	);

	or_bi _2033_ (
		.a(new_net_485),
		.b(new_net_227),
		.c(_0074_)
	);

	and_bi _2034_ (
		.a(new_net_486),
		.b(new_net_225),
		.c(_0075_)
	);

	or_bi _2035_ (
		.a(new_net_2227),
		.b(new_net_218),
		.c(_0076_)
	);

	and_ii _2036_ (
		.a(new_net_739),
		.b(new_net_489),
		.c(_0077_)
	);

	and_bb _2037_ (
		.a(new_net_740),
		.b(new_net_490),
		.c(_0078_)
	);

	and_ii _2038_ (
		.a(_0078_),
		.b(_0077_),
		.c(_0079_)
	);

	or_bb _2039_ (
		.a(new_net_1028),
		.b(new_net_161),
		.c(_0080_)
	);

	and_bb _2040_ (
		.a(new_net_1029),
		.b(new_net_162),
		.c(_0081_)
	);

	or_bb _2041_ (
		.a(_0081_),
		.b(new_net_588),
		.c(_0082_)
	);

	and_bi _2042_ (
		.a(new_net_2228),
		.b(_0082_),
		.c(_0083_)
	);

	or_bb _2043_ (
		.a(_0083_),
		.b(new_net_622),
		.c(_0084_)
	);

	and_bi _2044_ (
		.a(_0028_),
		.b(new_net_2229),
		.c(_0085_)
	);

	and_bi _2045_ (
		.a(new_net_2230),
		.b(new_net_223),
		.c(_0086_)
	);

	or_bb _2046_ (
		.a(new_net_2231),
		.b(new_net_1715),
		.c(_0087_)
	);

	and_bi _2047_ (
		.a(new_net_658),
		.b(new_net_480),
		.c(_0088_)
	);

	or_bb _2048_ (
		.a(_0088_),
		.b(new_net_800),
		.c(_0089_)
	);

	or_bb _2049_ (
		.a(new_net_2232),
		.b(_1227_),
		.c(_0090_)
	);

	or_bb _2050_ (
		.a(new_net_664),
		.b(new_net_1454),
		.c(_0091_)
	);

	and_bi _2051_ (
		.a(new_net_1717),
		.b(new_net_568),
		.c(_0092_)
	);

	or_bi _2052_ (
		.a(new_net_1455),
		.b(new_net_665),
		.c(_0093_)
	);

	and_bi _2053_ (
		.a(new_net_1478),
		.b(new_net_760),
		.c(_0094_)
	);

	or_bb _2054_ (
		.a(_0094_),
		.b(_0092_),
		.c(_0095_)
	);

	and_bi _2055_ (
		.a(_0090_),
		.b(new_net_2233),
		.c(_0096_)
	);

	or_bb _2056_ (
		.a(_0096_),
		.b(new_net_1129),
		.c(new_net_2453)
	);

	inv _2057_ (
		.din(new_net_1493),
		.dout(_0097_)
	);

	and_bi _2058_ (
		.a(new_net_1153),
		.b(new_net_552),
		.c(_0098_)
	);

	inv _2059_ (
		.din(new_net_1532),
		.dout(_0099_)
	);

	and_bi _2060_ (
		.a(new_net_1500),
		.b(new_net_482),
		.c(_0100_)
	);

	or_bb _2061_ (
		.a(_0100_),
		.b(new_net_672),
		.c(_0101_)
	);

	or_bb _2062_ (
		.a(new_net_2234),
		.b(_0098_),
		.c(_0102_)
	);

	or_bb _2063_ (
		.a(new_net_1534),
		.b(new_net_1494),
		.c(_0103_)
	);

	and_bi _2064_ (
		.a(new_net_1718),
		.b(new_net_730),
		.c(_0104_)
	);

	or_bi _2065_ (
		.a(new_net_1533),
		.b(new_net_1495),
		.c(_0105_)
	);

	and_bi _2066_ (
		.a(new_net_1479),
		.b(new_net_299),
		.c(_0106_)
	);

	or_bb _2067_ (
		.a(_0106_),
		.b(_0104_),
		.c(_0107_)
	);

	and_bi _2068_ (
		.a(_0102_),
		.b(new_net_2235),
		.c(_0108_)
	);

	or_bb _2069_ (
		.a(_0108_),
		.b(new_net_1130),
		.c(new_net_2357)
	);

	and_bb _2070_ (
		.a(new_net_2236),
		.b(new_net_57),
		.c(new_net_2435)
	);

	and_ii _2071_ (
		.a(new_net_1636),
		.b(new_net_174),
		.c(_0109_)
	);

	and_bb _2072_ (
		.a(new_net_1638),
		.b(new_net_176),
		.c(_0110_)
	);

	and_ii _2073_ (
		.a(_0110_),
		.b(_0109_),
		.c(_0111_)
	);

	and_bi _2074_ (
		.a(new_net_1399),
		.b(new_net_1418),
		.c(_0112_)
	);

	and_bi _2075_ (
		.a(new_net_1415),
		.b(new_net_1395),
		.c(_0113_)
	);

	and_ii _2076_ (
		.a(_0113_),
		.b(_0112_),
		.c(_0114_)
	);

	and_ii _2077_ (
		.a(new_net_187),
		.b(new_net_139),
		.c(_0115_)
	);

	and_bb _2078_ (
		.a(new_net_188),
		.b(new_net_140),
		.c(_0116_)
	);

	and_ii _2079_ (
		.a(_0116_),
		.b(_0115_),
		.c(_0117_)
	);

	inv _2080_ (
		.din(_0117_),
		.dout(_0118_)
	);

	and_bi _2081_ (
		.a(new_net_1030),
		.b(new_net_851),
		.c(_0119_)
	);

	and_bi _2082_ (
		.a(new_net_853),
		.b(new_net_1034),
		.c(_0120_)
	);

	or_bb _2083_ (
		.a(_0120_),
		.b(_0119_),
		.c(_0121_)
	);

	and_bi _2084_ (
		.a(new_net_1475),
		.b(new_net_1159),
		.c(_0122_)
	);

	and_bi _2085_ (
		.a(new_net_1160),
		.b(new_net_1470),
		.c(_0123_)
	);

	and_ii _2086_ (
		.a(_0123_),
		.b(_0122_),
		.c(_0124_)
	);

	and_bi _2087_ (
		.a(new_net_1607),
		.b(new_net_1660),
		.c(_0125_)
	);

	and_bi _2088_ (
		.a(new_net_1665),
		.b(new_net_1612),
		.c(_0126_)
	);

	and_ii _2089_ (
		.a(_0126_),
		.b(_0125_),
		.c(_0127_)
	);

	and_bi _2090_ (
		.a(new_net_135),
		.b(new_net_394),
		.c(_0128_)
	);

	and_bi _2091_ (
		.a(new_net_395),
		.b(new_net_136),
		.c(_0129_)
	);

	and_ii _2092_ (
		.a(_0129_),
		.b(_0128_),
		.c(_0130_)
	);

	and_bi _2093_ (
		.a(new_net_493),
		.b(new_net_255),
		.c(_0131_)
	);

	and_bi _2094_ (
		.a(new_net_256),
		.b(new_net_494),
		.c(_0132_)
	);

	or_bb _2095_ (
		.a(_0132_),
		.b(_0131_),
		.c(new_net_15)
	);

	and_ii _2096_ (
		.a(new_net_841),
		.b(new_net_881),
		.c(_0133_)
	);

	and_bb _2097_ (
		.a(new_net_837),
		.b(new_net_876),
		.c(_0134_)
	);

	and_ii _2098_ (
		.a(_0134_),
		.b(_0133_),
		.c(_0135_)
	);

	and_bi _2099_ (
		.a(new_net_754),
		.b(new_net_956),
		.c(_0136_)
	);

	and_bi _2100_ (
		.a(new_net_961),
		.b(new_net_759),
		.c(_0137_)
	);

	and_ii _2101_ (
		.a(_0137_),
		.b(_0136_),
		.c(_0138_)
	);

	and_ii _2102_ (
		.a(new_net_1188),
		.b(new_net_566),
		.c(_0139_)
	);

	and_bb _2103_ (
		.a(new_net_1189),
		.b(new_net_567),
		.c(_0140_)
	);

	and_ii _2104_ (
		.a(_0140_),
		.b(_0139_),
		.c(_0141_)
	);

	and_ii _2105_ (
		.a(new_net_1070),
		.b(new_net_1141),
		.c(_0142_)
	);

	and_bb _2106_ (
		.a(new_net_1076),
		.b(new_net_1147),
		.c(_0143_)
	);

	and_ii _2107_ (
		.a(_0143_),
		.b(_0142_),
		.c(_0144_)
	);

	and_bi _2108_ (
		.a(new_net_1253),
		.b(new_net_1296),
		.c(_0145_)
	);

	and_bi _2109_ (
		.a(new_net_1297),
		.b(new_net_1248),
		.c(_0146_)
	);

	and_ii _2110_ (
		.a(_0146_),
		.b(_0145_),
		.c(_0147_)
	);

	and_bi _2111_ (
		.a(new_net_430),
		.b(new_net_703),
		.c(_0148_)
	);

	and_bi _2112_ (
		.a(new_net_704),
		.b(new_net_431),
		.c(_0149_)
	);

	or_bb _2113_ (
		.a(_0149_),
		.b(_0148_),
		.c(_0150_)
	);

	and_bi _2114_ (
		.a(new_net_1118),
		.b(new_net_1179),
		.c(_0151_)
	);

	and_bi _2115_ (
		.a(new_net_1173),
		.b(new_net_1112),
		.c(_0152_)
	);

	or_bb _2116_ (
		.a(_0152_),
		.b(_0151_),
		.c(_0153_)
	);

	and_ii _2117_ (
		.a(new_net_1127),
		.b(new_net_829),
		.c(_0154_)
	);

	and_bb _2118_ (
		.a(new_net_1128),
		.b(new_net_830),
		.c(_0155_)
	);

	and_ii _2119_ (
		.a(_0155_),
		.b(_0154_),
		.c(_0156_)
	);

	and_ii _2120_ (
		.a(new_net_921),
		.b(new_net_1460),
		.c(_0157_)
	);

	and_bb _2121_ (
		.a(new_net_922),
		.b(new_net_1461),
		.c(_0158_)
	);

	and_ii _2122_ (
		.a(_0158_),
		.b(_0157_),
		.c(_0159_)
	);

	inv _2123_ (
		.din(new_net_80),
		.dout(new_net_2411)
	);

	and_ii _2124_ (
		.a(new_net_683),
		.b(new_net_308),
		.c(_0160_)
	);

	and_bb _2125_ (
		.a(new_net_684),
		.b(new_net_307),
		.c(_0161_)
	);

	or_bb _2126_ (
		.a(_0161_),
		.b(_0160_),
		.c(_0162_)
	);

	or_bb _2127_ (
		.a(new_net_396),
		.b(new_net_168),
		.c(_0163_)
	);

	and_bb _2128_ (
		.a(new_net_397),
		.b(new_net_170),
		.c(_0164_)
	);

	and_bi _2129_ (
		.a(_0163_),
		.b(_0164_),
		.c(_0165_)
	);

	and_bb _2130_ (
		.a(new_net_852),
		.b(new_net_1522),
		.c(_0166_)
	);

	and_bi _2131_ (
		.a(new_net_2237),
		.b(new_net_1526),
		.c(_0167_)
	);

	and_ii _2132_ (
		.a(_0167_),
		.b(_0166_),
		.c(_0168_)
	);

	and_bi _2133_ (
		.a(new_net_62),
		.b(new_net_1093),
		.c(_0169_)
	);

	and_bi _2134_ (
		.a(new_net_1092),
		.b(new_net_64),
		.c(_0170_)
	);

	and_ii _2135_ (
		.a(_0170_),
		.b(_0169_),
		.c(_0171_)
	);

	and_bi _2136_ (
		.a(new_net_886),
		.b(new_net_1316),
		.c(_0172_)
	);

	and_bi _2137_ (
		.a(new_net_1317),
		.b(new_net_887),
		.c(_0173_)
	);

	or_bb _2138_ (
		.a(_0173_),
		.b(_0172_),
		.c(_0174_)
	);

	and_ii _2139_ (
		.a(new_net_1686),
		.b(new_net_1120),
		.c(_0175_)
	);

	and_bi _2140_ (
		.a(new_net_1621),
		.b(new_net_1388),
		.c(_0176_)
	);

	and_ii _2141_ (
		.a(new_net_2238),
		.b(_0175_),
		.c(_0177_)
	);

	and_bi _2142_ (
		.a(new_net_193),
		.b(new_net_105),
		.c(_0178_)
	);

	and_bi _2143_ (
		.a(new_net_106),
		.b(new_net_194),
		.c(_0179_)
	);

	or_bb _2144_ (
		.a(_0179_),
		.b(_0178_),
		.c(_0180_)
	);

	and_ii _2145_ (
		.a(new_net_1441),
		.b(new_net_1363),
		.c(_0181_)
	);

	and_bb _2146_ (
		.a(new_net_1442),
		.b(new_net_1364),
		.c(_0182_)
	);

	and_ii _2147_ (
		.a(_0182_),
		.b(_0181_),
		.c(_0183_)
	);

	and_bi _2148_ (
		.a(new_net_1184),
		.b(new_net_1535),
		.c(_0184_)
	);

	and_bi _2149_ (
		.a(new_net_1536),
		.b(new_net_1185),
		.c(_0185_)
	);

	or_bb _2150_ (
		.a(_0185_),
		.b(_0184_),
		.c(_0186_)
	);

	inv _2151_ (
		.din(new_net_1024),
		.dout(new_net_2505)
	);

	or_bb _2152_ (
		.a(new_net_264),
		.b(new_net_316),
		.c(_0187_)
	);

	and_bb _2153_ (
		.a(new_net_263),
		.b(new_net_315),
		.c(_0188_)
	);

	and_bi _2154_ (
		.a(_0187_),
		.b(_0188_),
		.c(_0189_)
	);

	and_bi _2155_ (
		.a(new_net_537),
		.b(new_net_203),
		.c(_0190_)
	);

	and_bi _2156_ (
		.a(new_net_204),
		.b(new_net_538),
		.c(_0191_)
	);

	and_ii _2157_ (
		.a(_0191_),
		.b(_0190_),
		.c(_0192_)
	);

	or_bi _2158_ (
		.a(new_net_1699),
		.b(new_net_180),
		.c(_0193_)
	);

	and_bi _2159_ (
		.a(new_net_1700),
		.b(new_net_181),
		.c(_0194_)
	);

	and_bi _2160_ (
		.a(_0193_),
		.b(_0194_),
		.c(_0195_)
	);

	and_ii _2161_ (
		.a(new_net_501),
		.b(new_net_1567),
		.c(_0196_)
	);

	and_bb _2162_ (
		.a(new_net_502),
		.b(new_net_1565),
		.c(_0197_)
	);

	and_ii _2163_ (
		.a(_0197_),
		.b(_0196_),
		.c(_0198_)
	);

	and_bb _2164_ (
		.a(new_net_1563),
		.b(new_net_1298),
		.c(_0199_)
	);

	and_bi _2165_ (
		.a(new_net_2239),
		.b(new_net_1560),
		.c(_0200_)
	);

	and_ii _2166_ (
		.a(_0200_),
		.b(_0199_),
		.c(_0201_)
	);

	and_bi _2167_ (
		.a(new_net_232),
		.b(new_net_159),
		.c(_0202_)
	);

	and_bi _2168_ (
		.a(new_net_160),
		.b(new_net_233),
		.c(_0203_)
	);

	or_bb _2169_ (
		.a(_0203_),
		.b(_0202_),
		.c(_0204_)
	);

	or_ii _2170_ (
		.a(new_net_778),
		.b(new_net_785),
		.c(_0205_)
	);

	and_bi _2171_ (
		.a(new_net_1384),
		.b(new_net_786),
		.c(_0206_)
	);

	and_bi _2172_ (
		.a(_0205_),
		.b(_0206_),
		.c(_0207_)
	);

	and_ii _2173_ (
		.a(new_net_1681),
		.b(new_net_291),
		.c(_0208_)
	);

	and_bb _2174_ (
		.a(new_net_1682),
		.b(new_net_292),
		.c(_0209_)
	);

	and_ii _2175_ (
		.a(_0209_),
		.b(_0208_),
		.c(_0210_)
	);

	and_ii _2176_ (
		.a(new_net_444),
		.b(new_net_189),
		.c(_0211_)
	);

	and_bb _2177_ (
		.a(new_net_445),
		.b(new_net_190),
		.c(_0212_)
	);

	and_ii _2178_ (
		.a(_0212_),
		.b(_0211_),
		.c(_0213_)
	);

	or_bb _2179_ (
		.a(new_net_545),
		.b(new_net_137),
		.c(_0214_)
	);

	and_bb _2180_ (
		.a(new_net_546),
		.b(new_net_138),
		.c(_0215_)
	);

	and_bi _2181_ (
		.a(_0214_),
		.b(_0215_),
		.c(new_net_16)
	);

	and_bb _2182_ (
		.a(new_net_1405),
		.b(new_net_209),
		.c(new_net_14)
	);

	and_bb _2183_ (
		.a(new_net_2240),
		.b(new_net_1275),
		.c(new_net_2367)
	);

	and_bi _2184_ (
		.a(new_net_2241),
		.b(new_net_1627),
		.c(new_net_2393)
	);

	or_bi _2185_ (
		.a(new_net_1306),
		.b(new_net_2242),
		.c(_0216_)
	);

	and_bb _2186_ (
		.a(new_net_2243),
		.b(new_net_1312),
		.c(_0217_)
	);

	or_bb _2187_ (
		.a(new_net_2244),
		.b(new_net_909),
		.c(_0218_)
	);

	and_bi _2188_ (
		.a(new_net_2245),
		.b(_0218_),
		.c(_0219_)
	);

	and_bi _2189_ (
		.a(new_net_1273),
		.b(_0219_),
		.c(new_net_2399)
	);

	or_bi _2190_ (
		.a(new_net_1313),
		.b(new_net_2246),
		.c(_0220_)
	);

	and_bb _2191_ (
		.a(new_net_2247),
		.b(new_net_1307),
		.c(_0221_)
	);

	or_bb _2192_ (
		.a(new_net_2248),
		.b(new_net_915),
		.c(_0222_)
	);

	and_bi _2193_ (
		.a(new_net_2249),
		.b(_0222_),
		.c(_0223_)
	);

	and_bi _2194_ (
		.a(new_net_1278),
		.b(_0223_),
		.c(new_net_2503)
	);

	or_bi _2195_ (
		.a(new_net_1308),
		.b(new_net_2250),
		.c(_0224_)
	);

	and_bb _2196_ (
		.a(new_net_2251),
		.b(new_net_1314),
		.c(_0225_)
	);

	or_bb _2197_ (
		.a(new_net_2252),
		.b(new_net_910),
		.c(_0226_)
	);

	and_bi _2198_ (
		.a(new_net_2253),
		.b(_0226_),
		.c(_0227_)
	);

	and_bi _2199_ (
		.a(new_net_1274),
		.b(_0227_),
		.c(new_net_2459)
	);

	or_bi _2200_ (
		.a(new_net_1315),
		.b(new_net_2254),
		.c(_0228_)
	);

	and_bb _2201_ (
		.a(new_net_2255),
		.b(new_net_1309),
		.c(_0229_)
	);

	or_bb _2202_ (
		.a(new_net_2256),
		.b(new_net_916),
		.c(_0230_)
	);

	and_bi _2203_ (
		.a(new_net_2257),
		.b(_0230_),
		.c(_0231_)
	);

	and_bi _2204_ (
		.a(new_net_1279),
		.b(_0231_),
		.c(new_net_2477)
	);

	or_bb _2205_ (
		.a(new_net_1336),
		.b(new_net_687),
		.c(_0232_)
	);

	or_bb _2206_ (
		.a(new_net_2258),
		.b(new_net_219),
		.c(_0233_)
	);

	or_bb _2207_ (
		.a(_0233_),
		.b(new_net_443),
		.c(_0234_)
	);

	or_bb _2208_ (
		.a(new_net_654),
		.b(new_net_172),
		.c(_0235_)
	);

	or_bb _2209_ (
		.a(new_net_2259),
		.b(_0234_),
		.c(_0236_)
	);

	and_bi _2210_ (
		.a(new_net_288),
		.b(_0236_),
		.c(new_net_2447)
	);

	and_ii _2211_ (
		.a(new_net_695),
		.b(new_net_504),
		.c(_0237_)
	);

	and_bi _2212_ (
		.a(_0237_),
		.b(new_net_1057),
		.c(_0238_)
	);

	or_bb _2213_ (
		.a(new_net_950),
		.b(new_net_846),
		.c(_0239_)
	);

	or_bb _2214_ (
		.a(new_net_737),
		.b(new_net_926),
		.c(_0240_)
	);

	or_bb _2215_ (
		.a(new_net_1081),
		.b(new_net_1428),
		.c(_0241_)
	);

	or_bb _2216_ (
		.a(_0241_),
		.b(_0240_),
		.c(_0242_)
	);

	or_bb _2217_ (
		.a(_0242_),
		.b(new_net_2260),
		.c(_0243_)
	);

	and_bi _2218_ (
		.a(new_net_2261),
		.b(_0243_),
		.c(new_net_2499)
	);

	or_bi _2219_ (
		.a(new_net_1158),
		.b(new_net_1443),
		.c(_0244_)
	);

	and_ii _2220_ (
		.a(new_net_1285),
		.b(new_net_533),
		.c(new_net_2371)
	);

	and_ii _2221_ (
		.a(new_net_1448),
		.b(new_net_330),
		.c(_0245_)
	);

	or_ii _2222_ (
		.a(new_net_2262),
		.b(new_net_254),
		.c(_0246_)
	);

	and_bi _2223_ (
		.a(new_net_1263),
		.b(new_net_293),
		.c(new_net_2425)
	);

	and_bi _2224_ (
		.a(new_net_411),
		.b(new_net_1287),
		.c(_0247_)
	);

	and_ii _2225_ (
		.a(new_net_1580),
		.b(new_net_850),
		.c(_0248_)
	);

	or_bb _2226_ (
		.a(_0248_),
		.b(new_net_1390),
		.c(_0249_)
	);

	or_bb _2227_ (
		.a(new_net_354),
		.b(new_net_317),
		.c(new_net_2373)
	);

	or_bi _2228_ (
		.a(new_net_311),
		.b(new_net_250),
		.c(new_net_2443)
	);

	inv _2229_ (
		.din(new_net_146),
		.dout(_0250_)
	);

	or_ii _2230_ (
		.a(new_net_423),
		.b(new_net_382),
		.c(_0251_)
	);

	inv _2231_ (
		.din(new_net_141),
		.dout(_0252_)
	);

	and_bi _2232_ (
		.a(new_net_582),
		.b(new_net_384),
		.c(_0253_)
	);

	or_bb _2233_ (
		.a(_0253_),
		.b(new_net_432),
		.c(_0254_)
	);

	and_bi _2234_ (
		.a(_0251_),
		.b(new_net_2263),
		.c(_0255_)
	);

	or_bi _2235_ (
		.a(new_net_143),
		.b(new_net_147),
		.c(_0256_)
	);

	and_bi _2236_ (
		.a(new_net_505),
		.b(new_net_714),
		.c(_0257_)
	);

	or_bb _2237_ (
		.a(new_net_142),
		.b(new_net_149),
		.c(_0258_)
	);

	and_bi _2238_ (
		.a(new_net_352),
		.b(new_net_514),
		.c(_0259_)
	);

	or_bb _2239_ (
		.a(_0259_),
		.b(_0257_),
		.c(_0260_)
	);

	or_bb _2240_ (
		.a(new_net_2264),
		.b(_0255_),
		.c(new_net_2509)
	);

	or_bi _2241_ (
		.a(new_net_927),
		.b(new_net_420),
		.c(_0261_)
	);

	inv _2242_ (
		.din(new_net_1087),
		.dout(_0262_)
	);

	and_bb _2243_ (
		.a(new_net_580),
		.b(new_net_937),
		.c(_0263_)
	);

	or_bb _2244_ (
		.a(_0263_),
		.b(new_net_1357),
		.c(_0264_)
	);

	and_bi _2245_ (
		.a(_0261_),
		.b(new_net_2265),
		.c(_0265_)
	);

	or_bi _2246_ (
		.a(new_net_1089),
		.b(new_net_929),
		.c(_0266_)
	);

	and_bi _2247_ (
		.a(new_net_506),
		.b(new_net_643),
		.c(_0267_)
	);

	or_bb _2248_ (
		.a(new_net_1088),
		.b(new_net_947),
		.c(_0268_)
	);

	and_bi _2249_ (
		.a(new_net_353),
		.b(new_net_268),
		.c(_0269_)
	);

	or_bb _2250_ (
		.a(_0269_),
		.b(_0267_),
		.c(_0270_)
	);

	or_bb _2251_ (
		.a(new_net_2266),
		.b(_0265_),
		.c(new_net_2451)
	);

	or_bb _2252_ (
		.a(new_net_42),
		.b(new_net_1027),
		.c(_0271_)
	);

	or_bb _2253_ (
		.a(new_net_2267),
		.b(new_net_1281),
		.c(_0272_)
	);

	or_bb _2254_ (
		.a(_0272_),
		.b(new_net_1704),
		.c(_0273_)
	);

	or_bb _2255_ (
		.a(_0273_),
		.b(new_net_774),
		.c(_0274_)
	);

	or_bb _2256_ (
		.a(new_net_2268),
		.b(new_net_83),
		.c(_0275_)
	);

	and_bi _2257_ (
		.a(new_net_1720),
		.b(new_net_2269),
		.c(_0276_)
	);

	or_bb _2258_ (
		.a(new_net_1598),
		.b(new_net_1162),
		.c(_0277_)
	);

	and_bi _2259_ (
		.a(_0276_),
		.b(_0277_),
		.c(new_net_2417)
	);

	or_bi _2260_ (
		.a(new_net_719),
		.b(new_net_1167),
		.c(_0278_)
	);

	or_bb _2261_ (
		.a(new_net_2270),
		.b(new_net_217),
		.c(_0279_)
	);

	or_bb _2262_ (
		.a(new_net_2271),
		.b(new_net_492),
		.c(_0280_)
	);

	or_bb _2263_ (
		.a(new_net_2272),
		.b(new_net_235),
		.c(_0281_)
	);

	or_bb _2264_ (
		.a(new_net_2273),
		.b(new_net_563),
		.c(_0282_)
	);

	or_bb _2265_ (
		.a(new_net_2274),
		.b(new_net_351),
		.c(_0283_)
	);

	and_ii _2266_ (
		.a(new_net_2275),
		.b(new_net_402),
		.c(_0284_)
	);

	and_bi _2267_ (
		.a(_0284_),
		.b(new_net_164),
		.c(new_net_2469)
	);

	and_bi _2268_ (
		.a(new_net_422),
		.b(new_net_663),
		.c(_0285_)
	);

	and_bi _2269_ (
		.a(new_net_578),
		.b(new_net_1569),
		.c(_0286_)
	);

	or_bb _2270_ (
		.a(_0286_),
		.b(new_net_801),
		.c(_0287_)
	);

	or_bb _2271_ (
		.a(new_net_2276),
		.b(_0285_),
		.c(_0288_)
	);

	and_bi _2272_ (
		.a(new_net_1583),
		.b(new_net_569),
		.c(_0289_)
	);

	and_bi _2273_ (
		.a(new_net_1542),
		.b(new_net_767),
		.c(_0290_)
	);

	or_bb _2274_ (
		.a(_0290_),
		.b(_0289_),
		.c(_0291_)
	);

	and_bi _2275_ (
		.a(_0288_),
		.b(new_net_2277),
		.c(_0292_)
	);

	and_bi _2276_ (
		.a(new_net_107),
		.b(_0292_),
		.c(new_net_2427)
	);

	and_bi _2277_ (
		.a(new_net_424),
		.b(new_net_1501),
		.c(_0293_)
	);

	and_bi _2278_ (
		.a(new_net_579),
		.b(new_net_1148),
		.c(_0294_)
	);

	or_bb _2279_ (
		.a(_0294_),
		.b(new_net_677),
		.c(_0295_)
	);

	or_bb _2280_ (
		.a(new_net_2278),
		.b(_0293_),
		.c(_0296_)
	);

	and_bi _2281_ (
		.a(new_net_1584),
		.b(new_net_731),
		.c(_0297_)
	);

	and_bi _2282_ (
		.a(new_net_1543),
		.b(new_net_295),
		.c(_0298_)
	);

	or_bb _2283_ (
		.a(_0298_),
		.b(_0297_),
		.c(_0299_)
	);

	and_bi _2284_ (
		.a(_0296_),
		.b(new_net_2279),
		.c(_0300_)
	);

	and_bi _2285_ (
		.a(new_net_112),
		.b(_0300_),
		.c(new_net_2397)
	);

	or_ii _2286_ (
		.a(new_net_321),
		.b(new_net_376),
		.c(_0301_)
	);

	and_bi _2287_ (
		.a(new_net_416),
		.b(new_net_383),
		.c(_0302_)
	);

	or_bb _2288_ (
		.a(_0302_),
		.b(new_net_434),
		.c(_0303_)
	);

	and_bi _2289_ (
		.a(_0301_),
		.b(_0303_),
		.c(_0304_)
	);

	and_bi _2290_ (
		.a(new_net_1476),
		.b(new_net_708),
		.c(_0305_)
	);

	and_bi _2291_ (
		.a(new_net_1022),
		.b(new_net_515),
		.c(_0306_)
	);

	or_bb _2292_ (
		.a(_0306_),
		.b(_0305_),
		.c(_0307_)
	);

	or_bb _2293_ (
		.a(new_net_2280),
		.b(_0304_),
		.c(new_net_2437)
	);

	or_ii _2294_ (
		.a(new_net_894),
		.b(new_net_377),
		.c(_0308_)
	);

	and_bi _2295_ (
		.a(new_net_1086),
		.b(new_net_385),
		.c(_0309_)
	);

	or_bb _2296_ (
		.a(_0309_),
		.b(new_net_433),
		.c(_0310_)
	);

	and_bi _2297_ (
		.a(_0308_),
		.b(new_net_2281),
		.c(_0311_)
	);

	and_bi _2298_ (
		.a(new_net_1064),
		.b(new_net_511),
		.c(_0312_)
	);

	and_bi _2299_ (
		.a(new_net_790),
		.b(new_net_715),
		.c(_0313_)
	);

	or_bb _2300_ (
		.a(_0313_),
		.b(_0312_),
		.c(_0314_)
	);

	or_bb _2301_ (
		.a(new_net_2282),
		.b(_0311_),
		.c(new_net_2501)
	);

	or_ii _2302_ (
		.a(new_net_31),
		.b(new_net_378),
		.c(_0315_)
	);

	and_bi _2303_ (
		.a(new_net_186),
		.b(new_net_386),
		.c(_0316_)
	);

	or_bb _2304_ (
		.a(_0316_),
		.b(new_net_436),
		.c(_0317_)
	);

	and_bi _2305_ (
		.a(_0315_),
		.b(new_net_2283),
		.c(_0318_)
	);

	and_bi _2306_ (
		.a(new_net_450),
		.b(new_net_710),
		.c(_0319_)
	);

	and_bi _2307_ (
		.a(new_net_882),
		.b(new_net_517),
		.c(_0320_)
	);

	or_bb _2308_ (
		.a(_0320_),
		.b(_0319_),
		.c(_0321_)
	);

	or_bb _2309_ (
		.a(new_net_2284),
		.b(_0318_),
		.c(new_net_2383)
	);

	or_ii _2310_ (
		.a(new_net_1123),
		.b(new_net_379),
		.c(_0322_)
	);

	and_bi _2311_ (
		.a(new_net_823),
		.b(new_net_387),
		.c(_0323_)
	);

	or_bb _2312_ (
		.a(_0323_),
		.b(new_net_435),
		.c(_0324_)
	);

	and_bi _2313_ (
		.a(_0322_),
		.b(new_net_2285),
		.c(_0325_)
	);

	and_bi _2314_ (
		.a(new_net_403),
		.b(new_net_709),
		.c(_0326_)
	);

	and_bi _2315_ (
		.a(new_net_593),
		.b(new_net_516),
		.c(_0327_)
	);

	or_bb _2316_ (
		.a(_0327_),
		.b(_0326_),
		.c(_0328_)
	);

	or_bb _2317_ (
		.a(new_net_2286),
		.b(_0325_),
		.c(new_net_2369)
	);

	or_bi _2318_ (
		.a(new_net_938),
		.b(new_net_322),
		.c(_0329_)
	);

	and_bb _2319_ (
		.a(new_net_418),
		.b(new_net_933),
		.c(_0330_)
	);

	or_bb _2320_ (
		.a(_0330_),
		.b(new_net_1348),
		.c(_0331_)
	);

	and_bi _2321_ (
		.a(_0329_),
		.b(_0331_),
		.c(_0332_)
	);

	and_bi _2322_ (
		.a(new_net_1023),
		.b(new_net_269),
		.c(_0333_)
	);

	and_bi _2323_ (
		.a(new_net_1477),
		.b(new_net_649),
		.c(_0334_)
	);

	or_bb _2324_ (
		.a(_0334_),
		.b(_0333_),
		.c(_0335_)
	);

	or_bb _2325_ (
		.a(new_net_2287),
		.b(_0332_),
		.c(new_net_2473)
	);

	or_bi _2326_ (
		.a(new_net_942),
		.b(new_net_895),
		.c(_0336_)
	);

	and_bb _2327_ (
		.a(new_net_1085),
		.b(new_net_930),
		.c(_0337_)
	);

	or_bb _2328_ (
		.a(_0337_),
		.b(new_net_1349),
		.c(_0338_)
	);

	and_bi _2329_ (
		.a(_0336_),
		.b(new_net_2288),
		.c(_0339_)
	);

	and_bi _2330_ (
		.a(new_net_791),
		.b(new_net_645),
		.c(_0340_)
	);

	and_bi _2331_ (
		.a(new_net_1065),
		.b(new_net_274),
		.c(_0341_)
	);

	or_bb _2332_ (
		.a(_0341_),
		.b(_0340_),
		.c(_0342_)
	);

	or_bb _2333_ (
		.a(new_net_2289),
		.b(_0339_),
		.c(new_net_2467)
	);

	or_bi _2334_ (
		.a(new_net_939),
		.b(new_net_29),
		.c(_0343_)
	);

	and_bb _2335_ (
		.a(new_net_183),
		.b(new_net_934),
		.c(_0344_)
	);

	or_bb _2336_ (
		.a(_0344_),
		.b(new_net_1351),
		.c(_0345_)
	);

	and_bi _2337_ (
		.a(_0343_),
		.b(new_net_2290),
		.c(_0346_)
	);

	and_bi _2338_ (
		.a(new_net_883),
		.b(new_net_270),
		.c(_0347_)
	);

	and_bi _2339_ (
		.a(new_net_451),
		.b(new_net_650),
		.c(_0348_)
	);

	or_bb _2340_ (
		.a(_0348_),
		.b(_0347_),
		.c(_0349_)
	);

	or_bb _2341_ (
		.a(new_net_2291),
		.b(_0346_),
		.c(new_net_2481)
	);

	or_bi _2342_ (
		.a(new_net_940),
		.b(new_net_1124),
		.c(_0350_)
	);

	and_bb _2343_ (
		.a(new_net_824),
		.b(new_net_935),
		.c(_0351_)
	);

	or_bb _2344_ (
		.a(_0351_),
		.b(new_net_1350),
		.c(_0352_)
	);

	and_bi _2345_ (
		.a(_0350_),
		.b(new_net_2292),
		.c(_0353_)
	);

	and_bi _2346_ (
		.a(new_net_404),
		.b(new_net_644),
		.c(_0354_)
	);

	and_bi _2347_ (
		.a(new_net_594),
		.b(new_net_273),
		.c(_0355_)
	);

	or_bb _2348_ (
		.a(_0355_),
		.b(_0354_),
		.c(_0356_)
	);

	or_bb _2349_ (
		.a(new_net_2293),
		.b(_0353_),
		.c(new_net_2365)
	);

	and_bi _2350_ (
		.a(new_net_323),
		.b(new_net_659),
		.c(_0357_)
	);

	and_bi _2351_ (
		.a(new_net_419),
		.b(new_net_1576),
		.c(_0358_)
	);

	or_bb _2352_ (
		.a(_0358_),
		.b(new_net_797),
		.c(_0359_)
	);

	or_bb _2353_ (
		.a(_0359_),
		.b(_0357_),
		.c(_0360_)
	);

	and_bi _2354_ (
		.a(new_net_1425),
		.b(new_net_570),
		.c(_0361_)
	);

	and_bi _2355_ (
		.a(new_net_808),
		.b(new_net_768),
		.c(_0362_)
	);

	or_bb _2356_ (
		.a(_0362_),
		.b(_0361_),
		.c(_0363_)
	);

	and_bi _2357_ (
		.a(_0360_),
		.b(new_net_2294),
		.c(_0364_)
	);

	and_bi _2358_ (
		.a(new_net_117),
		.b(_0364_),
		.c(new_net_2461)
	);

	and_bi _2359_ (
		.a(new_net_1125),
		.b(new_net_666),
		.c(_0365_)
	);

	and_bi _2360_ (
		.a(new_net_821),
		.b(new_net_1568),
		.c(_0366_)
	);

	or_bb _2361_ (
		.a(_0366_),
		.b(new_net_802),
		.c(_0367_)
	);

	or_bb _2362_ (
		.a(new_net_2295),
		.b(_0365_),
		.c(_0368_)
	);

	and_bi _2363_ (
		.a(new_net_1385),
		.b(new_net_573),
		.c(_0369_)
	);

	and_bi _2364_ (
		.a(new_net_413),
		.b(new_net_761),
		.c(_0370_)
	);

	or_bb _2365_ (
		.a(_0370_),
		.b(_0369_),
		.c(_0371_)
	);

	and_bi _2366_ (
		.a(_0368_),
		.b(new_net_2296),
		.c(_0372_)
	);

	and_bi _2367_ (
		.a(new_net_125),
		.b(_0372_),
		.c(new_net_2407)
	);

	and_bi _2368_ (
		.a(new_net_32),
		.b(new_net_660),
		.c(_0373_)
	);

	and_bi _2369_ (
		.a(new_net_184),
		.b(new_net_1575),
		.c(_0374_)
	);

	or_bb _2370_ (
		.a(_0374_),
		.b(new_net_796),
		.c(_0375_)
	);

	or_bb _2371_ (
		.a(new_net_2297),
		.b(_0373_),
		.c(_0376_)
	);

	and_bi _2372_ (
		.a(new_net_745),
		.b(new_net_571),
		.c(_0377_)
	);

	and_bi _2373_ (
		.a(new_net_1358),
		.b(new_net_766),
		.c(_0378_)
	);

	or_bb _2374_ (
		.a(_0378_),
		.b(_0377_),
		.c(_0379_)
	);

	and_bi _2375_ (
		.a(_0376_),
		.b(new_net_2298),
		.c(_0380_)
	);

	and_bi _2376_ (
		.a(new_net_108),
		.b(_0380_),
		.c(new_net_2413)
	);

	and_bi _2377_ (
		.a(new_net_897),
		.b(new_net_667),
		.c(_0381_)
	);

	and_bi _2378_ (
		.a(new_net_1083),
		.b(new_net_1570),
		.c(_0382_)
	);

	or_bb _2379_ (
		.a(_0382_),
		.b(new_net_803),
		.c(_0383_)
	);

	or_bb _2380_ (
		.a(new_net_2299),
		.b(_0381_),
		.c(_0384_)
	);

	and_bi _2381_ (
		.a(new_net_1302),
		.b(new_net_574),
		.c(_0385_)
	);

	and_bi _2382_ (
		.a(new_net_1322),
		.b(new_net_762),
		.c(_0386_)
	);

	or_bb _2383_ (
		.a(_0386_),
		.b(_0385_),
		.c(_0387_)
	);

	and_bi _2384_ (
		.a(_0384_),
		.b(new_net_2300),
		.c(_0388_)
	);

	and_bi _2385_ (
		.a(new_net_113),
		.b(_0388_),
		.c(new_net_2387)
	);

	and_bi _2386_ (
		.a(new_net_320),
		.b(new_net_1496),
		.c(_0389_)
	);

	and_bi _2387_ (
		.a(new_net_417),
		.b(new_net_1155),
		.c(_0390_)
	);

	or_bb _2388_ (
		.a(_0390_),
		.b(new_net_674),
		.c(_0391_)
	);

	or_bb _2389_ (
		.a(_0391_),
		.b(_0389_),
		.c(_0392_)
	);

	and_bi _2390_ (
		.a(new_net_1426),
		.b(new_net_725),
		.c(_0393_)
	);

	and_bi _2391_ (
		.a(new_net_809),
		.b(new_net_301),
		.c(_0394_)
	);

	or_bb _2392_ (
		.a(_0394_),
		.b(_0393_),
		.c(_0395_)
	);

	and_bi _2393_ (
		.a(_0392_),
		.b(new_net_2301),
		.c(_0396_)
	);

	and_bi _2394_ (
		.a(new_net_118),
		.b(_0396_),
		.c(new_net_2445)
	);

	and_bi _2395_ (
		.a(new_net_1126),
		.b(new_net_1502),
		.c(_0397_)
	);

	and_bi _2396_ (
		.a(new_net_820),
		.b(new_net_1149),
		.c(_0398_)
	);

	or_bb _2397_ (
		.a(_0398_),
		.b(new_net_678),
		.c(_0399_)
	);

	or_bb _2398_ (
		.a(new_net_2302),
		.b(_0397_),
		.c(_0400_)
	);

	and_bi _2399_ (
		.a(new_net_1386),
		.b(new_net_732),
		.c(_0401_)
	);

	and_bi _2400_ (
		.a(new_net_414),
		.b(new_net_296),
		.c(_0402_)
	);

	or_bb _2401_ (
		.a(_0402_),
		.b(_0401_),
		.c(_0403_)
	);

	and_bi _2402_ (
		.a(_0400_),
		.b(new_net_2303),
		.c(_0404_)
	);

	and_bi _2403_ (
		.a(new_net_126),
		.b(_0404_),
		.c(new_net_2475)
	);

	and_bi _2404_ (
		.a(new_net_30),
		.b(new_net_1497),
		.c(_0405_)
	);

	and_bi _2405_ (
		.a(new_net_185),
		.b(new_net_1154),
		.c(_0406_)
	);

	or_bb _2406_ (
		.a(_0406_),
		.b(new_net_673),
		.c(_0407_)
	);

	or_bb _2407_ (
		.a(new_net_2304),
		.b(_0405_),
		.c(_0408_)
	);

	and_bi _2408_ (
		.a(new_net_746),
		.b(new_net_726),
		.c(_0409_)
	);

	and_bi _2409_ (
		.a(new_net_1359),
		.b(new_net_300),
		.c(_0410_)
	);

	or_bb _2410_ (
		.a(_0410_),
		.b(_0409_),
		.c(_0411_)
	);

	and_bi _2411_ (
		.a(_0408_),
		.b(new_net_2305),
		.c(_0412_)
	);

	and_bi _2412_ (
		.a(new_net_109),
		.b(_0412_),
		.c(new_net_2431)
	);

	and_bi _2413_ (
		.a(new_net_896),
		.b(new_net_1503),
		.c(_0413_)
	);

	and_bi _2414_ (
		.a(new_net_1082),
		.b(new_net_1150),
		.c(_0414_)
	);

	or_bb _2415_ (
		.a(_0414_),
		.b(new_net_679),
		.c(_0415_)
	);

	or_bb _2416_ (
		.a(new_net_2306),
		.b(_0413_),
		.c(_0416_)
	);

	and_bi _2417_ (
		.a(new_net_1303),
		.b(new_net_733),
		.c(_0417_)
	);

	and_bi _2418_ (
		.a(new_net_1323),
		.b(new_net_297),
		.c(_0418_)
	);

	or_bb _2419_ (
		.a(_0418_),
		.b(_0417_),
		.c(_0419_)
	);

	and_bi _2420_ (
		.a(_0416_),
		.b(new_net_2307),
		.c(_0420_)
	);

	and_bi _2421_ (
		.a(new_net_114),
		.b(_0420_),
		.c(new_net_2471)
	);

	or_ii _2422_ (
		.a(new_net_1164),
		.b(new_net_589),
		.c(_0421_)
	);

	and_ii _2423_ (
		.a(new_net_251),
		.b(new_net_1101),
		.c(_0422_)
	);

	and_bb _2424_ (
		.a(new_net_246),
		.b(new_net_1102),
		.c(_0423_)
	);

	and_ii _2425_ (
		.a(_0423_),
		.b(_0422_),
		.c(_0424_)
	);

	and_bi _2426_ (
		.a(new_net_1326),
		.b(new_net_592),
		.c(_0425_)
	);

	and_bi _2427_ (
		.a(_0421_),
		.b(new_net_2308),
		.c(_0426_)
	);

	and_bi _2428_ (
		.a(new_net_129),
		.b(_0426_),
		.c(_0427_)
	);

	or_ii _2429_ (
		.a(G178),
		.b(G62),
		.c(_0428_)
	);

	or_bi _2430_ (
		.a(new_net_907),
		.b(new_net_590),
		.c(_0429_)
	);

	and_ii _2431_ (
		.a(new_net_226),
		.b(new_net_591),
		.c(_0430_)
	);

	and_bi _2432_ (
		.a(new_net_2309),
		.b(_0430_),
		.c(_0431_)
	);

	or_bb _2433_ (
		.a(_0431_),
		.b(new_net_130),
		.c(_0432_)
	);

	or_ii _2434_ (
		.a(_0432_),
		.b(new_net_2310),
		.c(_0433_)
	);

	and_ii _2435_ (
		.a(new_net_2311),
		.b(_0427_),
		.c(new_net_2485)
	);

	and_bi _2436_ (
		.a(new_net_1166),
		.b(new_net_1327),
		.c(_0434_)
	);

	and_bi _2437_ (
		.a(new_net_1328),
		.b(new_net_1168),
		.c(_0435_)
	);

	or_bb _2438_ (
		.a(_0435_),
		.b(_0434_),
		.c(new_net_2377)
	);

	or_ii _2439_ (
		.a(new_net_1401),
		.b(new_net_1440),
		.c(_0436_)
	);

	and_ii _2440_ (
		.a(_0436_),
		.b(new_net_748),
		.c(_0437_)
	);

	and_bb _2441_ (
		.a(_0437_),
		.b(new_net_860),
		.c(_0438_)
	);

	or_ii _2442_ (
		.a(new_net_2312),
		.b(new_net_1000),
		.c(_0439_)
	);

	or_bb _2443_ (
		.a(_0439_),
		.b(new_net_81),
		.c(_0440_)
	);

	or_bb _2444_ (
		.a(new_net_2313),
		.b(new_net_1025),
		.c(_0441_)
	);

	and_bi _2445_ (
		.a(new_net_1334),
		.b(_0441_),
		.c(new_net_2423)
	);

	or_bi _2446_ (
		.a(new_net_943),
		.b(new_net_1481),
		.c(_0442_)
	);

	and_bb _2447_ (
		.a(new_net_1642),
		.b(new_net_936),
		.c(_0443_)
	);

	or_bb _2448_ (
		.a(_0443_),
		.b(new_net_1352),
		.c(_0444_)
	);

	and_bi _2449_ (
		.a(_0442_),
		.b(new_net_2314),
		.c(_0445_)
	);

	and_bi _2450_ (
		.a(new_net_692),
		.b(new_net_271),
		.c(_0446_)
	);

	and_bi _2451_ (
		.a(new_net_794),
		.b(new_net_651),
		.c(_0447_)
	);

	or_bb _2452_ (
		.a(_0447_),
		.b(_0446_),
		.c(_0448_)
	);

	or_bb _2453_ (
		.a(new_net_2315),
		.b(_0445_),
		.c(new_net_2439)
	);

	or_ii _2454_ (
		.a(new_net_1482),
		.b(new_net_380),
		.c(_0449_)
	);

	and_bi _2455_ (
		.a(new_net_1643),
		.b(new_net_388),
		.c(_0450_)
	);

	or_bb _2456_ (
		.a(_0450_),
		.b(new_net_437),
		.c(_0451_)
	);

	and_bi _2457_ (
		.a(_0449_),
		.b(new_net_2316),
		.c(_0452_)
	);

	and_bi _2458_ (
		.a(new_net_693),
		.b(new_net_512),
		.c(_0453_)
	);

	and_bi _2459_ (
		.a(new_net_795),
		.b(new_net_716),
		.c(_0454_)
	);

	or_bb _2460_ (
		.a(_0454_),
		.b(_0453_),
		.c(_0455_)
	);

	or_bb _2461_ (
		.a(new_net_2317),
		.b(_0452_),
		.c(new_net_2401)
	);

	or_ii _2462_ (
		.a(new_net_238),
		.b(new_net_148),
		.c(_0456_)
	);

	and_bi _2463_ (
		.a(new_net_428),
		.b(new_net_152),
		.c(_0457_)
	);

	or_bb _2464_ (
		.a(_0457_),
		.b(new_net_438),
		.c(_0458_)
	);

	and_bi _2465_ (
		.a(new_net_2318),
		.b(_0458_),
		.c(_0459_)
	);

	and_bi _2466_ (
		.a(new_net_523),
		.b(new_net_711),
		.c(_0460_)
	);

	and_bi _2467_ (
		.a(new_net_1489),
		.b(new_net_518),
		.c(_0461_)
	);

	or_bb _2468_ (
		.a(_0461_),
		.b(_0460_),
		.c(_0462_)
	);

	or_bb _2469_ (
		.a(new_net_2319),
		.b(_0459_),
		.c(new_net_2355)
	);

	or_bb _2470_ (
		.a(new_net_888),
		.b(new_net_381),
		.c(_0463_)
	);

	and_bi _2471_ (
		.a(new_net_968),
		.b(new_net_153),
		.c(_0464_)
	);

	or_bb _2472_ (
		.a(_0464_),
		.b(new_net_439),
		.c(_0465_)
	);

	and_bi _2473_ (
		.a(new_net_2320),
		.b(_0465_),
		.c(_0466_)
	);

	and_bi _2474_ (
		.a(new_net_468),
		.b(new_net_712),
		.c(_0467_)
	);

	and_bi _2475_ (
		.a(new_net_696),
		.b(new_net_519),
		.c(_0468_)
	);

	or_bb _2476_ (
		.a(_0468_),
		.b(_0467_),
		.c(_0469_)
	);

	or_bb _2477_ (
		.a(new_net_2321),
		.b(_0466_),
		.c(new_net_2457)
	);

	or_ii _2478_ (
		.a(new_net_283),
		.b(new_net_150),
		.c(_0470_)
	);

	and_bi _2479_ (
		.a(new_net_858),
		.b(new_net_154),
		.c(_0471_)
	);

	or_bb _2480_ (
		.a(_0471_),
		.b(new_net_440),
		.c(_0472_)
	);

	and_bi _2481_ (
		.a(new_net_2322),
		.b(_0472_),
		.c(_0473_)
	);

	and_bi _2482_ (
		.a(new_net_165),
		.b(new_net_713),
		.c(_0474_)
	);

	and_bi _2483_ (
		.a(new_net_1458),
		.b(new_net_520),
		.c(_0475_)
	);

	or_bb _2484_ (
		.a(_0475_),
		.b(_0474_),
		.c(_0476_)
	);

	or_bb _2485_ (
		.a(new_net_2323),
		.b(_0473_),
		.c(new_net_2483)
	);

	or_bi _2486_ (
		.a(new_net_944),
		.b(new_net_425),
		.c(_0477_)
	);

	and_bb _2487_ (
		.a(new_net_240),
		.b(new_net_931),
		.c(_0478_)
	);

	or_bb _2488_ (
		.a(_0478_),
		.b(new_net_1353),
		.c(_0479_)
	);

	and_bi _2489_ (
		.a(_0477_),
		.b(_0479_),
		.c(_0480_)
	);

	and_bi _2490_ (
		.a(new_net_524),
		.b(new_net_646),
		.c(_0481_)
	);

	and_bi _2491_ (
		.a(new_net_1490),
		.b(new_net_275),
		.c(_0482_)
	);

	or_bb _2492_ (
		.a(_0482_),
		.b(_0481_),
		.c(_0483_)
	);

	or_bb _2493_ (
		.a(new_net_2324),
		.b(_0480_),
		.c(new_net_2479)
	);

	or_bi _2494_ (
		.a(new_net_941),
		.b(new_net_965),
		.c(_0484_)
	);

	and_bi _2495_ (
		.a(new_net_948),
		.b(new_net_891),
		.c(_0485_)
	);

	or_bb _2496_ (
		.a(_0485_),
		.b(new_net_1354),
		.c(_0486_)
	);

	and_bi _2497_ (
		.a(_0484_),
		.b(_0486_),
		.c(_0487_)
	);

	and_bi _2498_ (
		.a(new_net_469),
		.b(new_net_647),
		.c(_0488_)
	);

	and_bi _2499_ (
		.a(new_net_697),
		.b(new_net_276),
		.c(_0489_)
	);

	or_bb _2500_ (
		.a(_0489_),
		.b(_0488_),
		.c(_0490_)
	);

	or_bb _2501_ (
		.a(new_net_2325),
		.b(_0487_),
		.c(new_net_2405)
	);

	or_bi _2502_ (
		.a(new_net_945),
		.b(new_net_855),
		.c(_0491_)
	);

	and_bb _2503_ (
		.a(new_net_286),
		.b(new_net_932),
		.c(_0492_)
	);

	or_bb _2504_ (
		.a(_0492_),
		.b(new_net_1355),
		.c(_0493_)
	);

	and_bi _2505_ (
		.a(_0491_),
		.b(_0493_),
		.c(_0494_)
	);

	and_bi _2506_ (
		.a(new_net_166),
		.b(new_net_648),
		.c(_0495_)
	);

	and_bi _2507_ (
		.a(new_net_1459),
		.b(new_net_277),
		.c(_0496_)
	);

	or_bb _2508_ (
		.a(_0496_),
		.b(_0495_),
		.c(_0497_)
	);

	or_bb _2509_ (
		.a(new_net_2326),
		.b(_0494_),
		.c(new_net_2511)
	);

	and_bi _2510_ (
		.a(new_net_284),
		.b(new_net_1571),
		.c(_0498_)
	);

	and_bi _2511_ (
		.a(new_net_857),
		.b(new_net_668),
		.c(_0499_)
	);

	or_bb _2512_ (
		.a(_0499_),
		.b(new_net_798),
		.c(_0500_)
	);

	or_bb _2513_ (
		.a(_0500_),
		.b(new_net_2327),
		.c(_0501_)
	);

	and_bi _2514_ (
		.a(new_net_1437),
		.b(new_net_572),
		.c(_0502_)
	);

	and_bi _2515_ (
		.a(new_net_816),
		.b(new_net_769),
		.c(_0503_)
	);

	or_bb _2516_ (
		.a(_0503_),
		.b(_0502_),
		.c(_0504_)
	);

	and_bi _2517_ (
		.a(_0501_),
		.b(new_net_2328),
		.c(_0505_)
	);

	and_bi _2518_ (
		.a(new_net_119),
		.b(_0505_),
		.c(new_net_2361)
	);

	and_bi _2519_ (
		.a(new_net_669),
		.b(new_net_892),
		.c(_0506_)
	);

	and_bi _2520_ (
		.a(new_net_966),
		.b(new_net_661),
		.c(_0507_)
	);

	or_bb _2521_ (
		.a(_0507_),
		.b(new_net_804),
		.c(_0508_)
	);

	or_bb _2522_ (
		.a(_0508_),
		.b(new_net_2329),
		.c(_0509_)
	);

	and_bi _2523_ (
		.a(new_net_1421),
		.b(new_net_575),
		.c(_0510_)
	);

	and_bi _2524_ (
		.a(new_net_1705),
		.b(new_net_763),
		.c(_0511_)
	);

	or_bb _2525_ (
		.a(_0511_),
		.b(_0510_),
		.c(_0512_)
	);

	and_bi _2526_ (
		.a(_0509_),
		.b(new_net_2330),
		.c(_0513_)
	);

	and_bi _2527_ (
		.a(new_net_123),
		.b(_0513_),
		.c(new_net_2381)
	);

	and_bi _2528_ (
		.a(new_net_237),
		.b(new_net_1572),
		.c(_0514_)
	);

	and_bi _2529_ (
		.a(new_net_427),
		.b(new_net_670),
		.c(_0515_)
	);

	or_bb _2530_ (
		.a(_0515_),
		.b(new_net_799),
		.c(_0516_)
	);

	or_bb _2531_ (
		.a(_0516_),
		.b(new_net_2331),
		.c(_0517_)
	);

	and_bi _2532_ (
		.a(new_net_1653),
		.b(new_net_764),
		.c(_0518_)
	);

	and_bi _2533_ (
		.a(new_net_1135),
		.b(new_net_576),
		.c(_0519_)
	);

	or_bb _2534_ (
		.a(_0519_),
		.b(_0518_),
		.c(_0520_)
	);

	and_bi _2535_ (
		.a(_0517_),
		.b(new_net_2332),
		.c(_0521_)
	);

	and_bi _2536_ (
		.a(new_net_110),
		.b(_0521_),
		.c(new_net_2395)
	);

	and_bi _2537_ (
		.a(new_net_1484),
		.b(new_net_671),
		.c(_0522_)
	);

	and_bi _2538_ (
		.a(new_net_1640),
		.b(new_net_1573),
		.c(_0523_)
	);

	or_bb _2539_ (
		.a(_0523_),
		.b(new_net_805),
		.c(_0524_)
	);

	or_bb _2540_ (
		.a(new_net_2333),
		.b(_0522_),
		.c(_0525_)
	);

	and_bi _2541_ (
		.a(new_net_1391),
		.b(new_net_577),
		.c(_0526_)
	);

	and_bi _2542_ (
		.a(new_net_1622),
		.b(new_net_765),
		.c(_0527_)
	);

	or_bb _2543_ (
		.a(_0527_),
		.b(_0526_),
		.c(_0528_)
	);

	and_bi _2544_ (
		.a(_0525_),
		.b(new_net_2334),
		.c(_0529_)
	);

	and_bi _2545_ (
		.a(new_net_115),
		.b(_0529_),
		.c(new_net_2449)
	);

	and_bi _2546_ (
		.a(new_net_854),
		.b(new_net_1498),
		.c(_0530_)
	);

	and_bi _2547_ (
		.a(new_net_285),
		.b(new_net_1156),
		.c(_0531_)
	);

	or_bb _2548_ (
		.a(_0531_),
		.b(new_net_675),
		.c(_0532_)
	);

	or_bb _2549_ (
		.a(_0532_),
		.b(_0530_),
		.c(_0533_)
	);

	and_bi _2550_ (
		.a(new_net_1438),
		.b(new_net_727),
		.c(_0534_)
	);

	and_bi _2551_ (
		.a(new_net_817),
		.b(new_net_302),
		.c(_0535_)
	);

	or_bb _2552_ (
		.a(_0535_),
		.b(_0534_),
		.c(_0536_)
	);

	and_bi _2553_ (
		.a(_0533_),
		.b(new_net_2335),
		.c(_0537_)
	);

	and_bi _2554_ (
		.a(new_net_120),
		.b(_0537_),
		.c(new_net_2491)
	);

	and_bi _2555_ (
		.a(new_net_969),
		.b(new_net_1504),
		.c(_0538_)
	);

	and_bi _2556_ (
		.a(new_net_1499),
		.b(new_net_889),
		.c(_0539_)
	);

	or_bb _2557_ (
		.a(_0539_),
		.b(new_net_680),
		.c(_0540_)
	);

	or_bb _2558_ (
		.a(_0540_),
		.b(_0538_),
		.c(_0541_)
	);

	and_bi _2559_ (
		.a(new_net_1706),
		.b(new_net_303),
		.c(_0542_)
	);

	and_bi _2560_ (
		.a(new_net_1422),
		.b(new_net_728),
		.c(_0543_)
	);

	or_bb _2561_ (
		.a(_0543_),
		.b(_0542_),
		.c(_0544_)
	);

	and_bi _2562_ (
		.a(_0541_),
		.b(new_net_2336),
		.c(_0545_)
	);

	and_bi _2563_ (
		.a(new_net_124),
		.b(_0545_),
		.c(new_net_2493)
	);

	and_bi _2564_ (
		.a(new_net_239),
		.b(new_net_1151),
		.c(_0546_)
	);

	and_bi _2565_ (
		.a(new_net_429),
		.b(new_net_1505),
		.c(_0547_)
	);

	or_bb _2566_ (
		.a(_0547_),
		.b(new_net_676),
		.c(_0548_)
	);

	or_bb _2567_ (
		.a(_0548_),
		.b(new_net_2337),
		.c(_0549_)
	);

	and_bi _2568_ (
		.a(new_net_1136),
		.b(new_net_729),
		.c(_0550_)
	);

	and_bi _2569_ (
		.a(new_net_1654),
		.b(new_net_304),
		.c(_0551_)
	);

	or_bb _2570_ (
		.a(_0551_),
		.b(_0550_),
		.c(_0552_)
	);

	and_bi _2571_ (
		.a(_0549_),
		.b(new_net_2338),
		.c(_0553_)
	);

	and_bi _2572_ (
		.a(new_net_111),
		.b(_0553_),
		.c(new_net_2363)
	);

	and_bi _2573_ (
		.a(new_net_1483),
		.b(new_net_1506),
		.c(_0554_)
	);

	and_bi _2574_ (
		.a(new_net_1639),
		.b(new_net_1152),
		.c(_0555_)
	);

	or_bb _2575_ (
		.a(_0555_),
		.b(new_net_681),
		.c(_0556_)
	);

	or_bb _2576_ (
		.a(new_net_2339),
		.b(_0554_),
		.c(_0557_)
	);

	and_bi _2577_ (
		.a(new_net_1392),
		.b(new_net_734),
		.c(_0558_)
	);

	and_bi _2578_ (
		.a(new_net_1623),
		.b(new_net_298),
		.c(_0559_)
	);

	or_bb _2579_ (
		.a(_0559_),
		.b(_0558_),
		.c(_0560_)
	);

	and_bi _2580_ (
		.a(_0557_),
		.b(new_net_2340),
		.c(_0561_)
	);

	and_bi _2581_ (
		.a(new_net_116),
		.b(_0561_),
		.c(new_net_2391)
	);

	or_bb _2582_ (
		.a(new_net_100),
		.b(new_net_2341),
		.c(_0562_)
	);

	and_bi _2583_ (
		.a(new_net_2342),
		.b(new_net_1716),
		.c(new_net_2353)
	);

	and_ii _2584_ (
		.a(new_net_87),
		.b(new_net_2343),
		.c(_0563_)
	);

	and_bi _2585_ (
		.a(new_net_510),
		.b(new_net_2344),
		.c(new_net_2409)
	);

	or_bb _2586_ (
		.a(new_net_551),
		.b(new_net_151),
		.c(_0564_)
	);

	and_bi _2587_ (
		.a(new_net_155),
		.b(new_net_481),
		.c(_0565_)
	);

	or_bb _2588_ (
		.a(_0565_),
		.b(new_net_441),
		.c(_0566_)
	);

	and_bi _2589_ (
		.a(_0564_),
		.b(new_net_2345),
		.c(_0567_)
	);

	and_bi _2590_ (
		.a(new_net_374),
		.b(new_net_513),
		.c(_0568_)
	);

	and_bi _2591_ (
		.a(new_net_525),
		.b(new_net_717),
		.c(_0569_)
	);

	or_bb _2592_ (
		.a(_0569_),
		.b(_0568_),
		.c(_0570_)
	);

	or_bb _2593_ (
		.a(new_net_2346),
		.b(_0567_),
		.c(new_net_2489)
	);

	or_bb _2594_ (
		.a(new_net_550),
		.b(new_net_928),
		.c(_0571_)
	);

	and_bi _2595_ (
		.a(new_net_946),
		.b(new_net_483),
		.c(_0572_)
	);

	or_bb _2596_ (
		.a(_0572_),
		.b(new_net_1356),
		.c(_0573_)
	);

	and_bi _2597_ (
		.a(_0571_),
		.b(new_net_2347),
		.c(_0574_)
	);

	and_bi _2598_ (
		.a(new_net_375),
		.b(new_net_272),
		.c(_0575_)
	);

	and_bi _2599_ (
		.a(new_net_526),
		.b(new_net_652),
		.c(_0576_)
	);

	or_bb _2600_ (
		.a(_0576_),
		.b(_0575_),
		.c(_0577_)
	);

	or_bb _2601_ (
		.a(new_net_2348),
		.b(_0574_),
		.c(new_net_2349)
	);

	and_bi _2602_ (
		.a(new_net_1264),
		.b(new_net_294),
		.c(new_net_2433)
	);

	and_ii _2603_ (
		.a(new_net_1286),
		.b(new_net_531),
		.c(new_net_2421)
	);

	or_bb _2604_ (
		.a(new_net_355),
		.b(new_net_318),
		.c(new_net_2385)
	);

	or_bi _2605_ (
		.a(new_net_312),
		.b(new_net_252),
		.c(new_net_2497)
	);

	spl2 new_net_1788_v_fanout (
		.a(new_net_1788),
		.b(G5219),
		.c(G5217)
	);

	spl4L _1226__v_fanout (
		.a(_1226_),
		.b(new_net_552),
		.c(new_net_551),
		.d(new_net_550),
		.e(new_net_549)
	);

	spl2 _1224__v_fanout (
		.a(_1224_),
		.b(new_net_509),
		.c(new_net_510)
	);

	bfr new_net_2513_bfr_before (
		.din(new_net_2513),
		.dout(G5291)
	);

	bfr new_net_2514_bfr_before (
		.din(new_net_2514),
		.dout(new_net_2513)
	);

	bfr new_net_2515_bfr_before (
		.din(new_net_2515),
		.dout(new_net_2514)
	);

	bfr new_net_2516_bfr_before (
		.din(new_net_2516),
		.dout(new_net_2515)
	);

	bfr new_net_2517_bfr_before (
		.din(new_net_2517),
		.dout(new_net_2516)
	);

	bfr new_net_2518_bfr_before (
		.din(new_net_2518),
		.dout(new_net_2517)
	);

	bfr new_net_2519_bfr_before (
		.din(new_net_2519),
		.dout(new_net_2518)
	);

	spl2 new_net_2103_v_fanout (
		.a(new_net_2103),
		.b(new_net_429),
		.c(new_net_2519)
	);

	bfr new_net_2520_bfr_before (
		.din(new_net_2520),
		.dout(G5214)
	);

	bfr new_net_2521_bfr_before (
		.din(new_net_2521),
		.dout(new_net_2520)
	);

	bfr new_net_2522_bfr_before (
		.din(new_net_2522),
		.dout(new_net_2521)
	);

	spl3L new_net_1861_v_fanout (
		.a(new_net_1861),
		.b(new_net_111),
		.c(new_net_110),
		.d(new_net_2522)
	);

	spl2 new_net_2105_v_fanout (
		.a(new_net_2105),
		.b(new_net_1483),
		.c(new_net_1481)
	);

	spl2 new_net_2101_v_fanout (
		.a(new_net_2101),
		.b(new_net_968),
		.c(new_net_969)
	);

	spl3L new_net_2104_v_fanout (
		.a(new_net_2104),
		.b(new_net_427),
		.c(new_net_428),
		.d(new_net_425)
	);

	bfr new_net_2523_bfr_before (
		.din(new_net_2523),
		.dout(G5290)
	);

	bfr new_net_2524_bfr_before (
		.din(new_net_2524),
		.dout(new_net_2523)
	);

	bfr new_net_2525_bfr_before (
		.din(new_net_2525),
		.dout(new_net_2524)
	);

	bfr new_net_2526_bfr_before (
		.din(new_net_2526),
		.dout(new_net_2525)
	);

	bfr new_net_2527_bfr_before (
		.din(new_net_2527),
		.dout(new_net_2526)
	);

	bfr new_net_2528_bfr_before (
		.din(new_net_2528),
		.dout(new_net_2527)
	);

	bfr new_net_2529_bfr_before (
		.din(new_net_2529),
		.dout(new_net_2528)
	);

	spl3L new_net_2106_v_fanout (
		.a(new_net_2106),
		.b(new_net_2529),
		.c(new_net_1484),
		.d(new_net_1482)
	);

	bfr new_net_2530_bfr_before (
		.din(new_net_2530),
		.dout(new_net_123)
	);

	spl2 new_net_1860_v_fanout (
		.a(new_net_1860),
		.b(new_net_2530),
		.c(new_net_124)
	);

	bfr new_net_2531_bfr_before (
		.din(new_net_2531),
		.dout(G5292)
	);

	bfr new_net_2532_bfr_before (
		.din(new_net_2532),
		.dout(new_net_2531)
	);

	bfr new_net_2533_bfr_before (
		.din(new_net_2533),
		.dout(new_net_2532)
	);

	bfr new_net_2534_bfr_before (
		.din(new_net_2534),
		.dout(new_net_2533)
	);

	bfr new_net_2535_bfr_before (
		.din(new_net_2535),
		.dout(new_net_2534)
	);

	bfr new_net_2536_bfr_before (
		.din(new_net_2536),
		.dout(new_net_2535)
	);

	bfr new_net_2537_bfr_before (
		.din(new_net_2537),
		.dout(new_net_2536)
	);

	spl3L new_net_2102_v_fanout (
		.a(new_net_2102),
		.b(new_net_965),
		.c(new_net_2537),
		.d(new_net_966)
	);

	spl2 new_net_21_v_fanout (
		.a(new_net_21),
		.b(new_net_2101),
		.c(new_net_2102)
	);

	spl2 new_net_20_v_fanout (
		.a(new_net_20),
		.b(new_net_2104),
		.c(new_net_2103)
	);

	spl3L new_net_2100_v_fanout (
		.a(new_net_2100),
		.b(new_net_888),
		.c(new_net_890),
		.d(new_net_889)
	);

	bfr new_net_2538_bfr_before (
		.din(new_net_2538),
		.dout(G5286)
	);

	bfr new_net_2539_bfr_before (
		.din(new_net_2539),
		.dout(new_net_2538)
	);

	bfr new_net_2540_bfr_before (
		.din(new_net_2540),
		.dout(new_net_2539)
	);

	bfr new_net_2541_bfr_before (
		.din(new_net_2541),
		.dout(new_net_2540)
	);

	bfr new_net_2542_bfr_before (
		.din(new_net_2542),
		.dout(new_net_2541)
	);

	bfr new_net_2543_bfr_before (
		.din(new_net_2543),
		.dout(new_net_2542)
	);

	bfr new_net_2544_bfr_before (
		.din(new_net_2544),
		.dout(new_net_2543)
	);

	bfr new_net_2545_bfr_before (
		.din(new_net_2545),
		.dout(new_net_2544)
	);

	spl3L new_net_2098_v_fanout (
		.a(new_net_2098),
		.b(new_net_2545),
		.c(new_net_239),
		.d(new_net_240)
	);

	bfr new_net_2546_bfr_before (
		.din(new_net_2546),
		.dout(new_net_1861)
	);

	bfr new_net_2547_bfr_before (
		.din(new_net_2547),
		.dout(new_net_115)
	);

	bfr new_net_2548_bfr_before (
		.din(new_net_2548),
		.dout(new_net_116)
	);

	spl4L new_net_1859_v_fanout (
		.a(new_net_1859),
		.b(new_net_2547),
		.c(new_net_2548),
		.d(new_net_1860),
		.e(new_net_2546)
	);

	spl2 new_net_2097_v_fanout (
		.a(new_net_2097),
		.b(new_net_237),
		.c(new_net_238)
	);

	spl2 new_net_2099_v_fanout (
		.a(new_net_2099),
		.b(new_net_892),
		.c(new_net_891)
	);

	spl2 new_net_17_v_fanout (
		.a(new_net_17),
		.b(new_net_2105),
		.c(new_net_2106)
	);

	bfr new_net_2549_bfr_before (
		.din(new_net_2549),
		.dout(new_net_680)
	);

	spl2 new_net_1966_v_fanout (
		.a(new_net_1966),
		.b(new_net_672),
		.c(new_net_2549)
	);

	spl2 new_net_19_v_fanout (
		.a(new_net_19),
		.b(new_net_2098),
		.c(new_net_2097)
	);

	bfr new_net_2550_bfr_before (
		.din(new_net_2550),
		.dout(new_net_1353)
	);

	bfr new_net_2551_bfr_before (
		.din(new_net_2551),
		.dout(new_net_1354)
	);

	spl3L new_net_1958_v_fanout (
		.a(new_net_1958),
		.b(new_net_2550),
		.c(new_net_2551),
		.d(new_net_1356)
	);

	spl2 _0910__v_fanout (
		.a(_0910_),
		.b(new_net_2100),
		.c(new_net_2099)
	);

	spl4L _0087__v_fanout (
		.a(_0087_),
		.b(new_net_482),
		.c(new_net_481),
		.d(new_net_483),
		.e(new_net_480)
	);

	bfr new_net_2552_bfr_before (
		.din(new_net_2552),
		.dout(G5293)
	);

	bfr new_net_2553_bfr_before (
		.din(new_net_2553),
		.dout(new_net_2552)
	);

	bfr new_net_2554_bfr_before (
		.din(new_net_2554),
		.dout(new_net_2553)
	);

	bfr new_net_2555_bfr_before (
		.din(new_net_2555),
		.dout(new_net_2554)
	);

	bfr new_net_2556_bfr_before (
		.din(new_net_2556),
		.dout(new_net_2555)
	);

	bfr new_net_2557_bfr_before (
		.din(new_net_2557),
		.dout(new_net_2556)
	);

	bfr new_net_2558_bfr_before (
		.din(new_net_2558),
		.dout(new_net_2557)
	);

	bfr new_net_2559_bfr_before (
		.din(new_net_2559),
		.dout(new_net_2558)
	);

	bfr new_net_2560_bfr_before (
		.din(new_net_2560),
		.dout(new_net_2559)
	);

	bfr new_net_2561_bfr_before (
		.din(new_net_2561),
		.dout(new_net_2560)
	);

	spl2 new_net_2095_v_fanout (
		.a(new_net_2095),
		.b(new_net_2561),
		.c(new_net_855)
	);

	spl3L new_net_2096_v_fanout (
		.a(new_net_2096),
		.b(new_net_854),
		.c(new_net_857),
		.d(new_net_858)
	);

	bfr new_net_2562_bfr_before (
		.din(new_net_2562),
		.dout(new_net_804)
	);

	bfr new_net_2563_bfr_before (
		.din(new_net_2563),
		.dout(new_net_2562)
	);

	bfr new_net_2564_bfr_before (
		.din(new_net_2564),
		.dout(new_net_799)
	);

	bfr new_net_2565_bfr_before (
		.din(new_net_2565),
		.dout(new_net_2564)
	);

	spl3L new_net_1973_v_fanout (
		.a(new_net_1973),
		.b(new_net_2563),
		.c(new_net_800),
		.d(new_net_2565)
	);

	bfr new_net_2566_bfr_before (
		.din(new_net_2566),
		.dout(new_net_1153)
	);

	bfr new_net_2567_bfr_before (
		.din(new_net_2567),
		.dout(new_net_2566)
	);

	bfr new_net_2568_bfr_before (
		.din(new_net_2568),
		.dout(new_net_2567)
	);

	spl2 new_net_1948_v_fanout (
		.a(new_net_1948),
		.b(new_net_1151),
		.c(new_net_2568)
	);

	bfr new_net_2569_bfr_before (
		.din(new_net_2569),
		.dout(new_net_438)
	);

	bfr new_net_2570_bfr_before (
		.din(new_net_2570),
		.dout(new_net_2569)
	);

	bfr new_net_2571_bfr_before (
		.din(new_net_2571),
		.dout(new_net_439)
	);

	bfr new_net_2572_bfr_before (
		.din(new_net_2572),
		.dout(new_net_2571)
	);

	spl3L new_net_1932_v_fanout (
		.a(new_net_1932),
		.b(new_net_2570),
		.c(new_net_2572),
		.d(new_net_441)
	);

	bfr new_net_2573_bfr_before (
		.din(new_net_2573),
		.dout(new_net_1574)
	);

	bfr new_net_2574_bfr_before (
		.din(new_net_2574),
		.dout(new_net_2573)
	);

	bfr new_net_2575_bfr_before (
		.din(new_net_2575),
		.dout(new_net_2574)
	);

	spl2 new_net_1988_v_fanout (
		.a(new_net_1988),
		.b(new_net_1572),
		.c(new_net_2575)
	);

	bfr new_net_2576_bfr_before (
		.din(new_net_2576),
		.dout(new_net_1499)
	);

	spl2 new_net_1900_v_fanout (
		.a(new_net_1900),
		.b(new_net_1500),
		.c(new_net_2576)
	);

	bfr new_net_2577_bfr_before (
		.din(new_net_2577),
		.dout(new_net_676)
	);

	bfr new_net_2578_bfr_before (
		.din(new_net_2578),
		.dout(new_net_2577)
	);

	bfr new_net_2579_bfr_before (
		.din(new_net_2579),
		.dout(new_net_2578)
	);

	spl2 new_net_1965_v_fanout (
		.a(new_net_1965),
		.b(new_net_1966),
		.c(new_net_2579)
	);

	bfr new_net_2580_bfr_before (
		.din(new_net_2580),
		.dout(new_net_119)
	);

	bfr new_net_2581_bfr_before (
		.din(new_net_2581),
		.dout(new_net_1859)
	);

	spl3L new_net_1858_v_fanout (
		.a(new_net_1858),
		.b(new_net_120),
		.c(new_net_2580),
		.d(new_net_2581)
	);

	bfr new_net_2582_bfr_before (
		.din(new_net_2582),
		.dout(G5288)
	);

	bfr new_net_2583_bfr_before (
		.din(new_net_2583),
		.dout(new_net_2582)
	);

	bfr new_net_2584_bfr_before (
		.din(new_net_2584),
		.dout(new_net_2583)
	);

	bfr new_net_2585_bfr_before (
		.din(new_net_2585),
		.dout(new_net_2584)
	);

	bfr new_net_2586_bfr_before (
		.din(new_net_2586),
		.dout(new_net_2585)
	);

	bfr new_net_2587_bfr_before (
		.din(new_net_2587),
		.dout(new_net_2586)
	);

	bfr new_net_2588_bfr_before (
		.din(new_net_2588),
		.dout(new_net_2587)
	);

	bfr new_net_2589_bfr_before (
		.din(new_net_2589),
		.dout(new_net_2588)
	);

	bfr new_net_2590_bfr_before (
		.din(new_net_2590),
		.dout(new_net_2589)
	);

	bfr new_net_2591_bfr_before (
		.din(new_net_2591),
		.dout(new_net_2590)
	);

	bfr new_net_2592_bfr_before (
		.din(new_net_2592),
		.dout(new_net_2591)
	);

	spl3L new_net_2094_v_fanout (
		.a(new_net_2094),
		.b(new_net_2592),
		.c(new_net_284),
		.d(new_net_285)
	);

	bfr new_net_2593_bfr_before (
		.din(new_net_2593),
		.dout(new_net_1505)
	);

	bfr new_net_2594_bfr_before (
		.din(new_net_2594),
		.dout(new_net_2593)
	);

	bfr new_net_2595_bfr_before (
		.din(new_net_2595),
		.dout(new_net_2594)
	);

	bfr new_net_2596_bfr_before (
		.din(new_net_2596),
		.dout(new_net_1506)
	);

	bfr new_net_2597_bfr_before (
		.din(new_net_2597),
		.dout(new_net_2596)
	);

	bfr new_net_2598_bfr_before (
		.din(new_net_2598),
		.dout(new_net_2597)
	);

	bfr new_net_2599_bfr_before (
		.din(new_net_2599),
		.dout(new_net_1504)
	);

	bfr new_net_2600_bfr_before (
		.din(new_net_2600),
		.dout(new_net_2599)
	);

	bfr new_net_2601_bfr_before (
		.din(new_net_2601),
		.dout(new_net_2600)
	);

	spl4L new_net_1899_v_fanout (
		.a(new_net_1899),
		.b(new_net_2598),
		.c(new_net_2601),
		.d(new_net_1900),
		.e(new_net_2595)
	);

	bfr new_net_2602_bfr_before (
		.din(new_net_2602),
		.dout(new_net_669)
	);

	spl2 new_net_1824_v_fanout (
		.a(new_net_1824),
		.b(new_net_658),
		.c(new_net_2602)
	);

	spl2 new_net_2093_v_fanout (
		.a(new_net_2093),
		.b(new_net_286),
		.c(new_net_283)
	);

	spl2 _0085__v_fanout (
		.a(_0085_),
		.b(new_net_1715),
		.c(new_net_1716)
	);

	bfr new_net_2603_bfr_before (
		.din(new_net_2603),
		.dout(new_net_380)
	);

	spl2 new_net_1981_v_fanout (
		.a(new_net_1981),
		.b(new_net_381),
		.c(new_net_2603)
	);

	bfr new_net_2604_bfr_before (
		.din(new_net_2604),
		.dout(new_net_928)
	);

	bfr new_net_2605_bfr_before (
		.din(new_net_2605),
		.dout(new_net_2604)
	);

	bfr new_net_2606_bfr_before (
		.din(new_net_2606),
		.dout(new_net_2605)
	);

	bfr new_net_2607_bfr_before (
		.din(new_net_2607),
		.dout(new_net_2606)
	);

	bfr new_net_2608_bfr_before (
		.din(new_net_2608),
		.dout(new_net_931)
	);

	bfr new_net_2609_bfr_before (
		.din(new_net_2609),
		.dout(new_net_948)
	);

	spl4L new_net_1800_v_fanout (
		.a(new_net_1800),
		.b(new_net_2607),
		.c(new_net_2608),
		.d(new_net_2609),
		.e(new_net_946)
	);

	spl2 new_net_23_v_fanout (
		.a(new_net_23),
		.b(new_net_2096),
		.c(new_net_2095)
	);

	bfr new_net_2610_bfr_before (
		.din(new_net_2610),
		.dout(new_net_153)
	);

	bfr new_net_2611_bfr_before (
		.din(new_net_2611),
		.dout(new_net_151)
	);

	bfr new_net_2612_bfr_before (
		.din(new_net_2612),
		.dout(new_net_2611)
	);

	bfr new_net_2613_bfr_before (
		.din(new_net_2613),
		.dout(new_net_2612)
	);

	spl3L new_net_1866_v_fanout (
		.a(new_net_1866),
		.b(new_net_2610),
		.c(new_net_2613),
		.d(new_net_148)
	);

	bfr new_net_2614_bfr_before (
		.din(new_net_2614),
		.dout(new_net_152)
	);

	bfr new_net_2615_bfr_before (
		.din(new_net_2615),
		.dout(new_net_2614)
	);

	spl2 new_net_1865_v_fanout (
		.a(new_net_1865),
		.b(new_net_155),
		.c(new_net_2615)
	);

	spl2 _1015__v_fanout (
		.a(_1015_),
		.b(new_net_1597),
		.c(new_net_1598)
	);

	spl2 _0994__v_fanout (
		.a(_0994_),
		.b(new_net_1161),
		.c(new_net_1162)
	);

	spl2 new_net_22_v_fanout (
		.a(new_net_22),
		.b(new_net_2094),
		.c(new_net_2093)
	);

	spl2 _1121__v_fanout (
		.a(_1121_),
		.b(new_net_806),
		.c(new_net_807)
	);

	bfr new_net_2616_bfr_before (
		.din(new_net_2616),
		.dout(new_net_1958)
	);

	spl2 new_net_1957_v_fanout (
		.a(new_net_1957),
		.b(new_net_1355),
		.c(new_net_2616)
	);

	spl2 _0975__v_fanout (
		.a(_0975_),
		.b(new_net_1719),
		.c(new_net_1720)
	);

	spl2 new_net_1964_v_fanout (
		.a(new_net_1964),
		.b(new_net_1965),
		.c(new_net_675)
	);

	bfr new_net_2617_bfr_before (
		.din(new_net_2617),
		.dout(new_net_1948)
	);

	bfr new_net_2618_bfr_before (
		.din(new_net_2618),
		.dout(new_net_2617)
	);

	spl2 new_net_1947_v_fanout (
		.a(new_net_1947),
		.b(new_net_1156),
		.c(new_net_2618)
	);

	bfr new_net_2619_bfr_before (
		.din(new_net_2619),
		.dout(new_net_1858)
	);

	bfr new_net_2620_bfr_before (
		.din(new_net_2620),
		.dout(new_net_2619)
	);

	bfr new_net_2621_bfr_before (
		.din(new_net_2621),
		.dout(new_net_2620)
	);

	spl3L new_net_1857_v_fanout (
		.a(new_net_1857),
		.b(new_net_2621),
		.c(new_net_117),
		.d(new_net_118)
	);

	bfr new_net_2622_bfr_before (
		.din(new_net_2622),
		.dout(new_net_1988)
	);

	bfr new_net_2623_bfr_before (
		.din(new_net_2623),
		.dout(new_net_2622)
	);

	spl2 new_net_1987_v_fanout (
		.a(new_net_1987),
		.b(new_net_1571),
		.c(new_net_2623)
	);

	spl2 new_net_1931_v_fanout (
		.a(new_net_1931),
		.b(new_net_440),
		.c(new_net_1932)
	);

	bfr new_net_2624_bfr_before (
		.din(new_net_2624),
		.dout(new_net_661)
	);

	bfr new_net_2625_bfr_before (
		.din(new_net_2625),
		.dout(new_net_2624)
	);

	bfr new_net_2626_bfr_before (
		.din(new_net_2626),
		.dout(new_net_2625)
	);

	bfr new_net_2627_bfr_before (
		.din(new_net_2627),
		.dout(new_net_670)
	);

	bfr new_net_2628_bfr_before (
		.din(new_net_2628),
		.dout(new_net_2627)
	);

	bfr new_net_2629_bfr_before (
		.din(new_net_2629),
		.dout(new_net_2628)
	);

	bfr new_net_2630_bfr_before (
		.din(new_net_2630),
		.dout(new_net_671)
	);

	bfr new_net_2631_bfr_before (
		.din(new_net_2631),
		.dout(new_net_2630)
	);

	bfr new_net_2632_bfr_before (
		.din(new_net_2632),
		.dout(new_net_2631)
	);

	spl4L new_net_1823_v_fanout (
		.a(new_net_1823),
		.b(new_net_2629),
		.c(new_net_2632),
		.d(new_net_1824),
		.e(new_net_2626)
	);

	spl2 new_net_1972_v_fanout (
		.a(new_net_1972),
		.b(new_net_798),
		.c(new_net_1973)
	);

	bfr new_net_2633_bfr_before (
		.din(new_net_2633),
		.dout(new_net_164)
	);

	spl2 _0895__v_fanout (
		.a(_0895_),
		.b(new_net_163),
		.c(new_net_2633)
	);

	bfr new_net_2634_bfr_before (
		.din(new_net_2634),
		.dout(new_net_941)
	);

	bfr new_net_2635_bfr_before (
		.din(new_net_2635),
		.dout(new_net_2634)
	);

	bfr new_net_2636_bfr_before (
		.din(new_net_2636),
		.dout(new_net_2635)
	);

	bfr new_net_2637_bfr_before (
		.din(new_net_2637),
		.dout(new_net_944)
	);

	bfr new_net_2638_bfr_before (
		.din(new_net_2638),
		.dout(new_net_2637)
	);

	bfr new_net_2639_bfr_before (
		.din(new_net_2639),
		.dout(new_net_2638)
	);

	bfr new_net_2640_bfr_before (
		.din(new_net_2640),
		.dout(new_net_943)
	);

	bfr new_net_2641_bfr_before (
		.din(new_net_2641),
		.dout(new_net_2640)
	);

	bfr new_net_2642_bfr_before (
		.din(new_net_2642),
		.dout(new_net_2641)
	);

	spl4L new_net_1799_v_fanout (
		.a(new_net_1799),
		.b(new_net_2639),
		.c(new_net_2642),
		.d(new_net_1800),
		.e(new_net_2636)
	);

	spl2 _0881__v_fanout (
		.a(_0881_),
		.b(new_net_401),
		.c(new_net_402)
	);

	spl3L new_net_1862_v_fanout (
		.a(new_net_1862),
		.b(new_net_114),
		.c(new_net_113),
		.d(new_net_109)
	);

	bfr new_net_2643_bfr_before (
		.din(new_net_2643),
		.dout(G5257)
	);

	bfr new_net_2644_bfr_before (
		.din(new_net_2644),
		.dout(new_net_2643)
	);

	bfr new_net_2645_bfr_before (
		.din(new_net_2645),
		.dout(new_net_2644)
	);

	bfr new_net_2646_bfr_before (
		.din(new_net_2646),
		.dout(new_net_2645)
	);

	bfr new_net_2647_bfr_before (
		.din(new_net_2647),
		.dout(new_net_2646)
	);

	bfr new_net_2648_bfr_before (
		.din(new_net_2648),
		.dout(new_net_2647)
	);

	bfr new_net_2649_bfr_before (
		.din(new_net_2649),
		.dout(new_net_2648)
	);

	bfr new_net_2650_bfr_before (
		.din(new_net_2650),
		.dout(new_net_2649)
	);

	bfr new_net_2651_bfr_before (
		.din(new_net_2651),
		.dout(new_net_2650)
	);

	bfr new_net_2652_bfr_before (
		.din(new_net_2652),
		.dout(new_net_2651)
	);

	bfr new_net_2653_bfr_before (
		.din(new_net_2653),
		.dout(new_net_2652)
	);

	bfr new_net_2654_bfr_before (
		.din(new_net_2654),
		.dout(new_net_2653)
	);

	bfr new_net_2655_bfr_before (
		.din(new_net_2655),
		.dout(new_net_2654)
	);

	bfr new_net_2656_bfr_before (
		.din(new_net_2656),
		.dout(new_net_2655)
	);

	spl3L new_net_2092_v_fanout (
		.a(new_net_2092),
		.b(new_net_2656),
		.c(new_net_321),
		.d(new_net_320)
	);

	bfr new_net_2657_bfr_before (
		.din(new_net_2657),
		.dout(new_net_154)
	);

	bfr new_net_2658_bfr_before (
		.din(new_net_2658),
		.dout(new_net_1866)
	);

	bfr new_net_2659_bfr_before (
		.din(new_net_2659),
		.dout(new_net_2658)
	);

	bfr new_net_2660_bfr_before (
		.din(new_net_2660),
		.dout(new_net_1865)
	);

	spl4L new_net_1864_v_fanout (
		.a(new_net_1864),
		.b(new_net_2657),
		.c(new_net_2659),
		.d(new_net_2660),
		.e(new_net_150)
	);

	spl2 new_net_2091_v_fanout (
		.a(new_net_2091),
		.b(new_net_323),
		.c(new_net_322)
	);

	spl2 new_net_1856_v_fanout (
		.a(new_net_1856),
		.b(new_net_1857),
		.c(new_net_108)
	);

	spl2 new_net_1798_v_fanout (
		.a(new_net_1798),
		.b(new_net_932),
		.c(new_net_1799)
	);

	bfr new_net_2661_bfr_before (
		.din(new_net_2661),
		.dout(new_net_1498)
	);

	spl2 new_net_1898_v_fanout (
		.a(new_net_1898),
		.b(new_net_2661),
		.c(new_net_1899)
	);

	spl2 _0991__v_fanout (
		.a(_0991_),
		.b(new_net_72),
		.c(new_net_73)
	);

	bfr new_net_2662_bfr_before (
		.din(new_net_2662),
		.dout(new_net_1972)
	);

	bfr new_net_2663_bfr_before (
		.din(new_net_2663),
		.dout(new_net_2662)
	);

	bfr new_net_2664_bfr_before (
		.din(new_net_2664),
		.dout(new_net_2663)
	);

	bfr new_net_2665_bfr_before (
		.din(new_net_2665),
		.dout(new_net_2664)
	);

	spl2 new_net_1971_v_fanout (
		.a(new_net_1971),
		.b(new_net_797),
		.c(new_net_2665)
	);

	bfr new_net_2666_bfr_before (
		.din(new_net_2666),
		.dout(G5258)
	);

	bfr new_net_2667_bfr_before (
		.din(new_net_2667),
		.dout(new_net_2666)
	);

	bfr new_net_2668_bfr_before (
		.din(new_net_2668),
		.dout(new_net_2667)
	);

	bfr new_net_2669_bfr_before (
		.din(new_net_2669),
		.dout(new_net_2668)
	);

	bfr new_net_2670_bfr_before (
		.din(new_net_2670),
		.dout(new_net_2669)
	);

	bfr new_net_2671_bfr_before (
		.din(new_net_2671),
		.dout(new_net_2670)
	);

	bfr new_net_2672_bfr_before (
		.din(new_net_2672),
		.dout(new_net_2671)
	);

	bfr new_net_2673_bfr_before (
		.din(new_net_2673),
		.dout(new_net_2672)
	);

	bfr new_net_2674_bfr_before (
		.din(new_net_2674),
		.dout(new_net_2673)
	);

	bfr new_net_2675_bfr_before (
		.din(new_net_2675),
		.dout(new_net_2674)
	);

	bfr new_net_2676_bfr_before (
		.din(new_net_2676),
		.dout(new_net_2675)
	);

	bfr new_net_2677_bfr_before (
		.din(new_net_2677),
		.dout(new_net_2676)
	);

	bfr new_net_2678_bfr_before (
		.din(new_net_2678),
		.dout(new_net_2677)
	);

	bfr new_net_2679_bfr_before (
		.din(new_net_2679),
		.dout(new_net_2678)
	);

	bfr new_net_2680_bfr_before (
		.din(new_net_2680),
		.dout(new_net_2679)
	);

	spl3L new_net_2086_v_fanout (
		.a(new_net_2086),
		.b(new_net_2680),
		.c(new_net_894),
		.d(new_net_897)
	);

	spl2 _1011__v_fanout (
		.a(_1011_),
		.b(new_net_1186),
		.c(new_net_1187)
	);

	spl2 _0972__v_fanout (
		.a(_0972_),
		.b(new_net_521),
		.c(new_net_522)
	);

	bfr new_net_2681_bfr_before (
		.din(new_net_2681),
		.dout(new_net_1931)
	);

	bfr new_net_2682_bfr_before (
		.din(new_net_2682),
		.dout(new_net_2681)
	);

	bfr new_net_2683_bfr_before (
		.din(new_net_2683),
		.dout(new_net_2682)
	);

	bfr new_net_2684_bfr_before (
		.din(new_net_2684),
		.dout(new_net_2683)
	);

	spl2 new_net_1930_v_fanout (
		.a(new_net_1930),
		.b(new_net_434),
		.c(new_net_2684)
	);

	bfr new_net_2685_bfr_before (
		.din(new_net_2685),
		.dout(G5253)
	);

	bfr new_net_2686_bfr_before (
		.din(new_net_2686),
		.dout(new_net_2685)
	);

	bfr new_net_2687_bfr_before (
		.din(new_net_2687),
		.dout(new_net_2686)
	);

	bfr new_net_2688_bfr_before (
		.din(new_net_2688),
		.dout(new_net_2687)
	);

	bfr new_net_2689_bfr_before (
		.din(new_net_2689),
		.dout(new_net_2688)
	);

	bfr new_net_2690_bfr_before (
		.din(new_net_2690),
		.dout(new_net_2689)
	);

	bfr new_net_2691_bfr_before (
		.din(new_net_2691),
		.dout(new_net_2690)
	);

	bfr new_net_2692_bfr_before (
		.din(new_net_2692),
		.dout(new_net_2691)
	);

	bfr new_net_2693_bfr_before (
		.din(new_net_2693),
		.dout(new_net_2692)
	);

	bfr new_net_2694_bfr_before (
		.din(new_net_2694),
		.dout(new_net_2693)
	);

	bfr new_net_2695_bfr_before (
		.din(new_net_2695),
		.dout(new_net_2694)
	);

	bfr new_net_2696_bfr_before (
		.din(new_net_2696),
		.dout(new_net_2695)
	);

	bfr new_net_2697_bfr_before (
		.din(new_net_2697),
		.dout(new_net_2696)
	);

	bfr new_net_2698_bfr_before (
		.din(new_net_2698),
		.dout(new_net_2697)
	);

	bfr new_net_2699_bfr_before (
		.din(new_net_2699),
		.dout(new_net_2698)
	);

	spl3L new_net_2090_v_fanout (
		.a(new_net_2090),
		.b(new_net_2699),
		.c(new_net_419),
		.d(new_net_418)
	);

	bfr new_net_2700_bfr_before (
		.din(new_net_2700),
		.dout(new_net_1957)
	);

	bfr new_net_2701_bfr_before (
		.din(new_net_2701),
		.dout(new_net_2700)
	);

	bfr new_net_2702_bfr_before (
		.din(new_net_2702),
		.dout(new_net_2701)
	);

	spl2 new_net_1956_v_fanout (
		.a(new_net_1956),
		.b(new_net_1348),
		.c(new_net_2702)
	);

	spl2 _1032__v_fanout (
		.a(_1032_),
		.b(new_net_82),
		.c(new_net_83)
	);

	bfr new_net_2703_bfr_after (
		.din(_1080_),
		.dout(new_net_2703)
	);

	bfr new_net_2704_bfr_after (
		.din(new_net_2703),
		.dout(new_net_2704)
	);

	bfr new_net_2705_bfr_after (
		.din(new_net_2704),
		.dout(new_net_2705)
	);

	spl2 _1080__v_fanout (
		.a(new_net_2705),
		.b(new_net_1683),
		.c(new_net_1684)
	);

	spl2 _1116__v_fanout (
		.a(_1116_),
		.b(new_net_833),
		.c(new_net_834)
	);

	spl2 new_net_2089_v_fanout (
		.a(new_net_2089),
		.b(new_net_416),
		.c(new_net_417)
	);

	spl2 new_net_5_v_fanout (
		.a(new_net_5),
		.b(new_net_2091),
		.c(new_net_2092)
	);

	spl2 new_net_2087_v_fanout (
		.a(new_net_2087),
		.b(new_net_30),
		.c(new_net_29)
	);

	bfr new_net_2706_bfr_before (
		.din(new_net_2706),
		.dout(new_net_1964)
	);

	bfr new_net_2707_bfr_before (
		.din(new_net_2707),
		.dout(new_net_2706)
	);

	bfr new_net_2708_bfr_before (
		.din(new_net_2708),
		.dout(new_net_2707)
	);

	spl2 new_net_1963_v_fanout (
		.a(new_net_1963),
		.b(new_net_674),
		.c(new_net_2708)
	);

	bfr new_net_2709_bfr_before (
		.din(new_net_2709),
		.dout(G5259)
	);

	bfr new_net_2710_bfr_before (
		.din(new_net_2710),
		.dout(new_net_2709)
	);

	bfr new_net_2711_bfr_before (
		.din(new_net_2711),
		.dout(new_net_2710)
	);

	bfr new_net_2712_bfr_before (
		.din(new_net_2712),
		.dout(new_net_2711)
	);

	bfr new_net_2713_bfr_before (
		.din(new_net_2713),
		.dout(new_net_2712)
	);

	bfr new_net_2714_bfr_before (
		.din(new_net_2714),
		.dout(new_net_2713)
	);

	bfr new_net_2715_bfr_before (
		.din(new_net_2715),
		.dout(new_net_2714)
	);

	bfr new_net_2716_bfr_before (
		.din(new_net_2716),
		.dout(new_net_2715)
	);

	bfr new_net_2717_bfr_before (
		.din(new_net_2717),
		.dout(new_net_2716)
	);

	bfr new_net_2718_bfr_before (
		.din(new_net_2718),
		.dout(new_net_2717)
	);

	bfr new_net_2719_bfr_before (
		.din(new_net_2719),
		.dout(new_net_2718)
	);

	bfr new_net_2720_bfr_before (
		.din(new_net_2720),
		.dout(new_net_2719)
	);

	bfr new_net_2721_bfr_before (
		.din(new_net_2721),
		.dout(new_net_2720)
	);

	bfr new_net_2722_bfr_before (
		.din(new_net_2722),
		.dout(new_net_2721)
	);

	bfr new_net_2723_bfr_before (
		.din(new_net_2723),
		.dout(new_net_2722)
	);

	spl3L new_net_2088_v_fanout (
		.a(new_net_2088),
		.b(new_net_31),
		.c(new_net_2723),
		.d(new_net_32)
	);

	spl2 new_net_2085_v_fanout (
		.a(new_net_2085),
		.b(new_net_895),
		.c(new_net_896)
	);

	bfr new_net_2724_bfr_before (
		.din(new_net_2724),
		.dout(new_net_1947)
	);

	bfr new_net_2725_bfr_before (
		.din(new_net_2725),
		.dout(new_net_2724)
	);

	bfr new_net_2726_bfr_before (
		.din(new_net_2726),
		.dout(new_net_2725)
	);

	spl2 new_net_1946_v_fanout (
		.a(new_net_1946),
		.b(new_net_1155),
		.c(new_net_2726)
	);

	bfr new_net_2727_bfr_before (
		.din(new_net_2727),
		.dout(new_net_668)
	);

	spl2 new_net_1822_v_fanout (
		.a(new_net_1822),
		.b(new_net_1823),
		.c(new_net_2727)
	);

	spl2 _0004__v_fanout (
		.a(_0004_),
		.b(new_net_497),
		.c(new_net_498)
	);

	spl2 _0914__v_fanout (
		.a(_0914_),
		.b(new_net_350),
		.c(new_net_351)
	);

	spl2 _0878__v_fanout (
		.a(_0878_),
		.b(new_net_144),
		.c(new_net_145)
	);

	bfr new_net_2728_bfr_before (
		.din(new_net_2728),
		.dout(new_net_945)
	);

	bfr new_net_2729_bfr_before (
		.din(new_net_2729),
		.dout(new_net_2728)
	);

	spl2 new_net_1797_v_fanout (
		.a(new_net_1797),
		.b(new_net_2729),
		.c(new_net_1798)
	);

	spl2 _0892__v_fanout (
		.a(_0892_),
		.b(new_net_1485),
		.c(new_net_1486)
	);

	spl2 new_net_6_v_fanout (
		.a(new_net_6),
		.b(new_net_2090),
		.c(new_net_2089)
	);

	spl2 new_net_9_v_fanout (
		.a(new_net_9),
		.b(new_net_2087),
		.c(new_net_2088)
	);

	bfr new_net_2730_bfr_before (
		.din(new_net_2730),
		.dout(new_net_1898)
	);

	bfr new_net_2731_bfr_before (
		.din(new_net_2731),
		.dout(new_net_2730)
	);

	spl2 new_net_1897_v_fanout (
		.a(new_net_1897),
		.b(new_net_1496),
		.c(new_net_2731)
	);

	spl2 new_net_7_v_fanout (
		.a(new_net_7),
		.b(new_net_2085),
		.c(new_net_2086)
	);

	bfr new_net_2732_bfr_before (
		.din(new_net_2732),
		.dout(new_net_1987)
	);

	bfr new_net_2733_bfr_before (
		.din(new_net_2733),
		.dout(new_net_2732)
	);

	bfr new_net_2734_bfr_before (
		.din(new_net_2734),
		.dout(new_net_2733)
	);

	spl2 new_net_1986_v_fanout (
		.a(new_net_1986),
		.b(new_net_2734),
		.c(new_net_1576)
	);

	bfr new_net_2735_bfr_before (
		.din(new_net_2735),
		.dout(new_net_376)
	);

	bfr new_net_2736_bfr_before (
		.din(new_net_2736),
		.dout(new_net_1981)
	);

	bfr new_net_2737_bfr_before (
		.din(new_net_2737),
		.dout(new_net_2736)
	);

	bfr new_net_2738_bfr_before (
		.din(new_net_2738),
		.dout(new_net_2737)
	);

	bfr new_net_2739_bfr_before (
		.din(new_net_2739),
		.dout(new_net_2738)
	);

	bfr new_net_2740_bfr_before (
		.din(new_net_2740),
		.dout(new_net_2739)
	);

	bfr new_net_2741_bfr_before (
		.din(new_net_2741),
		.dout(new_net_2740)
	);

	spl3L new_net_1980_v_fanout (
		.a(new_net_1980),
		.b(new_net_383),
		.c(new_net_2735),
		.d(new_net_2741)
	);

	bfr new_net_2742_bfr_before (
		.din(new_net_2742),
		.dout(new_net_1210)
	);

	spl3L new_net_1740_v_fanout (
		.a(new_net_1740),
		.b(new_net_1218),
		.c(new_net_1209),
		.d(new_net_2742)
	);

	bfr new_net_2743_bfr_before (
		.din(new_net_2743),
		.dout(new_net_1822)
	);

	bfr new_net_2744_bfr_before (
		.din(new_net_2744),
		.dout(new_net_2743)
	);

	spl2 new_net_1821_v_fanout (
		.a(new_net_1821),
		.b(new_net_2744),
		.c(new_net_659)
	);

	spl2 new_net_2083_v_fanout (
		.a(new_net_2083),
		.b(new_net_1086),
		.c(new_net_1083)
	);

	spl3L new_net_1896_v_fanout (
		.a(new_net_1896),
		.b(new_net_1503),
		.c(new_net_1497),
		.d(new_net_1897)
	);

	spl2 new_net_2011_v_fanout (
		.a(new_net_2011),
		.b(new_net_306),
		.c(new_net_310)
	);

	bfr new_net_2745_bfr_before (
		.din(new_net_2745),
		.dout(new_net_378)
	);

	bfr new_net_2746_bfr_before (
		.din(new_net_2746),
		.dout(new_net_377)
	);

	spl3L new_net_1979_v_fanout (
		.a(new_net_1979),
		.b(new_net_2745),
		.c(new_net_2746),
		.d(new_net_1980)
	);

	bfr new_net_2747_bfr_before (
		.din(new_net_2747),
		.dout(new_net_1956)
	);

	spl2 new_net_1955_v_fanout (
		.a(new_net_1955),
		.b(new_net_1349),
		.c(new_net_2747)
	);

	bfr new_net_2748_bfr_before (
		.din(new_net_2748),
		.dout(G5254)
	);

	bfr new_net_2749_bfr_before (
		.din(new_net_2749),
		.dout(new_net_2748)
	);

	bfr new_net_2750_bfr_before (
		.din(new_net_2750),
		.dout(new_net_2749)
	);

	bfr new_net_2751_bfr_before (
		.din(new_net_2751),
		.dout(new_net_2750)
	);

	bfr new_net_2752_bfr_before (
		.din(new_net_2752),
		.dout(new_net_2751)
	);

	bfr new_net_2753_bfr_before (
		.din(new_net_2753),
		.dout(new_net_2752)
	);

	bfr new_net_2754_bfr_before (
		.din(new_net_2754),
		.dout(new_net_2753)
	);

	bfr new_net_2755_bfr_before (
		.din(new_net_2755),
		.dout(new_net_2754)
	);

	bfr new_net_2756_bfr_before (
		.din(new_net_2756),
		.dout(new_net_2755)
	);

	bfr new_net_2757_bfr_before (
		.din(new_net_2757),
		.dout(new_net_2756)
	);

	bfr new_net_2758_bfr_before (
		.din(new_net_2758),
		.dout(new_net_2757)
	);

	bfr new_net_2759_bfr_before (
		.din(new_net_2759),
		.dout(new_net_2758)
	);

	bfr new_net_2760_bfr_before (
		.din(new_net_2760),
		.dout(new_net_2759)
	);

	bfr new_net_2761_bfr_before (
		.din(new_net_2761),
		.dout(new_net_2760)
	);

	bfr new_net_2762_bfr_before (
		.din(new_net_2762),
		.dout(new_net_2761)
	);

	bfr new_net_2763_bfr_before (
		.din(new_net_2763),
		.dout(new_net_2762)
	);

	bfr new_net_2764_bfr_before (
		.din(new_net_2764),
		.dout(new_net_2763)
	);

	spl3L new_net_2084_v_fanout (
		.a(new_net_2084),
		.b(new_net_1082),
		.c(new_net_1085),
		.d(new_net_2764)
	);

	bfr new_net_2765_bfr_before (
		.din(new_net_2765),
		.dout(new_net_1862)
	);

	bfr new_net_2766_bfr_before (
		.din(new_net_2766),
		.dout(new_net_2765)
	);

	bfr new_net_2767_bfr_before (
		.din(new_net_2767),
		.dout(new_net_2766)
	);

	bfr new_net_2768_bfr_before (
		.din(new_net_2768),
		.dout(new_net_1856)
	);

	bfr new_net_2769_bfr_before (
		.din(new_net_2769),
		.dout(new_net_2768)
	);

	bfr new_net_2770_bfr_before (
		.din(new_net_2770),
		.dout(new_net_2769)
	);

	spl4L new_net_1855_v_fanout (
		.a(new_net_1855),
		.b(new_net_125),
		.c(new_net_126),
		.d(new_net_2770),
		.e(new_net_2767)
	);

	bfr new_net_2771_bfr_before (
		.din(new_net_2771),
		.dout(new_net_938)
	);

	bfr new_net_2772_bfr_before (
		.din(new_net_2772),
		.dout(new_net_1797)
	);

	bfr new_net_2773_bfr_before (
		.din(new_net_2773),
		.dout(new_net_2772)
	);

	spl3L new_net_1796_v_fanout (
		.a(new_net_1796),
		.b(new_net_2771),
		.c(new_net_933),
		.d(new_net_2773)
	);

	bfr new_net_2774_bfr_before (
		.din(new_net_2774),
		.dout(new_net_1963)
	);

	spl2 new_net_1962_v_fanout (
		.a(new_net_1962),
		.b(new_net_679),
		.c(new_net_2774)
	);

	spl2 new_net_2041_v_fanout (
		.a(new_net_2041),
		.b(new_net_390),
		.c(new_net_392)
	);

	bfr new_net_2775_bfr_before (
		.din(new_net_2775),
		.dout(new_net_1971)
	);

	spl2 new_net_1970_v_fanout (
		.a(new_net_1970),
		.b(new_net_803),
		.c(new_net_2775)
	);

	bfr new_net_2776_bfr_before (
		.din(new_net_2776),
		.dout(new_net_1930)
	);

	spl2 new_net_1929_v_fanout (
		.a(new_net_1929),
		.b(new_net_433),
		.c(new_net_2776)
	);

	bfr new_net_2777_bfr_before (
		.din(new_net_2777),
		.dout(new_net_1212)
	);

	spl2 new_net_1739_v_fanout (
		.a(new_net_1739),
		.b(new_net_1222),
		.c(new_net_2777)
	);

	spl2 new_net_2054_v_fanout (
		.a(new_net_2054),
		.b(new_net_1444),
		.c(new_net_1446)
	);

	spl2 new_net_2052_v_fanout (
		.a(new_net_2052),
		.b(new_net_207),
		.c(new_net_206)
	);

	bfr new_net_2778_bfr_before (
		.din(new_net_2778),
		.dout(new_net_1986)
	);

	spl2 new_net_1985_v_fanout (
		.a(new_net_1985),
		.b(new_net_1570),
		.c(new_net_2778)
	);

	bfr new_net_2779_bfr_before (
		.din(new_net_2779),
		.dout(new_net_939)
	);

	spl2 new_net_1795_v_fanout (
		.a(new_net_1795),
		.b(new_net_2779),
		.c(new_net_1796)
	);

	spl2 new_net_1978_v_fanout (
		.a(new_net_1978),
		.b(new_net_385),
		.c(new_net_1979)
	);

	spl2 new_net_8_v_fanout (
		.a(new_net_8),
		.b(new_net_2084),
		.c(new_net_2083)
	);

	spl4L new_net_2082_v_fanout (
		.a(new_net_2082),
		.b(new_net_356),
		.c(new_net_358),
		.d(new_net_359),
		.e(new_net_357)
	);

	bfr new_net_2780_bfr_before (
		.din(new_net_2780),
		.dout(new_net_1946)
	);

	spl2 new_net_1945_v_fanout (
		.a(new_net_1945),
		.b(new_net_1150),
		.c(new_net_2780)
	);

	spl2 new_net_2081_v_fanout (
		.a(new_net_2081),
		.b(new_net_360),
		.c(new_net_361)
	);

	spl2 new_net_1820_v_fanout (
		.a(new_net_1820),
		.b(new_net_1821),
		.c(new_net_660)
	);

	bfr new_net_2781_bfr_after (
		.din(_0024_),
		.dout(new_net_2781)
	);

	bfr new_net_2782_bfr_after (
		.din(new_net_2781),
		.dout(new_net_2782)
	);

	bfr new_net_2783_bfr_after (
		.din(new_net_2782),
		.dout(new_net_2783)
	);

	spl2 _0024__v_fanout (
		.a(new_net_2783),
		.b(new_net_1324),
		.c(new_net_1325)
	);

	spl2 new_net_2079_v_fanout (
		.a(new_net_2079),
		.b(new_net_1125),
		.c(new_net_1123)
	);

	spl4L new_net_2076_v_fanout (
		.a(new_net_2076),
		.b(new_net_1615),
		.c(new_net_1614),
		.d(new_net_1617),
		.e(new_net_1613)
	);

	spl3L new_net_2075_v_fanout (
		.a(new_net_2075),
		.b(new_net_1616),
		.c(new_net_1618),
		.d(new_net_1619)
	);

	bfr new_net_2784_bfr_before (
		.din(new_net_2784),
		.dout(new_net_942)
	);

	bfr new_net_2785_bfr_before (
		.din(new_net_2785),
		.dout(new_net_2784)
	);

	spl3L new_net_1794_v_fanout (
		.a(new_net_1794),
		.b(new_net_930),
		.c(new_net_2785),
		.d(new_net_1795)
	);

	bfr new_net_2786_bfr_before (
		.din(new_net_2786),
		.dout(new_net_1740)
	);

	bfr new_net_2787_bfr_before (
		.din(new_net_2787),
		.dout(new_net_1739)
	);

	bfr new_net_2788_bfr_before (
		.din(new_net_2788),
		.dout(new_net_2787)
	);

	spl3L new_net_1738_v_fanout (
		.a(new_net_1738),
		.b(new_net_1219),
		.c(new_net_2786),
		.d(new_net_2788)
	);

	bfr new_net_2789_bfr_before (
		.din(new_net_2789),
		.dout(new_net_1962)
	);

	spl2 new_net_1961_v_fanout (
		.a(new_net_1961),
		.b(new_net_673),
		.c(new_net_2789)
	);

	bfr new_net_2790_bfr_before (
		.din(new_net_2790),
		.dout(G5260)
	);

	bfr new_net_2791_bfr_before (
		.din(new_net_2791),
		.dout(new_net_2790)
	);

	bfr new_net_2792_bfr_before (
		.din(new_net_2792),
		.dout(new_net_2791)
	);

	bfr new_net_2793_bfr_before (
		.din(new_net_2793),
		.dout(new_net_2792)
	);

	bfr new_net_2794_bfr_before (
		.din(new_net_2794),
		.dout(new_net_2793)
	);

	bfr new_net_2795_bfr_before (
		.din(new_net_2795),
		.dout(new_net_2794)
	);

	bfr new_net_2796_bfr_before (
		.din(new_net_2796),
		.dout(new_net_2795)
	);

	bfr new_net_2797_bfr_before (
		.din(new_net_2797),
		.dout(new_net_2796)
	);

	bfr new_net_2798_bfr_before (
		.din(new_net_2798),
		.dout(new_net_2797)
	);

	bfr new_net_2799_bfr_before (
		.din(new_net_2799),
		.dout(new_net_2798)
	);

	bfr new_net_2800_bfr_before (
		.din(new_net_2800),
		.dout(new_net_2799)
	);

	bfr new_net_2801_bfr_before (
		.din(new_net_2801),
		.dout(new_net_2800)
	);

	bfr new_net_2802_bfr_before (
		.din(new_net_2802),
		.dout(new_net_2801)
	);

	bfr new_net_2803_bfr_before (
		.din(new_net_2803),
		.dout(new_net_2802)
	);

	bfr new_net_2804_bfr_before (
		.din(new_net_2804),
		.dout(new_net_2803)
	);

	bfr new_net_2805_bfr_before (
		.din(new_net_2805),
		.dout(new_net_2804)
	);

	bfr new_net_2806_bfr_before (
		.din(new_net_2806),
		.dout(new_net_2805)
	);

	bfr new_net_2807_bfr_before (
		.din(new_net_2807),
		.dout(new_net_2806)
	);

	bfr new_net_2808_bfr_before (
		.din(new_net_2808),
		.dout(new_net_2807)
	);

	spl3L new_net_2080_v_fanout (
		.a(new_net_2080),
		.b(new_net_2808),
		.c(new_net_1126),
		.d(new_net_1124)
	);

	bfr new_net_2809_bfr_before (
		.din(new_net_2809),
		.dout(new_net_774)
	);

	spl2 _0776__v_fanout (
		.a(_0776_),
		.b(new_net_773),
		.c(new_net_2809)
	);

	spl2 _0963__v_fanout (
		.a(_0963_),
		.b(new_net_2082),
		.c(new_net_2081)
	);

	spl2 _1095__v_fanout (
		.a(_1095_),
		.b(new_net_1423),
		.c(new_net_1424)
	);

	bfr new_net_2810_bfr_before (
		.din(new_net_2810),
		.dout(G5255)
	);

	bfr new_net_2811_bfr_before (
		.din(new_net_2811),
		.dout(new_net_2810)
	);

	bfr new_net_2812_bfr_before (
		.din(new_net_2812),
		.dout(new_net_2811)
	);

	bfr new_net_2813_bfr_before (
		.din(new_net_2813),
		.dout(new_net_2812)
	);

	bfr new_net_2814_bfr_before (
		.din(new_net_2814),
		.dout(new_net_2813)
	);

	bfr new_net_2815_bfr_before (
		.din(new_net_2815),
		.dout(new_net_2814)
	);

	bfr new_net_2816_bfr_before (
		.din(new_net_2816),
		.dout(new_net_2815)
	);

	bfr new_net_2817_bfr_before (
		.din(new_net_2817),
		.dout(new_net_2816)
	);

	bfr new_net_2818_bfr_before (
		.din(new_net_2818),
		.dout(new_net_2817)
	);

	bfr new_net_2819_bfr_before (
		.din(new_net_2819),
		.dout(new_net_2818)
	);

	bfr new_net_2820_bfr_before (
		.din(new_net_2820),
		.dout(new_net_2819)
	);

	bfr new_net_2821_bfr_before (
		.din(new_net_2821),
		.dout(new_net_2820)
	);

	bfr new_net_2822_bfr_before (
		.din(new_net_2822),
		.dout(new_net_2821)
	);

	bfr new_net_2823_bfr_before (
		.din(new_net_2823),
		.dout(new_net_2822)
	);

	bfr new_net_2824_bfr_before (
		.din(new_net_2824),
		.dout(new_net_2823)
	);

	bfr new_net_2825_bfr_before (
		.din(new_net_2825),
		.dout(new_net_2824)
	);

	bfr new_net_2826_bfr_before (
		.din(new_net_2826),
		.dout(new_net_2825)
	);

	bfr new_net_2827_bfr_before (
		.din(new_net_2827),
		.dout(new_net_2826)
	);

	bfr new_net_2828_bfr_before (
		.din(new_net_2828),
		.dout(new_net_2827)
	);

	spl3L new_net_2078_v_fanout (
		.a(new_net_2078),
		.b(new_net_184),
		.c(new_net_185),
		.d(new_net_2828)
	);

	bfr new_net_2829_bfr_before (
		.din(new_net_2829),
		.dout(new_net_1955)
	);

	spl2 new_net_1954_v_fanout (
		.a(new_net_1954),
		.b(new_net_1351),
		.c(new_net_2829)
	);

	bfr new_net_2830_bfr_before (
		.din(new_net_2830),
		.dout(new_net_667)
	);

	spl2 new_net_1819_v_fanout (
		.a(new_net_1819),
		.b(new_net_2830),
		.c(new_net_1820)
	);

	bfr new_net_2831_bfr_before (
		.din(new_net_2831),
		.dout(new_net_1970)
	);

	spl2 new_net_1969_v_fanout (
		.a(new_net_1969),
		.b(new_net_796),
		.c(new_net_2831)
	);

	bfr new_net_2832_bfr_before (
		.din(new_net_2832),
		.dout(new_net_1929)
	);

	spl2 new_net_1928_v_fanout (
		.a(new_net_1928),
		.b(new_net_436),
		.c(new_net_2832)
	);

	spl2 new_net_2077_v_fanout (
		.a(new_net_2077),
		.b(new_net_186),
		.c(new_net_183)
	);

	spl2 _1057__v_fanout (
		.a(_1057_),
		.b(new_net_1381),
		.c(new_net_1382)
	);

	spl2 _1074__v_fanout (
		.a(_1074_),
		.b(new_net_997),
		.c(new_net_998)
	);

	bfr new_net_2833_bfr_before (
		.din(new_net_2833),
		.dout(new_net_1704)
	);

	spl2 _0819__v_fanout (
		.a(_0819_),
		.b(new_net_1703),
		.c(new_net_2833)
	);

	bfr new_net_2834_bfr_before (
		.din(new_net_2834),
		.dout(new_net_1985)
	);

	spl2 new_net_1984_v_fanout (
		.a(new_net_1984),
		.b(new_net_1575),
		.c(new_net_2834)
	);

	spl2 _1108__v_fanout (
		.a(_1108_),
		.b(new_net_690),
		.c(new_net_691)
	);

	spl2 _0798__v_fanout (
		.a(_0798_),
		.b(new_net_1280),
		.c(new_net_1281)
	);

	spl2 _0687__v_fanout (
		.a(_0687_),
		.b(new_net_562),
		.c(new_net_563)
	);

	spl2 new_net_11_v_fanout (
		.a(new_net_11),
		.b(new_net_2079),
		.c(new_net_2080)
	);

	spl2 _0876__v_fanout (
		.a(_0876_),
		.b(new_net_2075),
		.c(new_net_2076)
	);

	bfr new_net_2835_bfr_before (
		.din(new_net_2835),
		.dout(new_net_1945)
	);

	spl2 new_net_1944_v_fanout (
		.a(new_net_1944),
		.b(new_net_1154),
		.c(new_net_2835)
	);

	spl2 new_net_2047_v_fanout (
		.a(new_net_2047),
		.b(new_net_474),
		.c(new_net_473)
	);

	bfr new_net_2836_bfr_before (
		.din(new_net_2836),
		.dout(new_net_1978)
	);

	spl3L new_net_1977_v_fanout (
		.a(new_net_1977),
		.b(new_net_386),
		.c(new_net_379),
		.d(new_net_2836)
	);

	bfr new_net_2837_bfr_before (
		.din(new_net_2837),
		.dout(new_net_1224)
	);

	spl3L new_net_1737_v_fanout (
		.a(new_net_1737),
		.b(new_net_2837),
		.c(new_net_1228),
		.d(new_net_1738)
	);

	bfr new_net_2838_bfr_before (
		.din(new_net_2838),
		.dout(new_net_1896)
	);

	bfr new_net_2839_bfr_before (
		.din(new_net_2839),
		.dout(new_net_2838)
	);

	bfr new_net_2840_bfr_before (
		.din(new_net_2840),
		.dout(new_net_2839)
	);

	spl2 new_net_1895_v_fanout (
		.a(new_net_1895),
		.b(new_net_1502),
		.c(new_net_2840)
	);

	spl2 new_net_10_v_fanout (
		.a(new_net_10),
		.b(new_net_2078),
		.c(new_net_2077)
	);

	spl2 new_net_2049_v_fanout (
		.a(new_net_2049),
		.b(new_net_229),
		.c(new_net_231)
	);

	spl2 new_net_2074_v_fanout (
		.a(new_net_2074),
		.b(new_net_707),
		.c(new_net_706)
	);

	spl2 _0764__v_fanout (
		.a(_0764_),
		.b(new_net_867),
		.c(new_net_868)
	);

	bfr new_net_2841_bfr_before (
		.din(new_net_2841),
		.dout(new_net_1794)
	);

	spl3L new_net_1793_v_fanout (
		.a(new_net_1793),
		.b(new_net_940),
		.c(new_net_934),
		.d(new_net_2841)
	);

	bfr new_net_2842_bfr_before (
		.din(new_net_2842),
		.dout(new_net_1855)
	);

	bfr new_net_2843_bfr_before (
		.din(new_net_2843),
		.dout(new_net_2842)
	);

	bfr new_net_2844_bfr_before (
		.din(new_net_2844),
		.dout(new_net_2843)
	);

	spl3L new_net_1854_v_fanout (
		.a(new_net_1854),
		.b(new_net_112),
		.c(new_net_2844),
		.d(new_net_107)
	);

	bfr new_net_2845_bfr_before (
		.din(new_net_2845),
		.dout(new_net_1819)
	);

	bfr new_net_2846_bfr_before (
		.din(new_net_2846),
		.dout(new_net_2845)
	);

	spl2 new_net_1818_v_fanout (
		.a(new_net_1818),
		.b(new_net_2846),
		.c(new_net_666)
	);

	bfr new_net_2847_bfr_before (
		.din(new_net_2847),
		.dout(new_net_1928)
	);

	bfr new_net_2848_bfr_before (
		.din(new_net_2848),
		.dout(new_net_2847)
	);

	spl2 new_net_1927_v_fanout (
		.a(new_net_1927),
		.b(new_net_435),
		.c(new_net_2848)
	);

	bfr new_net_2849_bfr_before (
		.din(new_net_2849),
		.dout(new_net_1969)
	);

	bfr new_net_2850_bfr_before (
		.din(new_net_2850),
		.dout(new_net_2849)
	);

	spl2 new_net_1968_v_fanout (
		.a(new_net_1968),
		.b(new_net_802),
		.c(new_net_2850)
	);

	spl2 new_net_2072_v_fanout (
		.a(new_net_2072),
		.b(new_net_824),
		.c(new_net_823)
	);

	bfr new_net_2851_bfr_before (
		.din(new_net_2851),
		.dout(new_net_2074)
	);

	spl2 _0774__v_fanout (
		.a(_0774_),
		.b(new_net_705),
		.c(new_net_2851)
	);

	spl2 _1092__v_fanout (
		.a(_1092_),
		.b(new_net_446),
		.c(new_net_447)
	);

	spl2 _0706__v_fanout (
		.a(_0706_),
		.b(new_net_234),
		.c(new_net_235)
	);

	bfr new_net_2852_bfr_before (
		.din(new_net_2852),
		.dout(new_net_408)
	);

	bfr new_net_2853_bfr_before (
		.din(new_net_2853),
		.dout(new_net_2852)
	);

	spl2 new_net_2067_v_fanout (
		.a(new_net_2067),
		.b(new_net_2853),
		.c(new_net_409)
	);

	bfr new_net_2854_bfr_after (
		.din(_1067_),
		.dout(new_net_2854)
	);

	bfr new_net_2855_bfr_after (
		.din(new_net_2854),
		.dout(new_net_2855)
	);

	spl2 _1067__v_fanout (
		.a(new_net_2855),
		.b(new_net_1589),
		.c(new_net_1590)
	);

	bfr new_net_2856_bfr_before (
		.din(new_net_2856),
		.dout(new_net_1961)
	);

	bfr new_net_2857_bfr_before (
		.din(new_net_2857),
		.dout(new_net_2856)
	);

	spl2 new_net_1960_v_fanout (
		.a(new_net_1960),
		.b(new_net_678),
		.c(new_net_2857)
	);

	spl2 _0021__v_fanout (
		.a(_0021_),
		.b(new_net_788),
		.c(new_net_789)
	);

	spl2 _0007__v_fanout (
		.a(_0007_),
		.b(new_net_534),
		.c(new_net_535)
	);

	bfr new_net_2858_bfr_before (
		.din(new_net_2858),
		.dout(new_net_1737)
	);

	bfr new_net_2859_bfr_before (
		.din(new_net_2859),
		.dout(new_net_2858)
	);

	spl2 new_net_1736_v_fanout (
		.a(new_net_1736),
		.b(new_net_1225),
		.c(new_net_2859)
	);

	bfr new_net_2860_bfr_before (
		.din(new_net_2860),
		.dout(new_net_1954)
	);

	bfr new_net_2861_bfr_before (
		.din(new_net_2861),
		.dout(new_net_2860)
	);

	spl2 new_net_1953_v_fanout (
		.a(new_net_1953),
		.b(new_net_1350),
		.c(new_net_2861)
	);

	bfr new_net_2862_bfr_before (
		.din(new_net_2862),
		.dout(G5249)
	);

	bfr new_net_2863_bfr_before (
		.din(new_net_2863),
		.dout(new_net_2862)
	);

	bfr new_net_2864_bfr_before (
		.din(new_net_2864),
		.dout(new_net_2863)
	);

	bfr new_net_2865_bfr_before (
		.din(new_net_2865),
		.dout(new_net_2864)
	);

	bfr new_net_2866_bfr_before (
		.din(new_net_2866),
		.dout(new_net_2865)
	);

	bfr new_net_2867_bfr_before (
		.din(new_net_2867),
		.dout(new_net_2866)
	);

	bfr new_net_2868_bfr_before (
		.din(new_net_2868),
		.dout(new_net_2867)
	);

	bfr new_net_2869_bfr_before (
		.din(new_net_2869),
		.dout(new_net_2868)
	);

	bfr new_net_2870_bfr_before (
		.din(new_net_2870),
		.dout(new_net_2869)
	);

	bfr new_net_2871_bfr_before (
		.din(new_net_2871),
		.dout(new_net_2870)
	);

	bfr new_net_2872_bfr_before (
		.din(new_net_2872),
		.dout(new_net_2871)
	);

	bfr new_net_2873_bfr_before (
		.din(new_net_2873),
		.dout(new_net_2872)
	);

	bfr new_net_2874_bfr_before (
		.din(new_net_2874),
		.dout(new_net_2873)
	);

	bfr new_net_2875_bfr_before (
		.din(new_net_2875),
		.dout(new_net_2874)
	);

	bfr new_net_2876_bfr_before (
		.din(new_net_2876),
		.dout(new_net_2875)
	);

	bfr new_net_2877_bfr_before (
		.din(new_net_2877),
		.dout(new_net_2876)
	);

	bfr new_net_2878_bfr_before (
		.din(new_net_2878),
		.dout(new_net_2877)
	);

	bfr new_net_2879_bfr_before (
		.din(new_net_2879),
		.dout(new_net_2878)
	);

	bfr new_net_2880_bfr_before (
		.din(new_net_2880),
		.dout(new_net_2879)
	);

	bfr new_net_2881_bfr_before (
		.din(new_net_2881),
		.dout(new_net_2880)
	);

	bfr new_net_2882_bfr_before (
		.din(new_net_2882),
		.dout(new_net_2881)
	);

	bfr new_net_2883_bfr_before (
		.din(new_net_2883),
		.dout(new_net_2882)
	);

	spl3L new_net_2073_v_fanout (
		.a(new_net_2073),
		.b(new_net_820),
		.c(new_net_2883),
		.d(new_net_821)
	);

	bfr new_net_2884_bfr_before (
		.din(new_net_2884),
		.dout(new_net_1984)
	);

	bfr new_net_2885_bfr_before (
		.din(new_net_2885),
		.dout(new_net_2884)
	);

	spl2 new_net_1983_v_fanout (
		.a(new_net_1983),
		.b(new_net_1568),
		.c(new_net_2885)
	);

	spl2 _1070__v_fanout (
		.a(_1070_),
		.b(new_net_487),
		.c(new_net_488)
	);

	spl4L new_net_1735_v_fanout (
		.a(new_net_1735),
		.b(new_net_1206),
		.c(new_net_1220),
		.d(new_net_1205),
		.e(new_net_1736)
	);

	spl2 new_net_2042_v_fanout (
		.a(new_net_2042),
		.b(new_net_543),
		.c(new_net_541)
	);

	spl2 new_net_2068_v_fanout (
		.a(new_net_2068),
		.b(new_net_533),
		.c(new_net_531)
	);

	spl2 _0816__v_fanout (
		.a(_0816_),
		.b(new_net_1258),
		.c(new_net_1259)
	);

	spl3L _0678__v_fanout (
		.a(_0678_),
		.b(new_net_1360),
		.c(new_net_1362),
		.d(new_net_1361)
	);

	spl2 new_net_2046_v_fanout (
		.a(new_net_2046),
		.b(new_net_1648),
		.c(new_net_1650)
	);

	spl2 _0247__v_fanout (
		.a(_0247_),
		.b(new_net_317),
		.c(new_net_318)
	);

	bfr new_net_2886_bfr_before (
		.din(new_net_2886),
		.dout(new_net_1944)
	);

	bfr new_net_2887_bfr_before (
		.din(new_net_2887),
		.dout(new_net_2886)
	);

	spl2 new_net_1943_v_fanout (
		.a(new_net_1943),
		.b(new_net_1149),
		.c(new_net_2887)
	);

	bfr new_net_2888_bfr_before (
		.din(new_net_2888),
		.dout(new_net_1977)
	);

	bfr new_net_2889_bfr_before (
		.din(new_net_2889),
		.dout(new_net_2888)
	);

	spl2 new_net_1976_v_fanout (
		.a(new_net_1976),
		.b(new_net_387),
		.c(new_net_2889)
	);

	bfr new_net_2890_bfr_after (
		.din(new_net_16),
		.dout(new_net_2890)
	);

	bfr new_net_2891_bfr_before (
		.din(new_net_2891),
		.dout(G5262)
	);

	bfr new_net_2892_bfr_before (
		.din(new_net_2892),
		.dout(new_net_2891)
	);

	bfr new_net_2893_bfr_before (
		.din(new_net_2893),
		.dout(new_net_2892)
	);

	bfr new_net_2894_bfr_before (
		.din(new_net_2894),
		.dout(new_net_2893)
	);

	bfr new_net_2895_bfr_before (
		.din(new_net_2895),
		.dout(new_net_2894)
	);

	bfr new_net_2896_bfr_before (
		.din(new_net_2896),
		.dout(new_net_2895)
	);

	bfr new_net_2897_bfr_before (
		.din(new_net_2897),
		.dout(new_net_2896)
	);

	bfr new_net_2898_bfr_before (
		.din(new_net_2898),
		.dout(new_net_2897)
	);

	bfr new_net_2899_bfr_before (
		.din(new_net_2899),
		.dout(new_net_2898)
	);

	bfr new_net_2900_bfr_before (
		.din(new_net_2900),
		.dout(new_net_2899)
	);

	bfr new_net_2901_bfr_before (
		.din(new_net_2901),
		.dout(new_net_2900)
	);

	bfr new_net_2902_bfr_before (
		.din(new_net_2902),
		.dout(new_net_2901)
	);

	bfr new_net_2903_bfr_before (
		.din(new_net_2903),
		.dout(new_net_2902)
	);

	bfr new_net_2904_bfr_before (
		.din(new_net_2904),
		.dout(new_net_2903)
	);

	bfr new_net_2905_bfr_before (
		.din(new_net_2905),
		.dout(new_net_2904)
	);

	bfr new_net_2906_bfr_before (
		.din(new_net_2906),
		.dout(new_net_2905)
	);

	bfr new_net_2907_bfr_before (
		.din(new_net_2907),
		.dout(new_net_2906)
	);

	bfr new_net_2908_bfr_before (
		.din(new_net_2908),
		.dout(new_net_2907)
	);

	bfr new_net_2909_bfr_before (
		.din(new_net_2909),
		.dout(new_net_2908)
	);

	bfr new_net_2910_bfr_before (
		.din(new_net_2910),
		.dout(new_net_2909)
	);

	bfr new_net_2911_bfr_before (
		.din(new_net_2911),
		.dout(new_net_2910)
	);

	bfr new_net_2912_bfr_before (
		.din(new_net_2912),
		.dout(new_net_2911)
	);

	spl2 new_net_16_v_fanout (
		.a(new_net_2890),
		.b(new_net_2912),
		.c(new_net_1334)
	);

	spl2 new_net_2070_v_fanout (
		.a(new_net_2070),
		.b(new_net_422),
		.c(new_net_424)
	);

	spl2 new_net_12_v_fanout (
		.a(new_net_12),
		.b(new_net_2073),
		.c(new_net_2072)
	);

	spl2 _0795__v_fanout (
		.a(_0795_),
		.b(new_net_792),
		.c(new_net_793)
	);

	bfr new_net_2913_bfr_before (
		.din(new_net_2913),
		.dout(new_net_530)
	);

	bfr new_net_2914_bfr_before (
		.din(new_net_2914),
		.dout(new_net_2913)
	);

	bfr new_net_2915_bfr_before (
		.din(new_net_2915),
		.dout(new_net_2914)
	);

	spl3L new_net_2069_v_fanout (
		.a(new_net_2069),
		.b(new_net_529),
		.c(new_net_2915),
		.d(new_net_532)
	);

	bfr new_net_2916_bfr_before (
		.din(new_net_2916),
		.dout(new_net_2067)
	);

	spl2 new_net_2066_v_fanout (
		.a(new_net_2066),
		.b(new_net_2916),
		.c(new_net_410)
	);

	spl2 _1071__v_fanout (
		.a(_1071_),
		.b(new_net_1701),
		.c(new_net_1702)
	);

	spl2 new_net_2059_v_fanout (
		.a(new_net_2059),
		.b(new_net_635),
		.c(new_net_632)
	);

	bfr new_net_2917_bfr_before (
		.din(new_net_2917),
		.dout(G5250)
	);

	bfr new_net_2918_bfr_before (
		.din(new_net_2918),
		.dout(new_net_2917)
	);

	bfr new_net_2919_bfr_before (
		.din(new_net_2919),
		.dout(new_net_2918)
	);

	bfr new_net_2920_bfr_before (
		.din(new_net_2920),
		.dout(new_net_2919)
	);

	bfr new_net_2921_bfr_before (
		.din(new_net_2921),
		.dout(new_net_2920)
	);

	bfr new_net_2922_bfr_before (
		.din(new_net_2922),
		.dout(new_net_2921)
	);

	bfr new_net_2923_bfr_before (
		.din(new_net_2923),
		.dout(new_net_2922)
	);

	bfr new_net_2924_bfr_before (
		.din(new_net_2924),
		.dout(new_net_2923)
	);

	bfr new_net_2925_bfr_before (
		.din(new_net_2925),
		.dout(new_net_2924)
	);

	bfr new_net_2926_bfr_before (
		.din(new_net_2926),
		.dout(new_net_2925)
	);

	bfr new_net_2927_bfr_before (
		.din(new_net_2927),
		.dout(new_net_2926)
	);

	bfr new_net_2928_bfr_before (
		.din(new_net_2928),
		.dout(new_net_2927)
	);

	bfr new_net_2929_bfr_before (
		.din(new_net_2929),
		.dout(new_net_2928)
	);

	bfr new_net_2930_bfr_before (
		.din(new_net_2930),
		.dout(new_net_2929)
	);

	bfr new_net_2931_bfr_before (
		.din(new_net_2931),
		.dout(new_net_2930)
	);

	bfr new_net_2932_bfr_before (
		.din(new_net_2932),
		.dout(new_net_2931)
	);

	bfr new_net_2933_bfr_before (
		.din(new_net_2933),
		.dout(new_net_2932)
	);

	bfr new_net_2934_bfr_before (
		.din(new_net_2934),
		.dout(new_net_2933)
	);

	bfr new_net_2935_bfr_before (
		.din(new_net_2935),
		.dout(new_net_2934)
	);

	bfr new_net_2936_bfr_before (
		.din(new_net_2936),
		.dout(new_net_2935)
	);

	bfr new_net_2937_bfr_before (
		.din(new_net_2937),
		.dout(new_net_2936)
	);

	bfr new_net_2938_bfr_before (
		.din(new_net_2938),
		.dout(new_net_2937)
	);

	bfr new_net_2939_bfr_before (
		.din(new_net_2939),
		.dout(new_net_2938)
	);

	spl3L new_net_2071_v_fanout (
		.a(new_net_2071),
		.b(new_net_423),
		.c(new_net_420),
		.d(new_net_2939)
	);

	spl2 _0186__v_fanout (
		.a(_0186_),
		.b(new_net_1024),
		.c(new_net_1025)
	);

	spl2 _0249__v_fanout (
		.a(_0249_),
		.b(new_net_354),
		.c(new_net_355)
	);

	spl2 new_net_2055_v_fanout (
		.a(new_net_2055),
		.b(new_net_1451),
		.c(new_net_1450)
	);

	spl2 _1054__v_fanout (
		.a(_1054_),
		.b(new_net_1329),
		.c(new_net_1330)
	);

	spl2 new_net_3_v_fanout (
		.a(new_net_3),
		.b(new_net_2071),
		.c(new_net_2070)
	);

	bfr new_net_2940_bfr_before (
		.din(new_net_2940),
		.dout(new_net_1895)
	);

	bfr new_net_2941_bfr_before (
		.din(new_net_2941),
		.dout(new_net_2940)
	);

	bfr new_net_2942_bfr_before (
		.din(new_net_2942),
		.dout(new_net_2941)
	);

	spl2 new_net_1894_v_fanout (
		.a(new_net_1894),
		.b(new_net_1501),
		.c(new_net_2942)
	);

	bfr new_net_2943_bfr_before (
		.din(new_net_2943),
		.dout(new_net_412)
	);

	spl2 new_net_2065_v_fanout (
		.a(new_net_2065),
		.b(new_net_2943),
		.c(new_net_2066)
	);

	bfr new_net_2944_bfr_before (
		.din(new_net_2944),
		.dout(new_net_1793)
	);

	bfr new_net_2945_bfr_before (
		.din(new_net_2945),
		.dout(new_net_2944)
	);

	spl2 new_net_1792_v_fanout (
		.a(new_net_1792),
		.b(new_net_935),
		.c(new_net_2945)
	);

	spl2 _0836__v_fanout (
		.a(_0836_),
		.b(new_net_41),
		.c(new_net_42)
	);

	spl2 _0763__v_fanout (
		.a(_0763_),
		.b(new_net_2069),
		.c(new_net_2068)
	);

	bfr new_net_2946_bfr_before (
		.din(new_net_2946),
		.dout(new_net_587)
	);

	bfr new_net_2947_bfr_before (
		.din(new_net_2947),
		.dout(new_net_2946)
	);

	bfr new_net_2948_bfr_before (
		.din(new_net_2948),
		.dout(new_net_2947)
	);

	bfr new_net_2949_bfr_before (
		.din(new_net_2949),
		.dout(new_net_2948)
	);

	bfr new_net_2950_bfr_before (
		.din(new_net_2950),
		.dout(new_net_2949)
	);

	bfr new_net_2951_bfr_before (
		.din(new_net_2951),
		.dout(new_net_2950)
	);

	bfr new_net_2952_bfr_before (
		.din(new_net_2952),
		.dout(new_net_2951)
	);

	bfr new_net_2953_bfr_before (
		.din(new_net_2953),
		.dout(new_net_2952)
	);

	bfr new_net_2954_bfr_before (
		.din(new_net_2954),
		.dout(new_net_2953)
	);

	bfr new_net_2955_bfr_before (
		.din(new_net_2955),
		.dout(new_net_2954)
	);

	bfr new_net_2956_bfr_before (
		.din(new_net_2956),
		.dout(new_net_2955)
	);

	bfr new_net_2957_bfr_before (
		.din(new_net_2957),
		.dout(new_net_2956)
	);

	spl2 new_net_1919_v_fanout (
		.a(new_net_1919),
		.b(new_net_586),
		.c(new_net_2957)
	);

	spl2 _0718__v_fanout (
		.a(_0718_),
		.b(new_net_491),
		.c(new_net_492)
	);

	bfr new_net_2958_bfr_before (
		.din(new_net_2958),
		.dout(new_net_626)
	);

	bfr new_net_2959_bfr_before (
		.din(new_net_2959),
		.dout(new_net_2958)
	);

	spl2 new_net_1999_v_fanout (
		.a(new_net_1999),
		.b(new_net_2959),
		.c(new_net_622)
	);

	spl2 new_net_1975_v_fanout (
		.a(new_net_1975),
		.b(new_net_382),
		.c(new_net_1976)
	);

	spl2 new_net_2064_v_fanout (
		.a(new_net_2064),
		.b(new_net_1285),
		.c(new_net_1286)
	);

	spl2 _1104__v_fanout (
		.a(_1104_),
		.b(new_net_638),
		.c(new_net_639)
	);

	spl4L _0703__v_fanout (
		.a(_0703_),
		.b(new_net_600),
		.c(new_net_599),
		.d(new_net_598),
		.e(new_net_597)
	);

	bfr new_net_2960_bfr_before (
		.din(new_net_2960),
		.dout(new_net_1735)
	);

	spl2 new_net_1734_v_fanout (
		.a(new_net_1734),
		.b(new_net_1236),
		.c(new_net_2960)
	);

	spl2 new_net_2036_v_fanout (
		.a(new_net_2036),
		.b(new_net_977),
		.c(new_net_975)
	);

	bfr new_net_2961_bfr_after (
		.din(_1083_),
		.dout(new_net_2961)
	);

	bfr new_net_2962_bfr_after (
		.din(new_net_2961),
		.dout(new_net_2962)
	);

	bfr new_net_2963_bfr_after (
		.din(new_net_2962),
		.dout(new_net_2963)
	);

	spl2 _1083__v_fanout (
		.a(new_net_2963),
		.b(new_net_266),
		.c(new_net_267)
	);

	spl2 _1088__v_fanout (
		.a(_1088_),
		.b(new_net_701),
		.c(new_net_702)
	);

	spl2 _1218__v_fanout (
		.a(_1218_),
		.b(new_net_1491),
		.c(new_net_1492)
	);

	spl3L _0672__v_fanout (
		.a(_0672_),
		.b(new_net_1262),
		.c(new_net_1264),
		.d(new_net_1263)
	);

	spl2 new_net_1791_v_fanout (
		.a(new_net_1791),
		.b(new_net_927),
		.c(new_net_1792)
	);

	spl2 _0962__v_fanout (
		.a(_0962_),
		.b(new_net_2065),
		.c(new_net_411)
	);

	bfr new_net_2964_bfr_before (
		.din(new_net_2964),
		.dout(new_net_1818)
	);

	bfr new_net_2965_bfr_before (
		.din(new_net_2965),
		.dout(new_net_2964)
	);

	bfr new_net_2966_bfr_before (
		.din(new_net_2966),
		.dout(new_net_2965)
	);

	spl2 new_net_1817_v_fanout (
		.a(new_net_1817),
		.b(new_net_663),
		.c(new_net_2966)
	);

	spl3L _0793__v_fanout (
		.a(_0793_),
		.b(new_net_1105),
		.c(new_net_1107),
		.d(new_net_1106)
	);

	spl2 new_net_2062_v_fanout (
		.a(new_net_2062),
		.b(new_net_1642),
		.c(new_net_1643)
	);

	bfr new_net_2967_bfr_before (
		.din(new_net_2967),
		.dout(G5285)
	);

	bfr new_net_2968_bfr_before (
		.din(new_net_2968),
		.dout(new_net_2967)
	);

	bfr new_net_2969_bfr_before (
		.din(new_net_2969),
		.dout(new_net_2968)
	);

	bfr new_net_2970_bfr_before (
		.din(new_net_2970),
		.dout(new_net_2969)
	);

	bfr new_net_2971_bfr_before (
		.din(new_net_2971),
		.dout(new_net_2970)
	);

	bfr new_net_2972_bfr_before (
		.din(new_net_2972),
		.dout(new_net_2971)
	);

	bfr new_net_2973_bfr_before (
		.din(new_net_2973),
		.dout(new_net_2972)
	);

	bfr new_net_2974_bfr_before (
		.din(new_net_2974),
		.dout(new_net_2973)
	);

	bfr new_net_2975_bfr_before (
		.din(new_net_2975),
		.dout(new_net_2974)
	);

	bfr new_net_2976_bfr_before (
		.din(new_net_2976),
		.dout(new_net_2975)
	);

	bfr new_net_2977_bfr_before (
		.din(new_net_2977),
		.dout(new_net_2976)
	);

	bfr new_net_2978_bfr_before (
		.din(new_net_2978),
		.dout(new_net_2977)
	);

	bfr new_net_2979_bfr_before (
		.din(new_net_2979),
		.dout(new_net_2978)
	);

	bfr new_net_2980_bfr_before (
		.din(new_net_2980),
		.dout(new_net_2979)
	);

	bfr new_net_2981_bfr_before (
		.din(new_net_2981),
		.dout(new_net_2980)
	);

	bfr new_net_2982_bfr_before (
		.din(new_net_2982),
		.dout(new_net_2981)
	);

	bfr new_net_2983_bfr_before (
		.din(new_net_2983),
		.dout(new_net_2982)
	);

	bfr new_net_2984_bfr_before (
		.din(new_net_2984),
		.dout(new_net_2983)
	);

	bfr new_net_2985_bfr_before (
		.din(new_net_2985),
		.dout(new_net_2984)
	);

	bfr new_net_2986_bfr_before (
		.din(new_net_2986),
		.dout(new_net_2985)
	);

	bfr new_net_2987_bfr_before (
		.din(new_net_2987),
		.dout(new_net_2986)
	);

	bfr new_net_2988_bfr_before (
		.din(new_net_2988),
		.dout(new_net_2987)
	);

	bfr new_net_2989_bfr_before (
		.din(new_net_2989),
		.dout(new_net_2988)
	);

	bfr new_net_2990_bfr_before (
		.din(new_net_2990),
		.dout(new_net_2989)
	);

	bfr new_net_2991_bfr_before (
		.din(new_net_2991),
		.dout(new_net_2990)
	);

	spl3L new_net_2063_v_fanout (
		.a(new_net_2063),
		.b(new_net_1639),
		.c(new_net_1640),
		.d(new_net_2991)
	);

	spl2 new_net_2057_v_fanout (
		.a(new_net_2057),
		.b(new_net_78),
		.c(new_net_77)
	);

	spl2 _0018__v_fanout (
		.a(_0018_),
		.b(new_net_1058),
		.c(new_net_1059)
	);

	spl3L _0771__v_fanout (
		.a(_0771_),
		.b(new_net_1678),
		.c(new_net_1679),
		.d(new_net_1680)
	);

	bfr new_net_2992_bfr_before (
		.din(new_net_2992),
		.dout(new_net_1579)
	);

	bfr new_net_2993_bfr_before (
		.din(new_net_2993),
		.dout(new_net_2992)
	);

	bfr new_net_2994_bfr_before (
		.din(new_net_2994),
		.dout(new_net_2993)
	);

	bfr new_net_2995_bfr_before (
		.din(new_net_2995),
		.dout(new_net_2994)
	);

	bfr new_net_2996_bfr_before (
		.din(new_net_2996),
		.dout(new_net_2995)
	);

	bfr new_net_2997_bfr_before (
		.din(new_net_2997),
		.dout(new_net_2996)
	);

	bfr new_net_2998_bfr_before (
		.din(new_net_2998),
		.dout(new_net_2997)
	);

	bfr new_net_2999_bfr_before (
		.din(new_net_2999),
		.dout(new_net_2998)
	);

	bfr new_net_3000_bfr_before (
		.din(new_net_3000),
		.dout(new_net_2999)
	);

	spl2 _0957__v_fanout (
		.a(_0957_),
		.b(new_net_3000),
		.c(new_net_1580)
	);

	bfr new_net_3001_bfr_before (
		.din(new_net_3001),
		.dout(new_net_1734)
	);

	spl2 new_net_1733_v_fanout (
		.a(new_net_1733),
		.b(new_net_1227),
		.c(new_net_3001)
	);

	spl3L _1050__v_fanout (
		.a(_1050_),
		.b(new_net_195),
		.c(new_net_197),
		.d(new_net_196)
	);

	bfr new_net_3002_bfr_before (
		.din(new_net_3002),
		.dout(new_net_1919)
	);

	spl2 new_net_1918_v_fanout (
		.a(new_net_1918),
		.b(new_net_3002),
		.c(new_net_588)
	);

	bfr new_net_3003_bfr_before (
		.din(new_net_3003),
		.dout(new_net_700)
	);

	spl3L _0762__v_fanout (
		.a(_0762_),
		.b(new_net_698),
		.c(new_net_3003),
		.d(new_net_699)
	);

	bfr new_net_3004_bfr_before (
		.din(new_net_3004),
		.dout(new_net_1581)
	);

	spl2 _0815__v_fanout (
		.a(_0815_),
		.b(new_net_3004),
		.c(new_net_1582)
	);

	spl2 new_net_18_v_fanout (
		.a(new_net_18),
		.b(new_net_2062),
		.c(new_net_2063)
	);

	bfr new_net_3005_bfr_after (
		.din(_0244_),
		.dout(new_net_3005)
	);

	bfr new_net_3006_bfr_before (
		.din(new_net_3006),
		.dout(new_net_2064)
	);

	spl2 _0244__v_fanout (
		.a(new_net_3005),
		.b(new_net_3006),
		.c(new_net_1287)
	);

	bfr new_net_3007_bfr_after (
		.din(_1098_),
		.dout(new_net_3007)
	);

	bfr new_net_3008_bfr_after (
		.din(new_net_3007),
		.dout(new_net_3008)
	);

	spl2 _1098__v_fanout (
		.a(new_net_3008),
		.b(new_net_70),
		.c(new_net_71)
	);

	spl2 _0183__v_fanout (
		.a(_0183_),
		.b(new_net_1535),
		.c(new_net_1536)
	);

	spl2 _0213__v_fanout (
		.a(_0213_),
		.b(new_net_545),
		.c(new_net_546)
	);

	spl2 _0620__v_fanout (
		.a(_0620_),
		.b(new_net_216),
		.c(new_net_217)
	);

	bfr new_net_3009_bfr_before (
		.din(new_net_3009),
		.dout(new_net_1927)
	);

	bfr new_net_3010_bfr_before (
		.din(new_net_3010),
		.dout(new_net_3009)
	);

	spl2 new_net_1926_v_fanout (
		.a(new_net_1926),
		.b(new_net_437),
		.c(new_net_3010)
	);

	spl2 new_net_2038_v_fanout (
		.a(new_net_2038),
		.b(new_net_167),
		.c(new_net_169)
	);

	spl2 _0671__v_fanout (
		.a(_0671_),
		.b(new_net_608),
		.c(new_net_609)
	);

	bfr new_net_3011_bfr_before (
		.din(new_net_3011),
		.dout(new_net_1182)
	);

	bfr new_net_3012_bfr_before (
		.din(new_net_3012),
		.dout(new_net_3011)
	);

	spl3L new_net_2048_v_fanout (
		.a(new_net_2048),
		.b(new_net_1183),
		.c(new_net_1181),
		.d(new_net_3012)
	);

	bfr new_net_3013_bfr_before (
		.din(new_net_3013),
		.dout(new_net_1960)
	);

	bfr new_net_3014_bfr_before (
		.din(new_net_3014),
		.dout(new_net_3013)
	);

	spl2 new_net_1959_v_fanout (
		.a(new_net_1959),
		.b(new_net_3014),
		.c(new_net_681)
	);

	bfr new_net_3015_bfr_before (
		.din(new_net_3015),
		.dout(new_net_2059)
	);

	bfr new_net_3016_bfr_before (
		.din(new_net_3016),
		.dout(new_net_3015)
	);

	bfr new_net_3017_bfr_before (
		.din(new_net_3017),
		.dout(new_net_3016)
	);

	spl2 new_net_2058_v_fanout (
		.a(new_net_2058),
		.b(new_net_631),
		.c(new_net_3017)
	);

	bfr new_net_3018_bfr_after (
		.din(_0246_),
		.dout(new_net_3018)
	);

	bfr new_net_3019_bfr_after (
		.din(new_net_3018),
		.dout(new_net_3019)
	);

	spl2 _0246__v_fanout (
		.a(new_net_3019),
		.b(new_net_293),
		.c(new_net_294)
	);

	spl2 _0079__v_fanout (
		.a(_0079_),
		.b(new_net_1028),
		.c(new_net_1029)
	);

	bfr new_net_3020_bfr_before (
		.din(new_net_3020),
		.dout(new_net_2036)
	);

	spl2 new_net_2035_v_fanout (
		.a(new_net_2035),
		.b(new_net_973),
		.c(new_net_3020)
	);

	spl2 _0159__v_fanout (
		.a(_0159_),
		.b(new_net_80),
		.c(new_net_81)
	);

	spl3L new_net_2061_v_fanout (
		.a(new_net_2061),
		.b(new_net_578),
		.c(new_net_582),
		.d(new_net_579)
	);

	bfr new_net_3021_bfr_before (
		.din(new_net_3021),
		.dout(G5248)
	);

	bfr new_net_3022_bfr_before (
		.din(new_net_3022),
		.dout(new_net_3021)
	);

	bfr new_net_3023_bfr_before (
		.din(new_net_3023),
		.dout(new_net_3022)
	);

	bfr new_net_3024_bfr_before (
		.din(new_net_3024),
		.dout(new_net_3023)
	);

	bfr new_net_3025_bfr_before (
		.din(new_net_3025),
		.dout(new_net_3024)
	);

	bfr new_net_3026_bfr_before (
		.din(new_net_3026),
		.dout(new_net_3025)
	);

	bfr new_net_3027_bfr_before (
		.din(new_net_3027),
		.dout(new_net_3026)
	);

	bfr new_net_3028_bfr_before (
		.din(new_net_3028),
		.dout(new_net_3027)
	);

	bfr new_net_3029_bfr_before (
		.din(new_net_3029),
		.dout(new_net_3028)
	);

	bfr new_net_3030_bfr_before (
		.din(new_net_3030),
		.dout(new_net_3029)
	);

	bfr new_net_3031_bfr_before (
		.din(new_net_3031),
		.dout(new_net_3030)
	);

	bfr new_net_3032_bfr_before (
		.din(new_net_3032),
		.dout(new_net_3031)
	);

	bfr new_net_3033_bfr_before (
		.din(new_net_3033),
		.dout(new_net_3032)
	);

	bfr new_net_3034_bfr_before (
		.din(new_net_3034),
		.dout(new_net_3033)
	);

	bfr new_net_3035_bfr_before (
		.din(new_net_3035),
		.dout(new_net_3034)
	);

	bfr new_net_3036_bfr_before (
		.din(new_net_3036),
		.dout(new_net_3035)
	);

	bfr new_net_3037_bfr_before (
		.din(new_net_3037),
		.dout(new_net_3036)
	);

	bfr new_net_3038_bfr_before (
		.din(new_net_3038),
		.dout(new_net_3037)
	);

	bfr new_net_3039_bfr_before (
		.din(new_net_3039),
		.dout(new_net_3038)
	);

	bfr new_net_3040_bfr_before (
		.din(new_net_3040),
		.dout(new_net_3039)
	);

	bfr new_net_3041_bfr_before (
		.din(new_net_3041),
		.dout(new_net_3040)
	);

	bfr new_net_3042_bfr_before (
		.din(new_net_3042),
		.dout(new_net_3041)
	);

	bfr new_net_3043_bfr_before (
		.din(new_net_3043),
		.dout(new_net_3042)
	);

	bfr new_net_3044_bfr_before (
		.din(new_net_3044),
		.dout(new_net_3043)
	);

	bfr new_net_3045_bfr_before (
		.din(new_net_3045),
		.dout(new_net_3044)
	);

	bfr new_net_3046_bfr_before (
		.din(new_net_3046),
		.dout(new_net_3045)
	);

	bfr new_net_3047_bfr_before (
		.din(new_net_3047),
		.dout(new_net_3046)
	);

	spl2 new_net_2060_v_fanout (
		.a(new_net_2060),
		.b(new_net_3047),
		.c(new_net_580)
	);

	spl2 _1235__v_fanout (
		.a(_1235_),
		.b(new_net_1507),
		.c(new_net_1508)
	);

	bfr new_net_3048_bfr_before (
		.din(new_net_3048),
		.dout(new_net_1953)
	);

	bfr new_net_3049_bfr_before (
		.din(new_net_3049),
		.dout(new_net_3048)
	);

	spl2 new_net_1952_v_fanout (
		.a(new_net_1952),
		.b(new_net_3049),
		.c(new_net_1352)
	);

	bfr new_net_3050_bfr_before (
		.din(new_net_3050),
		.dout(new_net_1968)
	);

	bfr new_net_3051_bfr_before (
		.din(new_net_3051),
		.dout(new_net_3050)
	);

	spl2 new_net_1967_v_fanout (
		.a(new_net_1967),
		.b(new_net_3051),
		.c(new_net_805)
	);

	bfr new_net_3052_bfr_before (
		.din(new_net_3052),
		.dout(new_net_884)
	);

	bfr new_net_3053_bfr_before (
		.din(new_net_3053),
		.dout(new_net_3052)
	);

	spl2 _1090__v_fanout (
		.a(_1090_),
		.b(new_net_3053),
		.c(new_net_885)
	);

	spl2 _0715__v_fanout (
		.a(_0715_),
		.b(new_net_178),
		.c(new_net_179)
	);

	bfr new_net_3054_bfr_before (
		.din(new_net_3054),
		.dout(new_net_1204)
	);

	spl2 new_net_1732_v_fanout (
		.a(new_net_1732),
		.b(new_net_1733),
		.c(new_net_3054)
	);

	bfr new_net_3055_bfr_before (
		.din(new_net_3055),
		.dout(new_net_547)
	);

	bfr new_net_3056_bfr_before (
		.din(new_net_3056),
		.dout(new_net_3055)
	);

	spl2 _1086__v_fanout (
		.a(_1086_),
		.b(new_net_3056),
		.c(new_net_548)
	);

	bfr new_net_3057_bfr_before (
		.din(new_net_3057),
		.dout(new_net_2054)
	);

	bfr new_net_3058_bfr_before (
		.din(new_net_3058),
		.dout(new_net_3057)
	);

	bfr new_net_3059_bfr_before (
		.din(new_net_3059),
		.dout(new_net_3058)
	);

	bfr new_net_3060_bfr_before (
		.din(new_net_3060),
		.dout(new_net_3059)
	);

	bfr new_net_3061_bfr_before (
		.din(new_net_3061),
		.dout(new_net_3060)
	);

	bfr new_net_3062_bfr_before (
		.din(new_net_3062),
		.dout(new_net_3061)
	);

	bfr new_net_3063_bfr_before (
		.din(new_net_3063),
		.dout(new_net_3062)
	);

	bfr new_net_3064_bfr_before (
		.din(new_net_3064),
		.dout(new_net_3063)
	);

	bfr new_net_3065_bfr_before (
		.din(new_net_3065),
		.dout(new_net_3064)
	);

	bfr new_net_3066_bfr_before (
		.din(new_net_3066),
		.dout(new_net_3065)
	);

	bfr new_net_3067_bfr_before (
		.din(new_net_3067),
		.dout(new_net_3066)
	);

	bfr new_net_3068_bfr_before (
		.din(new_net_3068),
		.dout(new_net_3067)
	);

	spl2 new_net_2053_v_fanout (
		.a(new_net_2053),
		.b(new_net_1443),
		.c(new_net_3068)
	);

	bfr new_net_3069_bfr_before (
		.din(new_net_3069),
		.dout(new_net_1983)
	);

	bfr new_net_3070_bfr_before (
		.din(new_net_3070),
		.dout(new_net_3069)
	);

	spl2 new_net_1982_v_fanout (
		.a(new_net_1982),
		.b(new_net_1573),
		.c(new_net_3070)
	);

	bfr new_net_3071_bfr_before (
		.din(new_net_3071),
		.dout(new_net_1791)
	);

	spl2 new_net_1790_v_fanout (
		.a(new_net_1790),
		.b(new_net_936),
		.c(new_net_3071)
	);

	bfr new_net_3072_bfr_before (
		.din(new_net_3072),
		.dout(new_net_1943)
	);

	bfr new_net_3073_bfr_before (
		.din(new_net_3073),
		.dout(new_net_3072)
	);

	spl2 new_net_1942_v_fanout (
		.a(new_net_1942),
		.b(new_net_1152),
		.c(new_net_3073)
	);

	bfr new_net_3074_bfr_before (
		.din(new_net_3074),
		.dout(G5242)
	);

	bfr new_net_3075_bfr_before (
		.din(new_net_3075),
		.dout(new_net_3074)
	);

	bfr new_net_3076_bfr_before (
		.din(new_net_3076),
		.dout(new_net_3075)
	);

	bfr new_net_3077_bfr_before (
		.din(new_net_3077),
		.dout(new_net_3076)
	);

	bfr new_net_3078_bfr_before (
		.din(new_net_3078),
		.dout(new_net_3077)
	);

	bfr new_net_3079_bfr_before (
		.din(new_net_3079),
		.dout(new_net_3078)
	);

	bfr new_net_3080_bfr_before (
		.din(new_net_3080),
		.dout(new_net_3079)
	);

	bfr new_net_3081_bfr_before (
		.din(new_net_3081),
		.dout(new_net_3080)
	);

	bfr new_net_3082_bfr_before (
		.din(new_net_3082),
		.dout(new_net_3081)
	);

	bfr new_net_3083_bfr_before (
		.din(new_net_3083),
		.dout(new_net_3082)
	);

	bfr new_net_3084_bfr_before (
		.din(new_net_3084),
		.dout(new_net_3083)
	);

	bfr new_net_3085_bfr_before (
		.din(new_net_3085),
		.dout(new_net_3084)
	);

	bfr new_net_3086_bfr_before (
		.din(new_net_3086),
		.dout(new_net_3085)
	);

	bfr new_net_3087_bfr_before (
		.din(new_net_3087),
		.dout(new_net_3086)
	);

	bfr new_net_3088_bfr_before (
		.din(new_net_3088),
		.dout(new_net_3087)
	);

	bfr new_net_3089_bfr_before (
		.din(new_net_3089),
		.dout(new_net_3088)
	);

	bfr new_net_3090_bfr_before (
		.din(new_net_3090),
		.dout(new_net_3089)
	);

	bfr new_net_3091_bfr_before (
		.din(new_net_3091),
		.dout(new_net_3090)
	);

	bfr new_net_3092_bfr_before (
		.din(new_net_3092),
		.dout(new_net_3091)
	);

	bfr new_net_3093_bfr_before (
		.din(new_net_3093),
		.dout(new_net_3092)
	);

	bfr new_net_3094_bfr_before (
		.din(new_net_3094),
		.dout(new_net_3093)
	);

	bfr new_net_3095_bfr_before (
		.din(new_net_3095),
		.dout(new_net_3094)
	);

	bfr new_net_3096_bfr_before (
		.din(new_net_3096),
		.dout(new_net_3095)
	);

	bfr new_net_3097_bfr_before (
		.din(new_net_3097),
		.dout(new_net_3096)
	);

	bfr new_net_3098_bfr_before (
		.din(new_net_3098),
		.dout(new_net_3097)
	);

	bfr new_net_3099_bfr_before (
		.din(new_net_3099),
		.dout(new_net_3098)
	);

	bfr new_net_3100_bfr_before (
		.din(new_net_3100),
		.dout(new_net_3099)
	);

	bfr new_net_3101_bfr_before (
		.din(new_net_3101),
		.dout(new_net_3100)
	);

	spl2 new_net_15_v_fanout (
		.a(new_net_15),
		.b(new_net_3101),
		.c(new_net_1000)
	);

	spl4L _0769__v_fanout (
		.a(_0769_),
		.b(new_net_630),
		.c(new_net_633),
		.d(new_net_634),
		.e(new_net_2058)
	);

	spl2 _1215__v_fanout (
		.a(_1215_),
		.b(new_net_1241),
		.c(new_net_1242)
	);

	bfr new_net_3102_bfr_before (
		.din(new_net_3102),
		.dout(new_net_1157)
	);

	bfr new_net_3103_bfr_before (
		.din(new_net_3103),
		.dout(new_net_3102)
	);

	bfr new_net_3104_bfr_before (
		.din(new_net_3104),
		.dout(new_net_3103)
	);

	bfr new_net_3105_bfr_before (
		.din(new_net_3105),
		.dout(new_net_3104)
	);

	bfr new_net_3106_bfr_before (
		.din(new_net_3106),
		.dout(new_net_3105)
	);

	bfr new_net_3107_bfr_before (
		.din(new_net_3107),
		.dout(new_net_3106)
	);

	bfr new_net_3108_bfr_before (
		.din(new_net_3108),
		.dout(new_net_3107)
	);

	bfr new_net_3109_bfr_before (
		.din(new_net_3109),
		.dout(new_net_3108)
	);

	bfr new_net_3110_bfr_before (
		.din(new_net_3110),
		.dout(new_net_3109)
	);

	bfr new_net_3111_bfr_before (
		.din(new_net_3111),
		.dout(new_net_3110)
	);

	spl2 _0970__v_fanout (
		.a(_0970_),
		.b(new_net_3111),
		.c(new_net_1158)
	);

	bfr new_net_3112_bfr_before (
		.din(new_net_3112),
		.dout(new_net_1027)
	);

	bfr new_net_3113_bfr_before (
		.din(new_net_3113),
		.dout(new_net_3112)
	);

	bfr new_net_3114_bfr_before (
		.din(new_net_3114),
		.dout(new_net_3113)
	);

	bfr new_net_3115_bfr_before (
		.din(new_net_3115),
		.dout(new_net_3114)
	);

	spl2 _0643__v_fanout (
		.a(_0643_),
		.b(new_net_1026),
		.c(new_net_3115)
	);

	spl2 _0012__v_fanout (
		.a(_0012_),
		.b(new_net_601),
		.c(new_net_602)
	);

	bfr new_net_3116_bfr_after (
		.din(_0070_),
		.dout(new_net_3116)
	);

	spl2 _0070__v_fanout (
		.a(new_net_3116),
		.b(new_net_161),
		.c(new_net_162)
	);

	spl2 _0956__v_fanout (
		.a(_0956_),
		.b(new_net_1435),
		.c(new_net_1436)
	);

	bfr new_net_3117_bfr_before (
		.din(new_net_3117),
		.dout(new_net_2046)
	);

	bfr new_net_3118_bfr_before (
		.din(new_net_3118),
		.dout(new_net_3117)
	);

	bfr new_net_3119_bfr_before (
		.din(new_net_3119),
		.dout(new_net_3118)
	);

	bfr new_net_3120_bfr_before (
		.din(new_net_3120),
		.dout(new_net_3119)
	);

	spl2 new_net_2045_v_fanout (
		.a(new_net_2045),
		.b(new_net_1651),
		.c(new_net_3120)
	);

	bfr new_net_3121_bfr_before (
		.din(new_net_3121),
		.dout(new_net_1975)
	);

	spl2 new_net_1974_v_fanout (
		.a(new_net_1974),
		.b(new_net_388),
		.c(new_net_3121)
	);

	spl2 _0015__v_fanout (
		.a(_0015_),
		.b(new_net_775),
		.c(new_net_776)
	);

	spl2 _0814__v_fanout (
		.a(_0814_),
		.b(new_net_1540),
		.c(new_net_1541)
	);

	bfr new_net_3122_bfr_before (
		.din(new_net_3122),
		.dout(new_net_1134)
	);

	bfr new_net_3123_bfr_before (
		.din(new_net_3123),
		.dout(new_net_3122)
	);

	bfr new_net_3124_bfr_before (
		.din(new_net_3124),
		.dout(new_net_3123)
	);

	bfr new_net_3125_bfr_before (
		.din(new_net_3125),
		.dout(new_net_3124)
	);

	bfr new_net_3126_bfr_before (
		.din(new_net_3126),
		.dout(new_net_3125)
	);

	bfr new_net_3127_bfr_before (
		.din(new_net_3127),
		.dout(new_net_3126)
	);

	bfr new_net_3128_bfr_before (
		.din(new_net_3128),
		.dout(new_net_3127)
	);

	bfr new_net_3129_bfr_before (
		.din(new_net_3129),
		.dout(new_net_3128)
	);

	bfr new_net_3130_bfr_before (
		.din(new_net_3130),
		.dout(new_net_3129)
	);

	bfr new_net_3131_bfr_before (
		.din(new_net_3131),
		.dout(new_net_3130)
	);

	spl2 new_net_2028_v_fanout (
		.a(new_net_2028),
		.b(new_net_1132),
		.c(new_net_3131)
	);

	spl2 new_net_2056_v_fanout (
		.a(new_net_2056),
		.b(new_net_865),
		.c(new_net_864)
	);

	spl2 _1081__v_fanout (
		.a(_1081_),
		.b(new_net_68),
		.c(new_net_69)
	);

	spl2 new_net_4_v_fanout (
		.a(new_net_4),
		.b(new_net_2060),
		.c(new_net_2061)
	);

	spl2 new_net_2025_v_fanout (
		.a(new_net_2025),
		.b(new_net_1585),
		.c(new_net_1587)
	);

	bfr new_net_3132_bfr_after (
		.din(_1118_),
		.dout(new_net_3132)
	);

	bfr new_net_3133_bfr_after (
		.din(new_net_3132),
		.dout(new_net_3133)
	);

	bfr new_net_3134_bfr_after (
		.din(new_net_3133),
		.dout(new_net_3134)
	);

	bfr new_net_3135_bfr_after (
		.din(new_net_3134),
		.dout(new_net_3135)
	);

	bfr new_net_3136_bfr_after (
		.din(new_net_3135),
		.dout(new_net_3136)
	);

	bfr new_net_3137_bfr_after (
		.din(new_net_3136),
		.dout(new_net_3137)
	);

	bfr new_net_3138_bfr_after (
		.din(new_net_3137),
		.dout(new_net_3138)
	);

	bfr new_net_3139_bfr_after (
		.din(new_net_3138),
		.dout(new_net_3139)
	);

	bfr new_net_3140_bfr_after (
		.din(new_net_3139),
		.dout(new_net_3140)
	);

	bfr new_net_3141_bfr_after (
		.din(new_net_3140),
		.dout(new_net_3141)
	);

	bfr new_net_3142_bfr_after (
		.din(new_net_3141),
		.dout(new_net_3142)
	);

	bfr new_net_3143_bfr_after (
		.din(new_net_3142),
		.dout(new_net_3143)
	);

	bfr new_net_3144_bfr_after (
		.din(new_net_3143),
		.dout(new_net_3144)
	);

	spl2 _1118__v_fanout (
		.a(new_net_3144),
		.b(new_net_527),
		.c(new_net_528)
	);

	bfr new_net_3145_bfr_after (
		.din(_1161_),
		.dout(new_net_3145)
	);

	bfr new_net_3146_bfr_after (
		.din(new_net_3145),
		.dout(new_net_3146)
	);

	bfr new_net_3147_bfr_after (
		.din(new_net_3146),
		.dout(new_net_3147)
	);

	spl2 _1161__v_fanout (
		.a(new_net_3147),
		.b(new_net_869),
		.c(new_net_870)
	);

	spl3L _0748__v_fanout (
		.a(_0748_),
		.b(new_net_970),
		.c(new_net_971),
		.d(new_net_972)
	);

	bfr new_net_3148_bfr_before (
		.din(new_net_3148),
		.dout(new_net_253)
	);

	bfr new_net_3149_bfr_before (
		.din(new_net_3149),
		.dout(new_net_3148)
	);

	bfr new_net_3150_bfr_before (
		.din(new_net_3150),
		.dout(new_net_3149)
	);

	bfr new_net_3151_bfr_before (
		.din(new_net_3151),
		.dout(new_net_3150)
	);

	bfr new_net_3152_bfr_before (
		.din(new_net_3152),
		.dout(new_net_3151)
	);

	bfr new_net_3153_bfr_before (
		.din(new_net_3153),
		.dout(new_net_3152)
	);

	bfr new_net_3154_bfr_before (
		.din(new_net_3154),
		.dout(new_net_3153)
	);

	bfr new_net_3155_bfr_before (
		.din(new_net_3155),
		.dout(new_net_3154)
	);

	bfr new_net_3156_bfr_before (
		.din(new_net_3156),
		.dout(new_net_3155)
	);

	bfr new_net_3157_bfr_before (
		.din(new_net_3157),
		.dout(new_net_3156)
	);

	spl2 _0874__v_fanout (
		.a(_0874_),
		.b(new_net_3157),
		.c(new_net_254)
	);

	bfr new_net_3158_bfr_after (
		.din(_0195_),
		.dout(new_net_3158)
	);

	bfr new_net_3159_bfr_after (
		.din(new_net_3158),
		.dout(new_net_3159)
	);

	bfr new_net_3160_bfr_after (
		.din(new_net_3159),
		.dout(new_net_3160)
	);

	spl2 _0195__v_fanout (
		.a(new_net_3160),
		.b(new_net_137),
		.c(new_net_138)
	);

	bfr new_net_3161_bfr_after (
		.din(_1064_),
		.dout(new_net_3161)
	);

	bfr new_net_3162_bfr_after (
		.din(new_net_3161),
		.dout(new_net_3162)
	);

	bfr new_net_3163_bfr_after (
		.din(new_net_3162),
		.dout(new_net_3163)
	);

	bfr new_net_3164_bfr_after (
		.din(new_net_3163),
		.dout(new_net_3164)
	);

	spl2 _1064__v_fanout (
		.a(new_net_3164),
		.b(new_net_1577),
		.c(new_net_1578)
	);

	bfr new_net_3165_bfr_before (
		.din(new_net_3165),
		.dout(new_net_51)
	);

	bfr new_net_3166_bfr_before (
		.din(new_net_3166),
		.dout(new_net_3165)
	);

	bfr new_net_3167_bfr_before (
		.din(new_net_3167),
		.dout(new_net_3166)
	);

	spl2 new_net_1784_v_fanout (
		.a(new_net_1784),
		.b(new_net_52),
		.c(new_net_3167)
	);

	bfr new_net_3168_bfr_before (
		.din(new_net_3168),
		.dout(new_net_1347)
	);

	bfr new_net_3169_bfr_before (
		.din(new_net_3169),
		.dout(new_net_3168)
	);

	bfr new_net_3170_bfr_before (
		.din(new_net_3170),
		.dout(new_net_3169)
	);

	bfr new_net_3171_bfr_before (
		.din(new_net_3171),
		.dout(new_net_3170)
	);

	spl2 new_net_2023_v_fanout (
		.a(new_net_2023),
		.b(new_net_3171),
		.c(new_net_1346)
	);

	spl2 _0174__v_fanout (
		.a(_0174_),
		.b(new_net_1363),
		.c(new_net_1364)
	);

	bfr new_net_3172_bfr_before (
		.din(new_net_3172),
		.dout(new_net_1790)
	);

	spl2 new_net_1789_v_fanout (
		.a(new_net_1789),
		.b(new_net_937),
		.c(new_net_3172)
	);

	bfr new_net_3173_bfr_after (
		.din(_1101_),
		.dout(new_net_3173)
	);

	bfr new_net_3174_bfr_after (
		.din(new_net_3173),
		.dout(new_net_3174)
	);

	spl2 _1101__v_fanout (
		.a(new_net_3174),
		.b(new_net_372),
		.c(new_net_373)
	);

	spl2 _1084__v_fanout (
		.a(_1084_),
		.b(new_net_368),
		.c(new_net_369)
	);

	spl3L _0619__v_fanout (
		.a(_0619_),
		.b(new_net_398),
		.c(new_net_400),
		.d(new_net_399)
	);

	spl2 _0210__v_fanout (
		.a(_0210_),
		.b(new_net_444),
		.c(new_net_445)
	);

	spl2 _0180__v_fanout (
		.a(_0180_),
		.b(new_net_1441),
		.c(new_net_1442)
	);

	bfr new_net_3175_bfr_after (
		.din(_0165_),
		.dout(new_net_3175)
	);

	bfr new_net_3176_bfr_after (
		.din(new_net_3175),
		.dout(new_net_3176)
	);

	bfr new_net_3177_bfr_after (
		.din(new_net_3176),
		.dout(new_net_3177)
	);

	spl2 _0165__v_fanout (
		.a(new_net_3177),
		.b(new_net_1184),
		.c(new_net_1185)
	);

	spl2 _1085__v_fanout (
		.a(_1085_),
		.b(new_net_475),
		.c(new_net_476)
	);

	spl2 new_net_2044_v_fanout (
		.a(new_net_2044),
		.b(new_net_722),
		.c(new_net_723)
	);

	bfr new_net_3178_bfr_after (
		.din(_0739_),
		.dout(new_net_3178)
	);

	bfr new_net_3179_bfr_after (
		.din(new_net_3178),
		.dout(new_net_3179)
	);

	bfr new_net_3180_bfr_after (
		.din(new_net_3179),
		.dout(new_net_3180)
	);

	bfr new_net_3181_bfr_after (
		.din(new_net_3180),
		.dout(new_net_3181)
	);

	spl3L _0739__v_fanout (
		.a(new_net_3181),
		.b(new_net_76),
		.c(new_net_79),
		.d(new_net_2057)
	);

	bfr new_net_3182_bfr_before (
		.din(new_net_3182),
		.dout(new_net_2041)
	);

	bfr new_net_3183_bfr_before (
		.din(new_net_3183),
		.dout(new_net_3182)
	);

	bfr new_net_3184_bfr_before (
		.din(new_net_3184),
		.dout(new_net_3183)
	);

	bfr new_net_3185_bfr_before (
		.din(new_net_3185),
		.dout(new_net_3184)
	);

	bfr new_net_3186_bfr_before (
		.din(new_net_3186),
		.dout(new_net_3185)
	);

	bfr new_net_3187_bfr_before (
		.din(new_net_3187),
		.dout(new_net_3186)
	);

	bfr new_net_3188_bfr_before (
		.din(new_net_3188),
		.dout(new_net_3187)
	);

	bfr new_net_3189_bfr_before (
		.din(new_net_3189),
		.dout(new_net_3188)
	);

	bfr new_net_3190_bfr_before (
		.din(new_net_3190),
		.dout(new_net_3189)
	);

	bfr new_net_3191_bfr_before (
		.din(new_net_3191),
		.dout(new_net_3190)
	);

	bfr new_net_3192_bfr_before (
		.din(new_net_3192),
		.dout(new_net_3191)
	);

	bfr new_net_3193_bfr_before (
		.din(new_net_3193),
		.dout(new_net_3192)
	);

	bfr new_net_3194_bfr_before (
		.din(new_net_3194),
		.dout(new_net_3193)
	);

	bfr new_net_3195_bfr_before (
		.din(new_net_3195),
		.dout(new_net_3194)
	);

	spl2 new_net_2040_v_fanout (
		.a(new_net_2040),
		.b(new_net_389),
		.c(new_net_3195)
	);

	bfr new_net_3196_bfr_before (
		.din(new_net_3196),
		.dout(new_net_1321)
	);

	bfr new_net_3197_bfr_before (
		.din(new_net_3197),
		.dout(new_net_3196)
	);

	bfr new_net_3198_bfr_before (
		.din(new_net_3198),
		.dout(new_net_3197)
	);

	spl2 _0675__v_fanout (
		.a(_0675_),
		.b(new_net_1320),
		.c(new_net_3198)
	);

	bfr new_net_3199_bfr_before (
		.din(new_net_3199),
		.dout(new_net_199)
	);

	bfr new_net_3200_bfr_before (
		.din(new_net_3200),
		.dout(new_net_3199)
	);

	bfr new_net_3201_bfr_before (
		.din(new_net_3201),
		.dout(new_net_3200)
	);

	bfr new_net_3202_bfr_before (
		.din(new_net_3202),
		.dout(new_net_3201)
	);

	bfr new_net_3203_bfr_before (
		.din(new_net_3203),
		.dout(new_net_3202)
	);

	bfr new_net_3204_bfr_before (
		.din(new_net_3204),
		.dout(new_net_3203)
	);

	bfr new_net_3205_bfr_before (
		.din(new_net_3205),
		.dout(new_net_3204)
	);

	bfr new_net_3206_bfr_before (
		.din(new_net_3206),
		.dout(new_net_3205)
	);

	bfr new_net_3207_bfr_before (
		.din(new_net_3207),
		.dout(new_net_3206)
	);

	bfr new_net_3208_bfr_before (
		.din(new_net_3208),
		.dout(new_net_3207)
	);

	bfr new_net_3209_bfr_before (
		.din(new_net_3209),
		.dout(new_net_3208)
	);

	bfr new_net_3210_bfr_before (
		.din(new_net_3210),
		.dout(new_net_3209)
	);

	bfr new_net_3211_bfr_before (
		.din(new_net_3211),
		.dout(new_net_3210)
	);

	spl4L _0955__v_fanout (
		.a(_0955_),
		.b(new_net_200),
		.c(new_net_3211),
		.d(new_net_201),
		.e(new_net_198)
	);

	spl2 _1247__v_fanout (
		.a(_1247_),
		.b(new_net_1631),
		.c(new_net_1632)
	);

	bfr new_net_3212_bfr_before (
		.din(new_net_3212),
		.dout(new_net_1600)
	);

	bfr new_net_3213_bfr_before (
		.din(new_net_3213),
		.dout(new_net_3212)
	);

	bfr new_net_3214_bfr_before (
		.din(new_net_3214),
		.dout(new_net_3213)
	);

	spl2 new_net_2026_v_fanout (
		.a(new_net_2026),
		.b(new_net_1599),
		.c(new_net_3214)
	);

	bfr new_net_3215_bfr_before (
		.din(new_net_3215),
		.dout(new_net_606)
	);

	bfr new_net_3216_bfr_before (
		.din(new_net_3216),
		.dout(new_net_3215)
	);

	spl2 _0761__v_fanout (
		.a(_0761_),
		.b(new_net_3216),
		.c(new_net_607)
	);

	bfr new_net_3217_bfr_before (
		.din(new_net_3217),
		.dout(new_net_2056)
	);

	spl3L _0747__v_fanout (
		.a(_0747_),
		.b(new_net_863),
		.c(new_net_866),
		.d(new_net_3217)
	);

	bfr new_net_3218_bfr_after (
		.din(_0670_),
		.dout(new_net_3218)
	);

	bfr new_net_3219_bfr_before (
		.din(new_net_3219),
		.dout(new_net_1193)
	);

	bfr new_net_3220_bfr_before (
		.din(new_net_3220),
		.dout(new_net_3219)
	);

	bfr new_net_3221_bfr_before (
		.din(new_net_3221),
		.dout(new_net_3220)
	);

	bfr new_net_3222_bfr_before (
		.din(new_net_3222),
		.dout(new_net_3221)
	);

	spl2 _0670__v_fanout (
		.a(new_net_3218),
		.b(new_net_1192),
		.c(new_net_3222)
	);

	bfr new_net_3223_bfr_before (
		.din(new_net_3223),
		.dout(G5251)
	);

	bfr new_net_3224_bfr_before (
		.din(new_net_3224),
		.dout(new_net_3223)
	);

	bfr new_net_3225_bfr_before (
		.din(new_net_3225),
		.dout(new_net_3224)
	);

	bfr new_net_3226_bfr_before (
		.din(new_net_3226),
		.dout(new_net_3225)
	);

	bfr new_net_3227_bfr_before (
		.din(new_net_3227),
		.dout(new_net_3226)
	);

	bfr new_net_3228_bfr_before (
		.din(new_net_3228),
		.dout(new_net_3227)
	);

	bfr new_net_3229_bfr_before (
		.din(new_net_3229),
		.dout(new_net_3228)
	);

	bfr new_net_3230_bfr_before (
		.din(new_net_3230),
		.dout(new_net_3229)
	);

	bfr new_net_3231_bfr_before (
		.din(new_net_3231),
		.dout(new_net_3230)
	);

	bfr new_net_3232_bfr_before (
		.din(new_net_3232),
		.dout(new_net_3231)
	);

	bfr new_net_3233_bfr_before (
		.din(new_net_3233),
		.dout(new_net_3232)
	);

	bfr new_net_3234_bfr_before (
		.din(new_net_3234),
		.dout(new_net_3233)
	);

	bfr new_net_3235_bfr_before (
		.din(new_net_3235),
		.dout(new_net_3234)
	);

	bfr new_net_3236_bfr_before (
		.din(new_net_3236),
		.dout(new_net_3235)
	);

	bfr new_net_3237_bfr_before (
		.din(new_net_3237),
		.dout(new_net_3236)
	);

	bfr new_net_3238_bfr_before (
		.din(new_net_3238),
		.dout(new_net_3237)
	);

	bfr new_net_3239_bfr_before (
		.din(new_net_3239),
		.dout(new_net_3238)
	);

	bfr new_net_3240_bfr_before (
		.din(new_net_3240),
		.dout(new_net_3239)
	);

	bfr new_net_3241_bfr_before (
		.din(new_net_3241),
		.dout(new_net_3240)
	);

	bfr new_net_3242_bfr_before (
		.din(new_net_3242),
		.dout(new_net_3241)
	);

	bfr new_net_3243_bfr_before (
		.din(new_net_3243),
		.dout(new_net_3242)
	);

	bfr new_net_3244_bfr_before (
		.din(new_net_3244),
		.dout(new_net_3243)
	);

	bfr new_net_3245_bfr_before (
		.din(new_net_3245),
		.dout(new_net_3244)
	);

	bfr new_net_3246_bfr_before (
		.din(new_net_3246),
		.dout(new_net_3245)
	);

	bfr new_net_3247_bfr_before (
		.din(new_net_3247),
		.dout(new_net_3246)
	);

	bfr new_net_3248_bfr_before (
		.din(new_net_3248),
		.dout(new_net_3247)
	);

	bfr new_net_3249_bfr_before (
		.din(new_net_3249),
		.dout(new_net_3248)
	);

	bfr new_net_3250_bfr_before (
		.din(new_net_3250),
		.dout(new_net_3249)
	);

	bfr new_net_3251_bfr_before (
		.din(new_net_3251),
		.dout(new_net_3250)
	);

	bfr new_net_3252_bfr_before (
		.din(new_net_3252),
		.dout(new_net_3251)
	);

	spl4L new_net_2051_v_fanout (
		.a(new_net_2051),
		.b(new_net_1166),
		.c(new_net_3252),
		.d(new_net_1167),
		.e(new_net_1168)
	);

	bfr new_net_3253_bfr_before (
		.din(new_net_3253),
		.dout(new_net_1213)
	);

	bfr new_net_3254_bfr_before (
		.din(new_net_3254),
		.dout(new_net_1732)
	);

	bfr new_net_3255_bfr_before (
		.din(new_net_3255),
		.dout(new_net_3254)
	);

	spl3L new_net_1731_v_fanout (
		.a(new_net_1731),
		.b(new_net_1215),
		.c(new_net_3253),
		.d(new_net_3255)
	);

	spl2 _0641__v_fanout (
		.a(_0641_),
		.b(new_net_818),
		.c(new_net_819)
	);

	spl2 new_net_2050_v_fanout (
		.a(new_net_2050),
		.b(new_net_1164),
		.c(new_net_1165)
	);

	bfr new_net_3256_bfr_before (
		.din(new_net_3256),
		.dout(new_net_1036)
	);

	bfr new_net_3257_bfr_before (
		.din(new_net_3257),
		.dout(new_net_3256)
	);

	bfr new_net_3258_bfr_before (
		.din(new_net_3258),
		.dout(new_net_3257)
	);

	bfr new_net_3259_bfr_before (
		.din(new_net_3259),
		.dout(new_net_3258)
	);

	bfr new_net_3260_bfr_before (
		.din(new_net_3260),
		.dout(new_net_3259)
	);

	bfr new_net_3261_bfr_before (
		.din(new_net_3261),
		.dout(new_net_3260)
	);

	bfr new_net_3262_bfr_before (
		.din(new_net_3262),
		.dout(new_net_3261)
	);

	bfr new_net_3263_bfr_before (
		.din(new_net_3263),
		.dout(new_net_3262)
	);

	bfr new_net_3264_bfr_before (
		.din(new_net_3264),
		.dout(new_net_3263)
	);

	bfr new_net_3265_bfr_before (
		.din(new_net_3265),
		.dout(new_net_3264)
	);

	bfr new_net_3266_bfr_before (
		.din(new_net_3266),
		.dout(new_net_3265)
	);

	bfr new_net_3267_bfr_before (
		.din(new_net_3267),
		.dout(new_net_3266)
	);

	spl3L _0969__v_fanout (
		.a(_0969_),
		.b(new_net_1035),
		.c(new_net_3267),
		.d(new_net_1037)
	);

	bfr new_net_3268_bfr_before (
		.din(new_net_3268),
		.dout(new_net_2025)
	);

	spl2 new_net_2024_v_fanout (
		.a(new_net_2024),
		.b(new_net_1586),
		.c(new_net_3268)
	);

	bfr new_net_3269_bfr_before (
		.din(new_net_3269),
		.dout(new_net_1784)
	);

	spl2 new_net_1783_v_fanout (
		.a(new_net_1783),
		.b(new_net_3269),
		.c(new_net_54)
	);

	spl2 _0073__v_fanout (
		.a(_0073_),
		.b(new_net_489),
		.c(new_net_490)
	);

	spl2 _1244__v_fanout (
		.a(_1244_),
		.b(new_net_1331),
		.c(new_net_1332)
	);

	spl2 _0156__v_fanout (
		.a(_0156_),
		.b(new_net_921),
		.c(new_net_922)
	);

	spl2 new_net_2037_v_fanout (
		.a(new_net_2037),
		.b(new_net_1328),
		.c(new_net_1327)
	);

	bfr new_net_3270_bfr_before (
		.din(new_net_3270),
		.dout(new_net_2055)
	);

	bfr new_net_3271_bfr_before (
		.din(new_net_3271),
		.dout(new_net_3270)
	);

	bfr new_net_3272_bfr_before (
		.din(new_net_3272),
		.dout(new_net_3271)
	);

	bfr new_net_3273_bfr_before (
		.din(new_net_3273),
		.dout(new_net_3272)
	);

	bfr new_net_3274_bfr_before (
		.din(new_net_3274),
		.dout(new_net_3273)
	);

	bfr new_net_3275_bfr_before (
		.din(new_net_3275),
		.dout(new_net_3274)
	);

	bfr new_net_3276_bfr_before (
		.din(new_net_3276),
		.dout(new_net_3275)
	);

	spl4L _0684__v_fanout (
		.a(_0684_),
		.b(new_net_1448),
		.c(new_net_1449),
		.d(new_net_1452),
		.e(new_net_3276)
	);

	bfr new_net_3277_bfr_before (
		.din(new_net_3277),
		.dout(new_net_2049)
	);

	bfr new_net_3278_bfr_before (
		.din(new_net_3278),
		.dout(new_net_3277)
	);

	bfr new_net_3279_bfr_before (
		.din(new_net_3279),
		.dout(new_net_3278)
	);

	bfr new_net_3280_bfr_before (
		.din(new_net_3280),
		.dout(new_net_3279)
	);

	bfr new_net_3281_bfr_before (
		.din(new_net_3281),
		.dout(new_net_3280)
	);

	bfr new_net_3282_bfr_before (
		.din(new_net_3282),
		.dout(new_net_3281)
	);

	bfr new_net_3283_bfr_before (
		.din(new_net_3283),
		.dout(new_net_3282)
	);

	bfr new_net_3284_bfr_before (
		.din(new_net_3284),
		.dout(new_net_3283)
	);

	bfr new_net_3285_bfr_before (
		.din(new_net_3285),
		.dout(new_net_3284)
	);

	bfr new_net_3286_bfr_before (
		.din(new_net_3286),
		.dout(new_net_3285)
	);

	bfr new_net_3287_bfr_before (
		.din(new_net_3287),
		.dout(new_net_3286)
	);

	spl3L _0873__v_fanout (
		.a(_0873_),
		.b(new_net_228),
		.c(new_net_230),
		.d(new_net_3287)
	);

	spl2 _0046__v_fanout (
		.a(_0046_),
		.b(new_net_495),
		.c(new_net_496)
	);

	spl2 _1158__v_fanout (
		.a(_1158_),
		.b(new_net_831),
		.c(new_net_832)
	);

	spl2 new_net_1_v_fanout (
		.a(new_net_1),
		.b(new_net_2051),
		.c(new_net_2050)
	);

	bfr new_net_3288_bfr_before (
		.din(new_net_3288),
		.dout(new_net_2053)
	);

	bfr new_net_3289_bfr_before (
		.din(new_net_3289),
		.dout(new_net_3288)
	);

	spl3L _0936__v_fanout (
		.a(_0936_),
		.b(new_net_1447),
		.c(new_net_1445),
		.d(new_net_3289)
	);

	spl2 new_net_2043_v_fanout (
		.a(new_net_2043),
		.b(new_net_721),
		.c(new_net_2044)
	);

	spl2 _0618__v_fanout (
		.a(_0618_),
		.b(new_net_191),
		.c(new_net_192)
	);

	spl2 _0067__v_fanout (
		.a(_0067_),
		.b(new_net_74),
		.c(new_net_75)
	);

	bfr new_net_3290_bfr_after (
		.din(_1182_),
		.dout(new_net_3290)
	);

	bfr new_net_3291_bfr_after (
		.din(new_net_3290),
		.dout(new_net_3291)
	);

	bfr new_net_3292_bfr_after (
		.din(new_net_3291),
		.dout(new_net_3292)
	);

	spl2 _1182__v_fanout (
		.a(new_net_3292),
		.b(new_net_1097),
		.c(new_net_1098)
	);

	spl2 _1212__v_fanout (
		.a(_1212_),
		.b(new_net_289),
		.c(new_net_290)
	);

	spl2 _0130__v_fanout (
		.a(_0130_),
		.b(new_net_493),
		.c(new_net_494)
	);

	spl2 _1146__v_fanout (
		.a(_1146_),
		.b(new_net_1456),
		.c(new_net_1457)
	);

	bfr new_net_3293_bfr_before (
		.din(new_net_3293),
		.dout(new_net_406)
	);

	bfr new_net_3294_bfr_before (
		.din(new_net_3294),
		.dout(new_net_3293)
	);

	bfr new_net_3295_bfr_before (
		.din(new_net_3295),
		.dout(new_net_3294)
	);

	bfr new_net_3296_bfr_before (
		.din(new_net_3296),
		.dout(new_net_3295)
	);

	bfr new_net_3297_bfr_before (
		.din(new_net_3297),
		.dout(new_net_3296)
	);

	bfr new_net_3298_bfr_before (
		.din(new_net_3298),
		.dout(new_net_3297)
	);

	bfr new_net_3299_bfr_before (
		.din(new_net_3299),
		.dout(new_net_3298)
	);

	bfr new_net_3300_bfr_before (
		.din(new_net_3300),
		.dout(new_net_3299)
	);

	bfr new_net_3301_bfr_before (
		.din(new_net_3301),
		.dout(new_net_3300)
	);

	bfr new_net_3302_bfr_before (
		.din(new_net_3302),
		.dout(new_net_3301)
	);

	bfr new_net_3303_bfr_before (
		.din(new_net_3303),
		.dout(new_net_3302)
	);

	bfr new_net_3304_bfr_before (
		.din(new_net_3304),
		.dout(new_net_3303)
	);

	bfr new_net_3305_bfr_before (
		.din(new_net_3305),
		.dout(new_net_3304)
	);

	bfr new_net_3306_bfr_before (
		.din(new_net_3306),
		.dout(new_net_3305)
	);

	bfr new_net_3307_bfr_before (
		.din(new_net_3307),
		.dout(new_net_3306)
	);

	bfr new_net_3308_bfr_before (
		.din(new_net_3308),
		.dout(new_net_3307)
	);

	spl2 new_net_2039_v_fanout (
		.a(new_net_2039),
		.b(new_net_407),
		.c(new_net_3308)
	);

	bfr new_net_3309_bfr_before (
		.din(new_net_3309),
		.dout(new_net_211)
	);

	bfr new_net_3310_bfr_before (
		.din(new_net_3310),
		.dout(new_net_3309)
	);

	bfr new_net_3311_bfr_before (
		.din(new_net_3311),
		.dout(new_net_3310)
	);

	bfr new_net_3312_bfr_before (
		.din(new_net_3312),
		.dout(new_net_3311)
	);

	bfr new_net_3313_bfr_before (
		.din(new_net_3313),
		.dout(new_net_3312)
	);

	bfr new_net_3314_bfr_before (
		.din(new_net_3314),
		.dout(new_net_3313)
	);

	spl2 new_net_2032_v_fanout (
		.a(new_net_2032),
		.b(new_net_210),
		.c(new_net_3314)
	);

	bfr new_net_3315_bfr_before (
		.din(new_net_3315),
		.dout(new_net_2052)
	);

	bfr new_net_3316_bfr_before (
		.din(new_net_3316),
		.dout(new_net_3315)
	);

	bfr new_net_3317_bfr_before (
		.din(new_net_3317),
		.dout(new_net_3316)
	);

	bfr new_net_3318_bfr_before (
		.din(new_net_3318),
		.dout(new_net_3317)
	);

	bfr new_net_3319_bfr_before (
		.din(new_net_3319),
		.dout(new_net_3318)
	);

	bfr new_net_3320_bfr_before (
		.din(new_net_3320),
		.dout(new_net_3319)
	);

	bfr new_net_3321_bfr_before (
		.din(new_net_3321),
		.dout(new_net_3320)
	);

	bfr new_net_3322_bfr_before (
		.din(new_net_3322),
		.dout(new_net_3321)
	);

	bfr new_net_3323_bfr_before (
		.din(new_net_3323),
		.dout(new_net_3322)
	);

	bfr new_net_3324_bfr_before (
		.din(new_net_3324),
		.dout(new_net_3323)
	);

	bfr new_net_3325_bfr_before (
		.din(new_net_3325),
		.dout(new_net_3324)
	);

	bfr new_net_3326_bfr_before (
		.din(new_net_3326),
		.dout(new_net_3325)
	);

	bfr new_net_3327_bfr_before (
		.din(new_net_3327),
		.dout(new_net_3326)
	);

	bfr new_net_3328_bfr_before (
		.din(new_net_3328),
		.dout(new_net_3327)
	);

	spl2 _0871__v_fanout (
		.a(_0871_),
		.b(new_net_205),
		.c(new_net_3328)
	);

	bfr new_net_3329_bfr_after (
		.din(_1013_),
		.dout(new_net_3329)
	);

	bfr new_net_3330_bfr_before (
		.din(new_net_3330),
		.dout(new_net_507)
	);

	bfr new_net_3331_bfr_before (
		.din(new_net_3331),
		.dout(new_net_3330)
	);

	bfr new_net_3332_bfr_before (
		.din(new_net_3332),
		.dout(new_net_3331)
	);

	bfr new_net_3333_bfr_before (
		.din(new_net_3333),
		.dout(new_net_3332)
	);

	bfr new_net_3334_bfr_before (
		.din(new_net_3334),
		.dout(new_net_3333)
	);

	bfr new_net_3335_bfr_before (
		.din(new_net_3335),
		.dout(new_net_3334)
	);

	bfr new_net_3336_bfr_before (
		.din(new_net_3336),
		.dout(new_net_3335)
	);

	bfr new_net_3337_bfr_before (
		.din(new_net_3337),
		.dout(new_net_3336)
	);

	bfr new_net_3338_bfr_before (
		.din(new_net_3338),
		.dout(new_net_3337)
	);

	bfr new_net_3339_bfr_before (
		.din(new_net_3339),
		.dout(new_net_3338)
	);

	bfr new_net_3340_bfr_before (
		.din(new_net_3340),
		.dout(new_net_3339)
	);

	bfr new_net_3341_bfr_before (
		.din(new_net_3341),
		.dout(new_net_3340)
	);

	bfr new_net_3342_bfr_before (
		.din(new_net_3342),
		.dout(new_net_3341)
	);

	bfr new_net_3343_bfr_before (
		.din(new_net_3343),
		.dout(new_net_3342)
	);

	bfr new_net_3344_bfr_before (
		.din(new_net_3344),
		.dout(new_net_3343)
	);

	bfr new_net_3345_bfr_before (
		.din(new_net_3345),
		.dout(new_net_3344)
	);

	spl2 _1013__v_fanout (
		.a(new_net_3329),
		.b(new_net_3345),
		.c(new_net_508)
	);

	bfr new_net_3346_bfr_before (
		.din(new_net_3346),
		.dout(new_net_66)
	);

	bfr new_net_3347_bfr_before (
		.din(new_net_3347),
		.dout(new_net_3346)
	);

	bfr new_net_3348_bfr_before (
		.din(new_net_3348),
		.dout(new_net_3347)
	);

	bfr new_net_3349_bfr_before (
		.din(new_net_3349),
		.dout(new_net_3348)
	);

	bfr new_net_3350_bfr_before (
		.din(new_net_3350),
		.dout(new_net_3349)
	);

	bfr new_net_3351_bfr_before (
		.din(new_net_3351),
		.dout(new_net_3350)
	);

	spl3L _0738__v_fanout (
		.a(_0738_),
		.b(new_net_65),
		.c(new_net_67),
		.d(new_net_3351)
	);

	spl2 new_net_2033_v_fanout (
		.a(new_net_2033),
		.b(new_net_212),
		.c(new_net_215)
	);

	spl2 _0207__v_fanout (
		.a(_0207_),
		.b(new_net_1681),
		.c(new_net_1682)
	);

	bfr new_net_3352_bfr_before (
		.din(new_net_3352),
		.dout(new_net_2045)
	);

	bfr new_net_3353_bfr_before (
		.din(new_net_3353),
		.dout(new_net_3352)
	);

	bfr new_net_3354_bfr_before (
		.din(new_net_3354),
		.dout(new_net_3353)
	);

	spl3L _0754__v_fanout (
		.a(_0754_),
		.b(new_net_1649),
		.c(new_net_1652),
		.d(new_net_3354)
	);

	spl2 _0171__v_fanout (
		.a(_0171_),
		.b(new_net_1316),
		.c(new_net_1317)
	);

	bfr new_net_3355_bfr_before (
		.din(new_net_3355),
		.dout(new_net_288)
	);

	spl2 _0071__v_fanout (
		.a(_0071_),
		.b(new_net_287),
		.c(new_net_3355)
	);

	spl3L new_net_2034_v_fanout (
		.a(new_net_2034),
		.b(new_net_2032),
		.c(new_net_213),
		.d(new_net_214)
	);

	bfr new_net_3356_bfr_before (
		.din(new_net_3356),
		.dout(new_net_1295)
	);

	bfr new_net_3357_bfr_before (
		.din(new_net_3357),
		.dout(new_net_3356)
	);

	bfr new_net_3358_bfr_before (
		.din(new_net_3358),
		.dout(new_net_3357)
	);

	bfr new_net_3359_bfr_before (
		.din(new_net_3359),
		.dout(new_net_3358)
	);

	bfr new_net_3360_bfr_before (
		.din(new_net_3360),
		.dout(new_net_3359)
	);

	spl2 _0954__v_fanout (
		.a(_0954_),
		.b(new_net_1294),
		.c(new_net_3360)
	);

	bfr new_net_3361_bfr_before (
		.din(new_net_3361),
		.dout(new_net_2040)
	);

	spl3L _0964__v_fanout (
		.a(_0964_),
		.b(new_net_393),
		.c(new_net_391),
		.d(new_net_3361)
	);

	spl2 _0162__v_fanout (
		.a(_0162_),
		.b(new_net_396),
		.c(new_net_397)
	);

	bfr new_net_3362_bfr_before (
		.din(new_net_3362),
		.dout(new_net_455)
	);

	bfr new_net_3363_bfr_before (
		.din(new_net_3363),
		.dout(new_net_3362)
	);

	bfr new_net_3364_bfr_before (
		.din(new_net_3364),
		.dout(new_net_3363)
	);

	bfr new_net_3365_bfr_before (
		.din(new_net_3365),
		.dout(new_net_3364)
	);

	bfr new_net_3366_bfr_before (
		.din(new_net_3366),
		.dout(new_net_3365)
	);

	bfr new_net_3367_bfr_before (
		.din(new_net_3367),
		.dout(new_net_3366)
	);

	bfr new_net_3368_bfr_before (
		.din(new_net_3368),
		.dout(new_net_3367)
	);

	bfr new_net_3369_bfr_before (
		.din(new_net_3369),
		.dout(new_net_3368)
	);

	bfr new_net_3370_bfr_before (
		.din(new_net_3370),
		.dout(new_net_3369)
	);

	bfr new_net_3371_bfr_before (
		.din(new_net_3371),
		.dout(new_net_3370)
	);

	bfr new_net_3372_bfr_before (
		.din(new_net_3372),
		.dout(new_net_3371)
	);

	bfr new_net_3373_bfr_before (
		.din(new_net_3373),
		.dout(new_net_3372)
	);

	bfr new_net_3374_bfr_before (
		.din(new_net_3374),
		.dout(new_net_3373)
	);

	bfr new_net_3375_bfr_before (
		.din(new_net_3375),
		.dout(new_net_3374)
	);

	spl3L new_net_2021_v_fanout (
		.a(new_net_2021),
		.b(new_net_3375),
		.c(new_net_453),
		.d(new_net_454)
	);

	spl3L _0640__v_fanout (
		.a(_0640_),
		.b(new_net_720),
		.c(new_net_724),
		.d(new_net_2043)
	);

	bfr new_net_3376_bfr_before (
		.din(new_net_3376),
		.dout(new_net_2042)
	);

	bfr new_net_3377_bfr_before (
		.din(new_net_3377),
		.dout(new_net_3376)
	);

	bfr new_net_3378_bfr_before (
		.din(new_net_3378),
		.dout(new_net_3377)
	);

	bfr new_net_3379_bfr_before (
		.din(new_net_3379),
		.dout(new_net_3378)
	);

	bfr new_net_3380_bfr_before (
		.din(new_net_3380),
		.dout(new_net_3379)
	);

	bfr new_net_3381_bfr_before (
		.din(new_net_3381),
		.dout(new_net_3380)
	);

	bfr new_net_3382_bfr_before (
		.din(new_net_3382),
		.dout(new_net_3381)
	);

	bfr new_net_3383_bfr_before (
		.din(new_net_3383),
		.dout(new_net_3382)
	);

	spl4L _0760__v_fanout (
		.a(_0760_),
		.b(new_net_540),
		.c(new_net_544),
		.d(new_net_542),
		.e(new_net_3383)
	);

	bfr new_net_3384_bfr_after (
		.din(_0766_),
		.dout(new_net_3384)
	);

	spl2 _0766__v_fanout (
		.a(new_net_3384),
		.b(new_net_1099),
		.c(new_net_1100)
	);

	spl2 _0177__v_fanout (
		.a(_0177_),
		.b(new_net_193),
		.c(new_net_194)
	);

	spl2 _0965__v_fanout (
		.a(_0965_),
		.b(new_net_405),
		.c(new_net_2039)
	);

	spl2 _0192__v_fanout (
		.a(_0192_),
		.b(new_net_180),
		.c(new_net_181)
	);

	bfr new_net_3385_bfr_before (
		.din(new_net_3385),
		.dout(new_net_2038)
	);

	bfr new_net_3386_bfr_before (
		.din(new_net_3386),
		.dout(new_net_3385)
	);

	bfr new_net_3387_bfr_before (
		.din(new_net_3387),
		.dout(new_net_3386)
	);

	bfr new_net_3388_bfr_before (
		.din(new_net_3388),
		.dout(new_net_3387)
	);

	spl3L _1238__v_fanout (
		.a(_1238_),
		.b(new_net_170),
		.c(new_net_168),
		.d(new_net_3388)
	);

	bfr new_net_3389_bfr_before (
		.din(new_net_3389),
		.dout(new_net_719)
	);

	bfr new_net_3390_bfr_before (
		.din(new_net_3390),
		.dout(new_net_3389)
	);

	spl2 _0599__v_fanout (
		.a(_0599_),
		.b(new_net_718),
		.c(new_net_3390)
	);

	bfr new_net_3391_bfr_before (
		.din(new_net_3391),
		.dout(new_net_2047)
	);

	bfr new_net_3392_bfr_before (
		.din(new_net_3392),
		.dout(new_net_3391)
	);

	bfr new_net_3393_bfr_before (
		.din(new_net_3393),
		.dout(new_net_3392)
	);

	bfr new_net_3394_bfr_before (
		.din(new_net_3394),
		.dout(new_net_3393)
	);

	bfr new_net_3395_bfr_before (
		.din(new_net_3395),
		.dout(new_net_3394)
	);

	bfr new_net_3396_bfr_before (
		.din(new_net_3396),
		.dout(new_net_3395)
	);

	bfr new_net_3397_bfr_before (
		.din(new_net_3397),
		.dout(new_net_3396)
	);

	bfr new_net_3398_bfr_before (
		.din(new_net_3398),
		.dout(new_net_3397)
	);

	bfr new_net_3399_bfr_before (
		.din(new_net_3399),
		.dout(new_net_3398)
	);

	bfr new_net_3400_bfr_before (
		.din(new_net_3400),
		.dout(new_net_3399)
	);

	bfr new_net_3401_bfr_before (
		.din(new_net_3401),
		.dout(new_net_3400)
	);

	bfr new_net_3402_bfr_before (
		.din(new_net_3402),
		.dout(new_net_3401)
	);

	bfr new_net_3403_bfr_before (
		.din(new_net_3403),
		.dout(new_net_3402)
	);

	spl2 _0968__v_fanout (
		.a(_0968_),
		.b(new_net_472),
		.c(new_net_3403)
	);

	bfr new_net_3404_bfr_before (
		.din(new_net_3404),
		.dout(new_net_2048)
	);

	bfr new_net_3405_bfr_before (
		.din(new_net_3405),
		.dout(new_net_3404)
	);

	bfr new_net_3406_bfr_before (
		.din(new_net_3406),
		.dout(new_net_3405)
	);

	bfr new_net_3407_bfr_before (
		.din(new_net_3407),
		.dout(new_net_3406)
	);

	spl2 _0669__v_fanout (
		.a(_0669_),
		.b(new_net_1180),
		.c(new_net_3407)
	);

	bfr new_net_3408_bfr_after (
		.din(_0076_),
		.dout(new_net_3408)
	);

	bfr new_net_3409_bfr_after (
		.din(new_net_3408),
		.dout(new_net_3409)
	);

	spl2 _0076__v_fanout (
		.a(new_net_3409),
		.b(new_net_739),
		.c(new_net_740)
	);

	bfr new_net_3410_bfr_after (
		.din(_0662_),
		.dout(new_net_3410)
	);

	bfr new_net_3411_bfr_after (
		.din(new_net_3410),
		.dout(new_net_3411)
	);

	bfr new_net_3412_bfr_before (
		.din(new_net_3412),
		.dout(new_net_2035)
	);

	bfr new_net_3413_bfr_before (
		.din(new_net_3413),
		.dout(new_net_3412)
	);

	bfr new_net_3414_bfr_before (
		.din(new_net_3414),
		.dout(new_net_3413)
	);

	spl3L _0662__v_fanout (
		.a(new_net_3411),
		.b(new_net_974),
		.c(new_net_976),
		.d(new_net_3414)
	);

	bfr new_net_3415_bfr_before (
		.din(new_net_3415),
		.dout(new_net_1713)
	);

	bfr new_net_3416_bfr_before (
		.din(new_net_3416),
		.dout(new_net_3415)
	);

	spl4L _0615__v_fanout (
		.a(_0615_),
		.b(new_net_3416),
		.c(new_net_1712),
		.d(new_net_1714),
		.e(new_net_1711)
	);

	bfr new_net_3417_bfr_before (
		.din(new_net_3417),
		.dout(new_net_2037)
	);

	bfr new_net_3418_bfr_before (
		.din(new_net_3418),
		.dout(new_net_3417)
	);

	spl2 _0424__v_fanout (
		.a(_0424_),
		.b(new_net_1326),
		.c(new_net_3418)
	);

	bfr new_net_3419_bfr_before (
		.din(new_net_3419),
		.dout(new_net_330)
	);

	bfr new_net_3420_bfr_before (
		.din(new_net_3420),
		.dout(new_net_3419)
	);

	spl2 _0584__v_fanout (
		.a(_0584_),
		.b(new_net_329),
		.c(new_net_3420)
	);

	bfr new_net_3421_bfr_before (
		.din(new_net_3421),
		.dout(new_net_1433)
	);

	bfr new_net_3422_bfr_before (
		.din(new_net_3422),
		.dout(new_net_3421)
	);

	bfr new_net_3423_bfr_before (
		.din(new_net_3423),
		.dout(new_net_3422)
	);

	bfr new_net_3424_bfr_before (
		.din(new_net_3424),
		.dout(new_net_3423)
	);

	spl4L _0613__v_fanout (
		.a(_0613_),
		.b(new_net_3424),
		.c(new_net_1432),
		.d(new_net_1434),
		.e(new_net_1431)
	);

	bfr new_net_3425_bfr_before (
		.din(new_net_3425),
		.dout(new_net_324)
	);

	spl3L _0863__v_fanout (
		.a(_0863_),
		.b(new_net_3425),
		.c(new_net_326),
		.d(new_net_325)
	);

	bfr new_net_3426_bfr_before (
		.din(new_net_3426),
		.dout(new_net_560)
	);

	bfr new_net_3427_bfr_before (
		.din(new_net_3427),
		.dout(new_net_3426)
	);

	spl2 new_net_2027_v_fanout (
		.a(new_net_2027),
		.b(new_net_3427),
		.c(new_net_559)
	);

	bfr new_net_3428_bfr_after (
		.din(_0198_),
		.dout(new_net_3428)
	);

	bfr new_net_3429_bfr_after (
		.din(new_net_3428),
		.dout(new_net_3429)
	);

	bfr new_net_3430_bfr_after (
		.din(new_net_3429),
		.dout(new_net_3430)
	);

	bfr new_net_3431_bfr_after (
		.din(new_net_3430),
		.dout(new_net_3431)
	);

	spl2 _0198__v_fanout (
		.a(new_net_3431),
		.b(new_net_189),
		.c(new_net_190)
	);

	bfr new_net_3432_bfr_after (
		.din(_0609_),
		.dout(new_net_3432)
	);

	spl3L _0609__v_fanout (
		.a(new_net_3432),
		.b(new_net_104),
		.c(new_net_106),
		.d(new_net_105)
	);

	bfr new_net_3433_bfr_after (
		.din(_0204_),
		.dout(new_net_3433)
	);

	spl2 _0204__v_fanout (
		.a(new_net_3433),
		.b(new_net_291),
		.c(new_net_292)
	);

	bfr new_net_3434_bfr_after (
		.din(_0141_),
		.dout(new_net_3434)
	);

	bfr new_net_3435_bfr_after (
		.din(new_net_3434),
		.dout(new_net_3435)
	);

	bfr new_net_3436_bfr_after (
		.din(new_net_3435),
		.dout(new_net_3436)
	);

	spl2 _0141__v_fanout (
		.a(new_net_3436),
		.b(new_net_1460),
		.c(new_net_1461)
	);

	bfr new_net_3437_bfr_before (
		.din(new_net_3437),
		.dout(new_net_850)
	);

	bfr new_net_3438_bfr_before (
		.din(new_net_3438),
		.dout(new_net_3437)
	);

	bfr new_net_3439_bfr_before (
		.din(new_net_3439),
		.dout(new_net_3438)
	);

	bfr new_net_3440_bfr_before (
		.din(new_net_3440),
		.dout(new_net_3439)
	);

	bfr new_net_3441_bfr_before (
		.din(new_net_3441),
		.dout(new_net_3440)
	);

	bfr new_net_3442_bfr_before (
		.din(new_net_3442),
		.dout(new_net_3441)
	);

	bfr new_net_3443_bfr_before (
		.din(new_net_3443),
		.dout(new_net_3442)
	);

	spl2 _0935__v_fanout (
		.a(_0935_),
		.b(new_net_849),
		.c(new_net_3443)
	);

	bfr new_net_3444_bfr_before (
		.din(new_net_3444),
		.dout(new_net_1411)
	);

	bfr new_net_3445_bfr_before (
		.din(new_net_3445),
		.dout(new_net_3444)
	);

	bfr new_net_3446_bfr_before (
		.din(new_net_3446),
		.dout(new_net_3445)
	);

	bfr new_net_3447_bfr_before (
		.din(new_net_3447),
		.dout(new_net_3446)
	);

	bfr new_net_3448_bfr_before (
		.din(new_net_3448),
		.dout(new_net_3447)
	);

	bfr new_net_3449_bfr_before (
		.din(new_net_3449),
		.dout(new_net_3448)
	);

	bfr new_net_3450_bfr_before (
		.din(new_net_3450),
		.dout(new_net_3449)
	);

	bfr new_net_3451_bfr_before (
		.din(new_net_3451),
		.dout(new_net_3450)
	);

	bfr new_net_3452_bfr_before (
		.din(new_net_3452),
		.dout(new_net_3451)
	);

	bfr new_net_3453_bfr_before (
		.din(new_net_3453),
		.dout(new_net_3452)
	);

	bfr new_net_3454_bfr_before (
		.din(new_net_3454),
		.dout(new_net_3453)
	);

	spl2 _0682__v_fanout (
		.a(_0682_),
		.b(new_net_1410),
		.c(new_net_3454)
	);

	spl4L new_net_2001_v_fanout (
		.a(new_net_2001),
		.b(new_net_616),
		.c(new_net_619),
		.d(new_net_629),
		.e(new_net_625)
	);

	bfr new_net_3455_bfr_after (
		.din(_0189_),
		.dout(new_net_3455)
	);

	spl2 _0189__v_fanout (
		.a(new_net_3455),
		.b(new_net_1699),
		.c(new_net_1700)
	);

	bfr new_net_3456_bfr_after (
		.din(_0118_),
		.dout(new_net_3456)
	);

	bfr new_net_3457_bfr_after (
		.din(new_net_3456),
		.dout(new_net_3457)
	);

	spl2 _0118__v_fanout (
		.a(new_net_3457),
		.b(new_net_255),
		.c(new_net_256)
	);

	bfr new_net_3458_bfr_before (
		.din(new_net_3458),
		.dout(new_net_1200)
	);

	bfr new_net_3459_bfr_before (
		.din(new_net_3459),
		.dout(new_net_3458)
	);

	bfr new_net_3460_bfr_before (
		.din(new_net_3460),
		.dout(new_net_3459)
	);

	bfr new_net_3461_bfr_before (
		.din(new_net_3461),
		.dout(new_net_3460)
	);

	bfr new_net_3462_bfr_before (
		.din(new_net_3462),
		.dout(new_net_3461)
	);

	bfr new_net_3463_bfr_before (
		.din(new_net_3463),
		.dout(new_net_3462)
	);

	bfr new_net_3464_bfr_before (
		.din(new_net_3464),
		.dout(new_net_3463)
	);

	bfr new_net_3465_bfr_before (
		.din(new_net_3465),
		.dout(new_net_3464)
	);

	bfr new_net_3466_bfr_before (
		.din(new_net_3466),
		.dout(new_net_3465)
	);

	bfr new_net_3467_bfr_before (
		.din(new_net_3467),
		.dout(new_net_3466)
	);

	bfr new_net_3468_bfr_before (
		.din(new_net_3468),
		.dout(new_net_3467)
	);

	bfr new_net_3469_bfr_before (
		.din(new_net_3469),
		.dout(new_net_3468)
	);

	bfr new_net_3470_bfr_before (
		.din(new_net_3470),
		.dout(new_net_3469)
	);

	bfr new_net_3471_bfr_before (
		.din(new_net_3471),
		.dout(new_net_3470)
	);

	spl3L new_net_2031_v_fanout (
		.a(new_net_2031),
		.b(new_net_1198),
		.c(new_net_1202),
		.d(new_net_3471)
	);

	spl4L new_net_2000_v_fanout (
		.a(new_net_2000),
		.b(new_net_623),
		.c(new_net_615),
		.d(new_net_612),
		.e(new_net_610)
	);

	bfr new_net_3472_bfr_before (
		.din(new_net_3472),
		.dout(new_net_1999)
	);

	bfr new_net_3473_bfr_before (
		.din(new_net_3473),
		.dout(new_net_3472)
	);

	bfr new_net_3474_bfr_before (
		.din(new_net_3474),
		.dout(new_net_3473)
	);

	bfr new_net_3475_bfr_before (
		.din(new_net_3475),
		.dout(new_net_3474)
	);

	bfr new_net_3476_bfr_before (
		.din(new_net_3476),
		.dout(new_net_3475)
	);

	bfr new_net_3477_bfr_before (
		.din(new_net_3477),
		.dout(new_net_3476)
	);

	bfr new_net_3478_bfr_before (
		.din(new_net_3478),
		.dout(new_net_3477)
	);

	bfr new_net_3479_bfr_before (
		.din(new_net_3479),
		.dout(new_net_3478)
	);

	spl4L new_net_1998_v_fanout (
		.a(new_net_1998),
		.b(new_net_3479),
		.c(new_net_617),
		.d(new_net_618),
		.e(new_net_628)
	);

	bfr new_net_3480_bfr_before (
		.din(new_net_3480),
		.dout(new_net_783)
	);

	bfr new_net_3481_bfr_before (
		.din(new_net_3481),
		.dout(new_net_3480)
	);

	bfr new_net_3482_bfr_before (
		.din(new_net_3482),
		.dout(new_net_3481)
	);

	bfr new_net_3483_bfr_before (
		.din(new_net_3483),
		.dout(new_net_3482)
	);

	bfr new_net_3484_bfr_before (
		.din(new_net_3484),
		.dout(new_net_3483)
	);

	bfr new_net_3485_bfr_before (
		.din(new_net_3485),
		.dout(new_net_3484)
	);

	bfr new_net_3486_bfr_before (
		.din(new_net_3486),
		.dout(new_net_3485)
	);

	bfr new_net_3487_bfr_before (
		.din(new_net_3487),
		.dout(new_net_3486)
	);

	bfr new_net_3488_bfr_before (
		.din(new_net_3488),
		.dout(new_net_3487)
	);

	bfr new_net_3489_bfr_before (
		.din(new_net_3489),
		.dout(new_net_3488)
	);

	bfr new_net_3490_bfr_before (
		.din(new_net_3490),
		.dout(new_net_3489)
	);

	bfr new_net_3491_bfr_before (
		.din(new_net_3491),
		.dout(new_net_3490)
	);

	bfr new_net_3492_bfr_before (
		.din(new_net_3492),
		.dout(new_net_3491)
	);

	bfr new_net_3493_bfr_before (
		.din(new_net_3493),
		.dout(new_net_3492)
	);

	spl4L new_net_2029_v_fanout (
		.a(new_net_2029),
		.b(new_net_782),
		.c(new_net_780),
		.d(new_net_3493),
		.e(new_net_779)
	);

	spl2 _0150__v_fanout (
		.a(_0150_),
		.b(new_net_829),
		.c(new_net_830)
	);

	bfr new_net_3494_bfr_before (
		.din(new_net_3494),
		.dout(new_net_1390)
	);

	bfr new_net_3495_bfr_before (
		.din(new_net_3495),
		.dout(new_net_3494)
	);

	bfr new_net_3496_bfr_before (
		.din(new_net_3496),
		.dout(new_net_3495)
	);

	bfr new_net_3497_bfr_before (
		.din(new_net_3497),
		.dout(new_net_3496)
	);

	bfr new_net_3498_bfr_before (
		.din(new_net_3498),
		.dout(new_net_3497)
	);

	bfr new_net_3499_bfr_before (
		.din(new_net_3499),
		.dout(new_net_3498)
	);

	bfr new_net_3500_bfr_before (
		.din(new_net_3500),
		.dout(new_net_3499)
	);

	bfr new_net_3501_bfr_before (
		.din(new_net_3501),
		.dout(new_net_3500)
	);

	spl2 _0932__v_fanout (
		.a(_0932_),
		.b(new_net_1389),
		.c(new_net_3501)
	);

	bfr new_net_3502_bfr_before (
		.din(new_net_3502),
		.dout(new_net_589)
	);

	bfr new_net_3503_bfr_before (
		.din(new_net_3503),
		.dout(new_net_3502)
	);

	bfr new_net_3504_bfr_before (
		.din(new_net_3504),
		.dout(new_net_3503)
	);

	spl2 new_net_1802_v_fanout (
		.a(new_net_1802),
		.b(new_net_3504),
		.c(new_net_592)
	);

	spl2 new_net_2030_v_fanout (
		.a(new_net_2030),
		.b(new_net_1199),
		.c(new_net_1201)
	);

	bfr new_net_3505_bfr_after (
		.din(_0673_),
		.dout(new_net_3505)
	);

	bfr new_net_3506_bfr_after (
		.din(new_net_3505),
		.dout(new_net_3506)
	);

	bfr new_net_3507_bfr_after (
		.din(new_net_3506),
		.dout(new_net_3507)
	);

	bfr new_net_3508_bfr_before (
		.din(new_net_3508),
		.dout(new_net_815)
	);

	bfr new_net_3509_bfr_before (
		.din(new_net_3509),
		.dout(new_net_3508)
	);

	bfr new_net_3510_bfr_before (
		.din(new_net_3510),
		.dout(new_net_3509)
	);

	bfr new_net_3511_bfr_before (
		.din(new_net_3511),
		.dout(new_net_3510)
	);

	bfr new_net_3512_bfr_before (
		.din(new_net_3512),
		.dout(new_net_3511)
	);

	spl2 _0673__v_fanout (
		.a(new_net_3507),
		.b(new_net_814),
		.c(new_net_3512)
	);

	bfr new_net_3513_bfr_before (
		.din(new_net_3513),
		.dout(new_net_1430)
	);

	bfr new_net_3514_bfr_before (
		.din(new_net_3514),
		.dout(new_net_3513)
	);

	bfr new_net_3515_bfr_before (
		.din(new_net_3515),
		.dout(new_net_3514)
	);

	bfr new_net_3516_bfr_before (
		.din(new_net_3516),
		.dout(new_net_3515)
	);

	bfr new_net_3517_bfr_before (
		.din(new_net_3517),
		.dout(new_net_3516)
	);

	bfr new_net_3518_bfr_before (
		.din(new_net_3518),
		.dout(new_net_3517)
	);

	bfr new_net_3519_bfr_before (
		.din(new_net_3519),
		.dout(new_net_3518)
	);

	bfr new_net_3520_bfr_before (
		.din(new_net_3520),
		.dout(new_net_3519)
	);

	bfr new_net_3521_bfr_before (
		.din(new_net_3521),
		.dout(new_net_3520)
	);

	bfr new_net_3522_bfr_before (
		.din(new_net_3522),
		.dout(new_net_3521)
	);

	spl2 _0683__v_fanout (
		.a(_0683_),
		.b(new_net_1429),
		.c(new_net_3522)
	);

	spl2 _0746__v_fanout (
		.a(_0746_),
		.b(new_net_2033),
		.c(new_net_2034)
	);

	bfr new_net_3523_bfr_before (
		.din(new_net_3523),
		.dout(new_net_60)
	);

	spl3L _0864__v_fanout (
		.a(_0864_),
		.b(new_net_58),
		.c(new_net_3523),
		.d(new_net_59)
	);

	bfr new_net_3524_bfr_before (
		.din(new_net_3524),
		.dout(new_net_862)
	);

	spl2 _1229__v_fanout (
		.a(_1229_),
		.b(new_net_861),
		.c(new_net_3524)
	);

	spl2 _1004__v_fanout (
		.a(_1004_),
		.b(new_net_503),
		.c(new_net_504)
	);

	spl2 _0830__v_fanout (
		.a(_0830_),
		.b(new_net_1080),
		.c(new_net_1081)
	);

	spl3L _0948__v_fanout (
		.a(_0948_),
		.b(new_net_655),
		.c(new_net_657),
		.d(new_net_656)
	);

	bfr new_net_3525_bfr_before (
		.din(new_net_3525),
		.dout(new_net_334)
	);

	bfr new_net_3526_bfr_before (
		.din(new_net_3526),
		.dout(new_net_3525)
	);

	spl2 _0752__v_fanout (
		.a(_0752_),
		.b(new_net_333),
		.c(new_net_3526)
	);

	spl2 _1200__v_fanout (
		.a(_1200_),
		.b(new_net_1402),
		.c(new_net_1403)
	);

	spl4L new_net_2002_v_fanout (
		.a(new_net_2002),
		.b(new_net_613),
		.c(new_net_627),
		.d(new_net_621),
		.e(new_net_2000)
	);

	spl2 _1025__v_fanout (
		.a(_1025_),
		.b(new_net_694),
		.c(new_net_695)
	);

	spl2 _0043__v_fanout (
		.a(_0043_),
		.b(new_net_1487),
		.c(new_net_1488)
	);

	spl2 new_net_1997_v_fanout (
		.a(new_net_1997),
		.b(new_net_2001),
		.c(new_net_1998)
	);

	spl2 _0787__v_fanout (
		.a(_0787_),
		.b(new_net_949),
		.c(new_net_950)
	);

	spl2 _0698__v_fanout (
		.a(_0698_),
		.b(new_net_171),
		.c(new_net_172)
	);

	bfr new_net_3527_bfr_before (
		.din(new_net_3527),
		.dout(new_net_443)
	);

	spl2 _0630__v_fanout (
		.a(_0630_),
		.b(new_net_442),
		.c(new_net_3527)
	);

	bfr new_net_3528_bfr_before (
		.din(new_net_3528),
		.dout(new_net_1512)
	);

	bfr new_net_3529_bfr_before (
		.din(new_net_3529),
		.dout(new_net_3528)
	);

	bfr new_net_3530_bfr_before (
		.din(new_net_3530),
		.dout(new_net_3529)
	);

	bfr new_net_3531_bfr_before (
		.din(new_net_3531),
		.dout(new_net_3530)
	);

	spl2 _0753__v_fanout (
		.a(_0753_),
		.b(new_net_1511),
		.c(new_net_3531)
	);

	spl2 _0737__v_fanout (
		.a(_0737_),
		.b(new_net_1644),
		.c(new_net_1645)
	);

	bfr new_net_3532_bfr_before (
		.din(new_net_3532),
		.dout(new_net_2027)
	);

	spl3L _0638__v_fanout (
		.a(_0638_),
		.b(new_net_558),
		.c(new_net_561),
		.d(new_net_3532)
	);

	bfr new_net_3533_bfr_before (
		.din(new_net_3533),
		.dout(new_net_2028)
	);

	bfr new_net_3534_bfr_before (
		.din(new_net_3534),
		.dout(new_net_3533)
	);

	bfr new_net_3535_bfr_before (
		.din(new_net_3535),
		.dout(new_net_3534)
	);

	bfr new_net_3536_bfr_before (
		.din(new_net_3536),
		.dout(new_net_3535)
	);

	bfr new_net_3537_bfr_before (
		.din(new_net_3537),
		.dout(new_net_3536)
	);

	spl3L _0953__v_fanout (
		.a(_0953_),
		.b(new_net_3537),
		.c(new_net_1131),
		.d(new_net_1133)
	);

	spl2 _0846__v_fanout (
		.a(_0846_),
		.b(new_net_925),
		.c(new_net_926)
	);

	bfr new_net_3538_bfr_before (
		.din(new_net_3538),
		.dout(new_net_479)
	);

	bfr new_net_3539_bfr_before (
		.din(new_net_3539),
		.dout(new_net_3538)
	);

	bfr new_net_3540_bfr_before (
		.din(new_net_3540),
		.dout(new_net_3539)
	);

	bfr new_net_3541_bfr_before (
		.din(new_net_3541),
		.dout(new_net_3540)
	);

	bfr new_net_3542_bfr_before (
		.din(new_net_3542),
		.dout(new_net_3541)
	);

	bfr new_net_3543_bfr_before (
		.din(new_net_3543),
		.dout(new_net_3542)
	);

	bfr new_net_3544_bfr_before (
		.din(new_net_3544),
		.dout(new_net_3543)
	);

	spl3L _0759__v_fanout (
		.a(_0759_),
		.b(new_net_477),
		.c(new_net_3544),
		.d(new_net_478)
	);

	spl3L _0924__v_fanout (
		.a(_0924_),
		.b(new_net_1462),
		.c(new_net_1464),
		.d(new_net_1463)
	);

	spl2 _1179__v_fanout (
		.a(_1179_),
		.b(new_net_1318),
		.c(new_net_1319)
	);

	bfr new_net_3545_bfr_before (
		.din(new_net_3545),
		.dout(new_net_603)
	);

	bfr new_net_3546_bfr_before (
		.din(new_net_3546),
		.dout(new_net_3545)
	);

	spl3L _0744__v_fanout (
		.a(_0744_),
		.b(new_net_3546),
		.c(new_net_604),
		.d(new_net_605)
	);

	spl2 _0034__v_fanout (
		.a(_0034_),
		.b(new_net_241),
		.c(new_net_242)
	);

	bfr new_net_3547_bfr_before (
		.din(new_net_3547),
		.dout(new_net_365)
	);

	bfr new_net_3548_bfr_before (
		.din(new_net_3548),
		.dout(new_net_3547)
	);

	bfr new_net_3549_bfr_before (
		.din(new_net_3549),
		.dout(new_net_3548)
	);

	bfr new_net_3550_bfr_before (
		.din(new_net_3550),
		.dout(new_net_3549)
	);

	bfr new_net_3551_bfr_before (
		.din(new_net_3551),
		.dout(new_net_3550)
	);

	bfr new_net_3552_bfr_before (
		.din(new_net_3552),
		.dout(new_net_3551)
	);

	spl2 _0758__v_fanout (
		.a(_0758_),
		.b(new_net_364),
		.c(new_net_3552)
	);

	bfr new_net_3553_bfr_before (
		.din(new_net_3553),
		.dout(new_net_2024)
	);

	bfr new_net_3554_bfr_before (
		.din(new_net_3554),
		.dout(new_net_3553)
	);

	bfr new_net_3555_bfr_before (
		.din(new_net_3555),
		.dout(new_net_3554)
	);

	spl2 _0941__v_fanout (
		.a(_0941_),
		.b(new_net_1588),
		.c(new_net_3555)
	);

	bfr new_net_3556_bfr_before (
		.din(new_net_3556),
		.dout(new_net_1510)
	);

	spl2 _0736__v_fanout (
		.a(_0736_),
		.b(new_net_1509),
		.c(new_net_3556)
	);

	bfr new_net_3557_bfr_before (
		.din(new_net_3557),
		.dout(new_net_781)
	);

	spl2 _0868__v_fanout (
		.a(_0868_),
		.b(new_net_3557),
		.c(new_net_2029)
	);

	bfr new_net_3558_bfr_before (
		.din(new_net_3558),
		.dout(new_net_1104)
	);

	bfr new_net_3559_bfr_before (
		.din(new_net_3559),
		.dout(new_net_3558)
	);

	spl2 _0667__v_fanout (
		.a(_0667_),
		.b(new_net_1103),
		.c(new_net_3559)
	);

	spl2 _1170__v_fanout (
		.a(_1170_),
		.b(new_net_1646),
		.c(new_net_1647)
	);

	spl2 _0872__v_fanout (
		.a(_0872_),
		.b(new_net_2030),
		.c(new_net_2031)
	);

	bfr new_net_3560_bfr_before (
		.din(new_net_3560),
		.dout(new_net_641)
	);

	bfr new_net_3561_bfr_before (
		.din(new_net_3561),
		.dout(new_net_3560)
	);

	spl3L _0639__v_fanout (
		.a(_0639_),
		.b(new_net_640),
		.c(new_net_642),
		.d(new_net_3561)
	);

	spl2 _0124__v_fanout (
		.a(_0124_),
		.b(new_net_394),
		.c(new_net_395)
	);

	spl2 _0055__v_fanout (
		.a(_0055_),
		.b(new_net_636),
		.c(new_net_637)
	);

	bfr new_net_3562_bfr_before (
		.din(new_net_3562),
		.dout(new_net_43)
	);

	bfr new_net_3563_bfr_before (
		.din(new_net_3563),
		.dout(new_net_3562)
	);

	spl3L _0947__v_fanout (
		.a(_0947_),
		.b(new_net_3563),
		.c(new_net_45),
		.d(new_net_44)
	);

	spl2 _0809__v_fanout (
		.a(_0809_),
		.b(new_net_1427),
		.c(new_net_1428)
	);

	bfr new_net_3564_bfr_before (
		.din(new_net_3564),
		.dout(new_net_371)
	);

	spl2 _0668__v_fanout (
		.a(_0668_),
		.b(new_net_370),
		.c(new_net_3564)
	);

	bfr new_net_3565_bfr_after (
		.din(_1191_),
		.dout(new_net_3565)
	);

	bfr new_net_3566_bfr_after (
		.din(new_net_3565),
		.dout(new_net_3566)
	);

	bfr new_net_3567_bfr_after (
		.din(new_net_3566),
		.dout(new_net_3567)
	);

	spl2 _1191__v_fanout (
		.a(new_net_3567),
		.b(new_net_366),
		.c(new_net_367)
	);

	spl2 _0074__v_fanout (
		.a(_0074_),
		.b(new_net_218),
		.c(new_net_219)
	);

	spl2 _1143__v_fanout (
		.a(_1143_),
		.b(new_net_1408),
		.c(new_net_1409)
	);

	spl2 _1209__v_fanout (
		.a(_1209_),
		.b(new_net_595),
		.c(new_net_596)
	);

	spl2 new_net_2016_v_fanout (
		.a(new_net_2016),
		.b(new_net_245),
		.c(new_net_247)
	);

	spl2 _0654__v_fanout (
		.a(_0654_),
		.b(new_net_845),
		.c(new_net_846)
	);

	spl2 _1134__v_fanout (
		.a(_1134_),
		.b(new_net_470),
		.c(new_net_471)
	);

	bfr new_net_3568_bfr_before (
		.din(new_net_3568),
		.dout(new_net_2026)
	);

	bfr new_net_3569_bfr_before (
		.din(new_net_3569),
		.dout(new_net_3568)
	);

	bfr new_net_3570_bfr_before (
		.din(new_net_3570),
		.dout(new_net_3569)
	);

	spl2 _0942__v_fanout (
		.a(_0942_),
		.b(new_net_3570),
		.c(new_net_1601)
	);

	spl4L _0985__v_fanout (
		.a(_0985_),
		.b(new_net_736),
		.c(new_net_737),
		.d(new_net_738),
		.e(new_net_735)
	);

	spl2 new_net_2022_v_fanout (
		.a(new_net_2022),
		.b(new_net_844),
		.c(new_net_843)
	);

	bfr new_net_3571_bfr_after (
		.din(_0967_),
		.dout(new_net_3571)
	);

	bfr new_net_3572_bfr_before (
		.din(new_net_3572),
		.dout(new_net_2021)
	);

	spl2 _0967__v_fanout (
		.a(new_net_3571),
		.b(new_net_3572),
		.c(new_net_452)
	);

	spl3L _0681__v_fanout (
		.a(_0681_),
		.b(new_net_1685),
		.c(new_net_1686),
		.d(new_net_1687)
	);

	bfr new_net_3573_bfr_before (
		.din(new_net_3573),
		.dout(new_net_2011)
	);

	bfr new_net_3574_bfr_before (
		.din(new_net_3574),
		.dout(new_net_3573)
	);

	bfr new_net_3575_bfr_before (
		.din(new_net_3575),
		.dout(new_net_3574)
	);

	bfr new_net_3576_bfr_before (
		.din(new_net_3576),
		.dout(new_net_3575)
	);

	bfr new_net_3577_bfr_before (
		.din(new_net_3577),
		.dout(new_net_3576)
	);

	bfr new_net_3578_bfr_before (
		.din(new_net_3578),
		.dout(new_net_3577)
	);

	bfr new_net_3579_bfr_before (
		.din(new_net_3579),
		.dout(new_net_3578)
	);

	bfr new_net_3580_bfr_before (
		.din(new_net_3580),
		.dout(new_net_3579)
	);

	bfr new_net_3581_bfr_before (
		.din(new_net_3581),
		.dout(new_net_3580)
	);

	bfr new_net_3582_bfr_before (
		.din(new_net_3582),
		.dout(new_net_3581)
	);

	bfr new_net_3583_bfr_before (
		.din(new_net_3583),
		.dout(new_net_3582)
	);

	bfr new_net_3584_bfr_before (
		.din(new_net_3584),
		.dout(new_net_3583)
	);

	bfr new_net_3585_bfr_before (
		.din(new_net_3585),
		.dout(new_net_3584)
	);

	bfr new_net_3586_bfr_before (
		.din(new_net_3586),
		.dout(new_net_3585)
	);

	bfr new_net_3587_bfr_before (
		.din(new_net_3587),
		.dout(new_net_3586)
	);

	bfr new_net_3588_bfr_before (
		.din(new_net_3588),
		.dout(new_net_3587)
	);

	bfr new_net_3589_bfr_before (
		.din(new_net_3589),
		.dout(new_net_3588)
	);

	bfr new_net_3590_bfr_before (
		.din(new_net_3590),
		.dout(new_net_3589)
	);

	spl4L new_net_2013_v_fanout (
		.a(new_net_2013),
		.b(new_net_307),
		.c(new_net_3590),
		.d(new_net_308),
		.e(new_net_312)
	);

	bfr new_net_3591_bfr_before (
		.din(new_net_3591),
		.dout(new_net_1057)
	);

	bfr new_net_3592_bfr_before (
		.din(new_net_3592),
		.dout(new_net_3591)
	);

	spl2 _1042__v_fanout (
		.a(_1042_),
		.b(new_net_1056),
		.c(new_net_3592)
	);

	spl2 new_net_1778_v_fanout (
		.a(new_net_1778),
		.b(new_net_1254),
		.c(new_net_1256)
	);

	spl2 _0906__v_fanout (
		.a(_0906_),
		.b(new_net_842),
		.c(new_net_2022)
	);

	spl2 _0660__v_fanout (
		.a(_0660_),
		.b(new_net_923),
		.c(new_net_924)
	);

	bfr new_net_3593_bfr_after (
		.din(_1155_),
		.dout(new_net_3593)
	);

	spl2 _1155__v_fanout (
		.a(new_net_3593),
		.b(new_net_1709),
		.c(new_net_1710)
	);

	spl2 new_net_2007_v_fanout (
		.a(new_net_2007),
		.b(new_net_538),
		.c(new_net_537)
	);

	bfr new_net_3594_bfr_before (
		.din(new_net_3594),
		.dout(new_net_554)
	);

	bfr new_net_3595_bfr_before (
		.din(new_net_3595),
		.dout(new_net_3594)
	);

	spl2 new_net_2018_v_fanout (
		.a(new_net_2018),
		.b(new_net_3595),
		.c(new_net_555)
	);

	bfr new_net_3596_bfr_before (
		.din(new_net_3596),
		.dout(new_net_1731)
	);

	bfr new_net_3597_bfr_before (
		.din(new_net_3597),
		.dout(new_net_3596)
	);

	bfr new_net_3598_bfr_before (
		.din(new_net_3598),
		.dout(new_net_3597)
	);

	bfr new_net_3599_bfr_before (
		.din(new_net_3599),
		.dout(new_net_3598)
	);

	bfr new_net_3600_bfr_before (
		.din(new_net_3600),
		.dout(new_net_3599)
	);

	bfr new_net_3601_bfr_before (
		.din(new_net_3601),
		.dout(new_net_1231)
	);

	bfr new_net_3602_bfr_before (
		.din(new_net_3602),
		.dout(new_net_3601)
	);

	spl4L new_net_1741_v_fanout (
		.a(new_net_1741),
		.b(new_net_3600),
		.c(new_net_1221),
		.d(new_net_3602),
		.e(new_net_1216)
	);

	bfr new_net_3603_bfr_before (
		.din(new_net_3603),
		.dout(new_net_2016)
	);

	spl3L new_net_2015_v_fanout (
		.a(new_net_2015),
		.b(new_net_250),
		.c(new_net_252),
		.d(new_net_3603)
	);

	bfr new_net_3604_bfr_after (
		.din(new_net_27),
		.dout(new_net_3604)
	);

	bfr new_net_3605_bfr_after (
		.din(new_net_3604),
		.dout(new_net_3605)
	);

	bfr new_net_3606_bfr_after (
		.din(new_net_3605),
		.dout(new_net_3606)
	);

	bfr new_net_3607_bfr_after (
		.din(new_net_3606),
		.dout(new_net_3607)
	);

	bfr new_net_3608_bfr_after (
		.din(new_net_3607),
		.dout(new_net_3608)
	);

	bfr new_net_3609_bfr_after (
		.din(new_net_3608),
		.dout(new_net_3609)
	);

	bfr new_net_3610_bfr_after (
		.din(new_net_3609),
		.dout(new_net_3610)
	);

	bfr new_net_3611_bfr_after (
		.din(new_net_3610),
		.dout(new_net_3611)
	);

	bfr new_net_3612_bfr_after (
		.din(new_net_3611),
		.dout(new_net_3612)
	);

	bfr new_net_3613_bfr_after (
		.din(new_net_3612),
		.dout(new_net_3613)
	);

	bfr new_net_3614_bfr_after (
		.din(new_net_3613),
		.dout(new_net_3614)
	);

	bfr new_net_3615_bfr_after (
		.din(new_net_3614),
		.dout(new_net_3615)
	);

	bfr new_net_3616_bfr_after (
		.din(new_net_3615),
		.dout(new_net_3616)
	);

	bfr new_net_3617_bfr_after (
		.din(new_net_3616),
		.dout(new_net_3617)
	);

	bfr new_net_3618_bfr_after (
		.din(new_net_3617),
		.dout(new_net_3618)
	);

	bfr new_net_3619_bfr_after (
		.din(new_net_3618),
		.dout(new_net_3619)
	);

	bfr new_net_3620_bfr_after (
		.din(new_net_3619),
		.dout(new_net_3620)
	);

	bfr new_net_3621_bfr_after (
		.din(new_net_3620),
		.dout(new_net_3621)
	);

	bfr new_net_3622_bfr_after (
		.din(new_net_3621),
		.dout(new_net_3622)
	);

	bfr new_net_3623_bfr_after (
		.din(new_net_3622),
		.dout(new_net_3623)
	);

	bfr new_net_3624_bfr_after (
		.din(new_net_3623),
		.dout(new_net_3624)
	);

	bfr new_net_3625_bfr_after (
		.din(new_net_3624),
		.dout(new_net_3625)
	);

	bfr new_net_3626_bfr_after (
		.din(new_net_3625),
		.dout(new_net_3626)
	);

	bfr new_net_3627_bfr_after (
		.din(new_net_3626),
		.dout(new_net_3627)
	);

	bfr new_net_3628_bfr_after (
		.din(new_net_3627),
		.dout(new_net_3628)
	);

	bfr new_net_3629_bfr_after (
		.din(new_net_3628),
		.dout(new_net_3629)
	);

	bfr new_net_3630_bfr_after (
		.din(new_net_3629),
		.dout(new_net_3630)
	);

	bfr new_net_3631_bfr_after (
		.din(new_net_3630),
		.dout(new_net_3631)
	);

	bfr new_net_3632_bfr_after (
		.din(new_net_3631),
		.dout(new_net_3632)
	);

	bfr new_net_3633_bfr_after (
		.din(new_net_3632),
		.dout(new_net_3633)
	);

	bfr new_net_3634_bfr_after (
		.din(new_net_3633),
		.dout(new_net_3634)
	);

	bfr new_net_3635_bfr_after (
		.din(new_net_3634),
		.dout(new_net_3635)
	);

	bfr new_net_3636_bfr_after (
		.din(new_net_3635),
		.dout(new_net_3636)
	);

	bfr new_net_3637_bfr_after (
		.din(new_net_3636),
		.dout(new_net_3637)
	);

	bfr new_net_3638_bfr_after (
		.din(new_net_3637),
		.dout(new_net_3638)
	);

	spl2 new_net_27_v_fanout (
		.a(new_net_3638),
		.b(G5229),
		.c(G5230)
	);

	spl4L new_net_2010_v_fanout (
		.a(new_net_2010),
		.b(new_net_35),
		.c(new_net_34),
		.d(new_net_33),
		.e(new_net_38)
	);

	bfr new_net_3639_bfr_before (
		.din(new_net_3639),
		.dout(new_net_654)
	);

	spl2 _0728__v_fanout (
		.a(_0728_),
		.b(new_net_653),
		.c(new_net_3639)
	);

	spl4L new_net_1742_v_fanout (
		.a(new_net_1742),
		.b(new_net_1238),
		.c(new_net_1207),
		.d(new_net_1237),
		.e(new_net_1214)
	);

	spl2 new_net_2008_v_fanout (
		.a(new_net_2008),
		.b(new_net_786),
		.c(new_net_785)
	);

	spl2 _0934__v_fanout (
		.a(_0934_),
		.b(new_net_777),
		.c(new_net_778)
	);

	spl2 _0931__v_fanout (
		.a(_0931_),
		.b(new_net_1383),
		.c(new_net_1384)
	);

	bfr new_net_3640_bfr_before (
		.din(new_net_3640),
		.dout(new_net_37)
	);

	bfr new_net_3641_bfr_before (
		.din(new_net_3641),
		.dout(new_net_3640)
	);

	bfr new_net_3642_bfr_before (
		.din(new_net_3642),
		.dout(new_net_3641)
	);

	bfr new_net_3643_bfr_before (
		.din(new_net_3643),
		.dout(new_net_3642)
	);

	spl2 new_net_2009_v_fanout (
		.a(new_net_2009),
		.b(new_net_36),
		.c(new_net_3643)
	);

	spl2 new_net_2014_v_fanout (
		.a(new_net_2014),
		.b(new_net_1093),
		.c(new_net_1092)
	);

	bfr new_net_3644_bfr_after (
		.din(_0064_),
		.dout(new_net_3644)
	);

	spl2 _0064__v_fanout (
		.a(new_net_3644),
		.b(new_net_39),
		.c(new_net_40)
	);

	spl3L _0745__v_fanout (
		.a(_0745_),
		.b(new_net_202),
		.c(new_net_203),
		.d(new_net_204)
	);

	spl4L _0612__v_fanout (
		.a(_0612_),
		.b(new_net_64),
		.c(new_net_62),
		.d(new_net_63),
		.e(new_net_61)
	);

	bfr new_net_3645_bfr_before (
		.din(new_net_3645),
		.dout(new_net_1211)
	);

	bfr new_net_3646_bfr_before (
		.din(new_net_3646),
		.dout(new_net_1203)
	);

	spl3L new_net_1743_v_fanout (
		.a(new_net_1743),
		.b(new_net_3645),
		.c(new_net_1226),
		.d(new_net_3646)
	);

	bfr new_net_3647_bfr_before (
		.din(new_net_3647),
		.dout(new_net_2023)
	);

	bfr new_net_3648_bfr_before (
		.din(new_net_3648),
		.dout(new_net_3647)
	);

	bfr new_net_3649_bfr_before (
		.din(new_net_3649),
		.dout(new_net_3648)
	);

	bfr new_net_3650_bfr_before (
		.din(new_net_3650),
		.dout(new_net_3649)
	);

	bfr new_net_3651_bfr_before (
		.din(new_net_3651),
		.dout(new_net_3650)
	);

	spl2 _0661__v_fanout (
		.a(_0661_),
		.b(new_net_1345),
		.c(new_net_3651)
	);

	spl3L new_net_2012_v_fanout (
		.a(new_net_2012),
		.b(new_net_309),
		.c(new_net_305),
		.d(new_net_311)
	);

	spl2 new_net_2020_v_fanout (
		.a(new_net_2020),
		.b(new_net_684),
		.c(new_net_683)
	);

	bfr new_net_3652_bfr_before (
		.din(new_net_3652),
		.dout(new_net_1223)
	);

	spl2 new_net_1730_v_fanout (
		.a(new_net_1730),
		.b(new_net_3652),
		.c(new_net_1235)
	);

	spl3L new_net_1996_v_fanout (
		.a(new_net_1996),
		.b(new_net_2002),
		.c(new_net_1997),
		.d(new_net_624)
	);

	spl3L new_net_2019_v_fanout (
		.a(new_net_2019),
		.b(new_net_553),
		.c(new_net_556),
		.d(new_net_557)
	);

	spl4L new_net_2017_v_fanout (
		.a(new_net_2017),
		.b(new_net_249),
		.c(new_net_248),
		.d(new_net_244),
		.e(new_net_243)
	);

	bfr new_net_3653_bfr_before (
		.din(new_net_3653),
		.dout(new_net_348)
	);

	bfr new_net_3654_bfr_before (
		.din(new_net_3654),
		.dout(new_net_3653)
	);

	spl2 new_net_1992_v_fanout (
		.a(new_net_1992),
		.b(new_net_3654),
		.c(new_net_347)
	);

	spl2 new_net_2006_v_fanout (
		.a(new_net_2006),
		.b(new_net_486),
		.c(new_net_485)
	);

	spl4L _0946__v_fanout (
		.a(_0946_),
		.b(new_net_501),
		.c(new_net_500),
		.d(new_net_502),
		.e(new_net_499)
	);

	spl2 _0862__v_fanout (
		.a(_0862_),
		.b(new_net_2009),
		.c(new_net_2010)
	);

	spl3L _0952__v_fanout (
		.a(_0952_),
		.b(new_net_158),
		.c(new_net_160),
		.d(new_net_159)
	);

	bfr new_net_3655_bfr_before (
		.din(new_net_3655),
		.dout(new_net_1234)
	);

	bfr new_net_3656_bfr_before (
		.din(new_net_3656),
		.dout(new_net_3655)
	);

	bfr new_net_3657_bfr_before (
		.din(new_net_3657),
		.dout(new_net_1741)
	);

	bfr new_net_3658_bfr_before (
		.din(new_net_3658),
		.dout(new_net_1742)
	);

	spl4L new_net_1744_v_fanout (
		.a(new_net_1744),
		.b(new_net_3657),
		.c(new_net_3658),
		.d(new_net_1743),
		.e(new_net_3656)
	);

	bfr new_net_3659_bfr_before (
		.din(new_net_3659),
		.dout(new_net_1229)
	);

	bfr new_net_3660_bfr_before (
		.din(new_net_3660),
		.dout(new_net_3659)
	);

	bfr new_net_3661_bfr_before (
		.din(new_net_3661),
		.dout(new_net_1240)
	);

	spl3L new_net_1729_v_fanout (
		.a(new_net_1729),
		.b(new_net_3660),
		.c(new_net_3661),
		.d(new_net_1730)
	);

	bfr new_net_3662_bfr_after (
		.din(_0153_),
		.dout(new_net_3662)
	);

	bfr new_net_3663_bfr_after (
		.din(new_net_3662),
		.dout(new_net_3663)
	);

	bfr new_net_3664_bfr_after (
		.din(new_net_3663),
		.dout(new_net_3664)
	);

	spl2 _0153__v_fanout (
		.a(new_net_3664),
		.b(new_net_1127),
		.c(new_net_1128)
	);

	spl3L _0735__v_fanout (
		.a(_0735_),
		.b(new_net_784),
		.c(new_net_2008),
		.d(new_net_787)
	);

	spl2 _0135__v_fanout (
		.a(_0135_),
		.b(new_net_566),
		.c(new_net_567)
	);

	spl4L _0757__v_fanout (
		.a(_0757_),
		.b(new_net_264),
		.c(new_net_263),
		.d(new_net_265),
		.e(new_net_262)
	);

	spl4L _0940__v_fanout (
		.a(_0940_),
		.b(new_net_1565),
		.c(new_net_1567),
		.d(new_net_1566),
		.e(new_net_1564)
	);

	spl2 new_net_1901_v_fanout (
		.a(new_net_1901),
		.b(new_net_962),
		.c(new_net_964)
	);

	spl2 _0583__v_fanout (
		.a(_0583_),
		.b(new_net_2013),
		.c(new_net_2012)
	);

	spl2 new_net_1840_v_fanout (
		.a(new_net_1840),
		.b(new_net_903),
		.c(new_net_904)
	);

	spl3L _0666__v_fanout (
		.a(_0666_),
		.b(new_net_2014),
		.c(new_net_1090),
		.d(new_net_1091)
	);

	spl2 new_net_1786_v_fanout (
		.a(new_net_1786),
		.b(new_net_1194),
		.c(new_net_1196)
	);

	spl4L _0580__v_fanout (
		.a(_0580_),
		.b(new_net_251),
		.c(new_net_2017),
		.d(new_net_2015),
		.e(new_net_246)
	);

	spl2 _0144__v_fanout (
		.a(_0144_),
		.b(new_net_703),
		.c(new_net_704)
	);

	bfr new_net_3665_bfr_after (
		.din(_0168_),
		.dout(new_net_3665)
	);

	bfr new_net_3666_bfr_after (
		.din(new_net_3665),
		.dout(new_net_3666)
	);

	bfr new_net_3667_bfr_after (
		.din(new_net_3666),
		.dout(new_net_3667)
	);

	bfr new_net_3668_bfr_after (
		.din(new_net_3667),
		.dout(new_net_3668)
	);

	spl2 _0168__v_fanout (
		.a(new_net_3668),
		.b(new_net_886),
		.c(new_net_887)
	);

	spl2 _0596__v_fanout (
		.a(_0596_),
		.b(new_net_2019),
		.c(new_net_2018)
	);

	spl2 new_net_1905_v_fanout (
		.a(new_net_1905),
		.b(new_net_917),
		.c(new_net_919)
	);

	spl3L _0637__v_fanout (
		.a(_0637_),
		.b(new_net_536),
		.c(new_net_539),
		.d(new_net_2007)
	);

	spl4L _0855__v_fanout (
		.a(_0855_),
		.b(new_net_227),
		.c(new_net_226),
		.d(new_net_225),
		.e(new_net_224)
	);

	spl4L _0751__v_fanout (
		.a(_0751_),
		.b(new_net_316),
		.c(new_net_315),
		.d(new_net_314),
		.e(new_net_313)
	);

	spl3L _0867__v_fanout (
		.a(_0867_),
		.b(new_net_682),
		.c(new_net_2020),
		.d(new_net_685)
	);

	spl2 new_net_1993_v_fanout (
		.a(new_net_1993),
		.b(new_net_1020),
		.c(new_net_1019)
	);

	spl2 new_net_1868_v_fanout (
		.a(new_net_1868),
		.b(new_net_1265),
		.c(new_net_1268)
	);

	spl4L _0604__v_fanout (
		.a(_0604_),
		.b(new_net_688),
		.c(new_net_687),
		.d(new_net_689),
		.e(new_net_686)
	);

	spl2 _0679__v_fanout (
		.a(_0679_),
		.b(new_net_1387),
		.c(new_net_1388)
	);

	spl4L new_net_1915_v_fanout (
		.a(new_net_1915),
		.b(new_net_89),
		.c(new_net_91),
		.d(new_net_103),
		.e(new_net_101)
	);

	spl2 new_net_1769_v_fanout (
		.a(new_net_1769),
		.b(new_net_1279),
		.c(new_net_1278)
	);

	spl2 _0111__v_fanout (
		.a(_0111_),
		.b(new_net_139),
		.c(new_net_140)
	);

	bfr new_net_3669_bfr_before (
		.din(new_net_3669),
		.dout(G5215)
	);

	bfr new_net_3670_bfr_before (
		.din(new_net_3670),
		.dout(new_net_3669)
	);

	bfr new_net_3671_bfr_before (
		.din(new_net_3671),
		.dout(new_net_3670)
	);

	bfr new_net_3672_bfr_before (
		.din(new_net_3672),
		.dout(new_net_3671)
	);

	bfr new_net_3673_bfr_before (
		.din(new_net_3673),
		.dout(new_net_3672)
	);

	bfr new_net_3674_bfr_before (
		.din(new_net_3674),
		.dout(new_net_3673)
	);

	bfr new_net_3675_bfr_before (
		.din(new_net_3675),
		.dout(new_net_3674)
	);

	bfr new_net_3676_bfr_before (
		.din(new_net_3676),
		.dout(new_net_3675)
	);

	bfr new_net_3677_bfr_before (
		.din(new_net_3677),
		.dout(new_net_3676)
	);

	bfr new_net_3678_bfr_before (
		.din(new_net_3678),
		.dout(new_net_3677)
	);

	bfr new_net_3679_bfr_before (
		.din(new_net_3679),
		.dout(new_net_3678)
	);

	bfr new_net_3680_bfr_before (
		.din(new_net_3680),
		.dout(new_net_3679)
	);

	bfr new_net_3681_bfr_before (
		.din(new_net_3681),
		.dout(new_net_3680)
	);

	bfr new_net_3682_bfr_before (
		.din(new_net_3682),
		.dout(new_net_3681)
	);

	bfr new_net_3683_bfr_before (
		.din(new_net_3683),
		.dout(new_net_3682)
	);

	bfr new_net_3684_bfr_before (
		.din(new_net_3684),
		.dout(new_net_3683)
	);

	bfr new_net_3685_bfr_before (
		.din(new_net_3685),
		.dout(new_net_3684)
	);

	bfr new_net_3686_bfr_before (
		.din(new_net_3686),
		.dout(new_net_3685)
	);

	bfr new_net_3687_bfr_before (
		.din(new_net_3687),
		.dout(new_net_3686)
	);

	bfr new_net_3688_bfr_before (
		.din(new_net_3688),
		.dout(new_net_3687)
	);

	bfr new_net_3689_bfr_before (
		.din(new_net_3689),
		.dout(new_net_3688)
	);

	bfr new_net_3690_bfr_before (
		.din(new_net_3690),
		.dout(new_net_3689)
	);

	bfr new_net_3691_bfr_before (
		.din(new_net_3691),
		.dout(new_net_3690)
	);

	bfr new_net_3692_bfr_before (
		.din(new_net_3692),
		.dout(new_net_3691)
	);

	bfr new_net_3693_bfr_before (
		.din(new_net_3693),
		.dout(new_net_3692)
	);

	bfr new_net_3694_bfr_before (
		.din(new_net_3694),
		.dout(new_net_3693)
	);

	bfr new_net_3695_bfr_before (
		.din(new_net_3695),
		.dout(new_net_3694)
	);

	bfr new_net_3696_bfr_before (
		.din(new_net_3696),
		.dout(new_net_3695)
	);

	bfr new_net_3697_bfr_before (
		.din(new_net_3697),
		.dout(new_net_3696)
	);

	bfr new_net_3698_bfr_before (
		.din(new_net_3698),
		.dout(new_net_3697)
	);

	bfr new_net_3699_bfr_before (
		.din(new_net_3699),
		.dout(new_net_3698)
	);

	bfr new_net_3700_bfr_before (
		.din(new_net_3700),
		.dout(new_net_3699)
	);

	bfr new_net_3701_bfr_before (
		.din(new_net_3701),
		.dout(new_net_3700)
	);

	bfr new_net_3702_bfr_before (
		.din(new_net_3702),
		.dout(new_net_3701)
	);

	bfr new_net_3703_bfr_before (
		.din(new_net_3703),
		.dout(new_net_3702)
	);

	bfr new_net_3704_bfr_before (
		.din(new_net_3704),
		.dout(new_net_3703)
	);

	spl3L new_net_1770_v_fanout (
		.a(new_net_1770),
		.b(new_net_1273),
		.c(new_net_1274),
		.d(new_net_3704)
	);

	bfr new_net_3705_bfr_before (
		.din(new_net_3705),
		.dout(new_net_1778)
	);

	spl2 new_net_1777_v_fanout (
		.a(new_net_1777),
		.b(new_net_3705),
		.c(new_net_1257)
	);

	spl2 new_net_1787_v_fanout (
		.a(new_net_1787),
		.b(new_net_898),
		.c(new_net_899)
	);

	spl4L new_net_1912_v_fanout (
		.a(new_net_1912),
		.b(new_net_88),
		.c(new_net_99),
		.d(new_net_86),
		.e(new_net_97)
	);

	spl2 _0885__v_fanout (
		.a(_0885_),
		.b(new_net_484),
		.c(new_net_2006)
	);

	bfr new_net_3706_bfr_after (
		.din(_0138_),
		.dout(new_net_3706)
	);

	spl2 _0138__v_fanout (
		.a(new_net_3706),
		.b(new_net_1188),
		.c(new_net_1189)
	);

	bfr new_net_3707_bfr_before (
		.din(new_net_3707),
		.dout(new_net_1120)
	);

	bfr new_net_3708_bfr_before (
		.din(new_net_3708),
		.dout(new_net_3707)
	);

	spl3L _0659__v_fanout (
		.a(_0659_),
		.b(new_net_1119),
		.c(new_net_1121),
		.d(new_net_3708)
	);

	spl2 _0114__v_fanout (
		.a(_0114_),
		.b(new_net_187),
		.c(new_net_188)
	);

	bfr new_net_3709_bfr_before (
		.din(new_net_3709),
		.dout(G5221)
	);

	bfr new_net_3710_bfr_before (
		.din(new_net_3710),
		.dout(new_net_3709)
	);

	bfr new_net_3711_bfr_before (
		.din(new_net_3711),
		.dout(new_net_3710)
	);

	bfr new_net_3712_bfr_before (
		.din(new_net_3712),
		.dout(new_net_3711)
	);

	bfr new_net_3713_bfr_before (
		.din(new_net_3713),
		.dout(new_net_3712)
	);

	bfr new_net_3714_bfr_before (
		.din(new_net_3714),
		.dout(new_net_3713)
	);

	bfr new_net_3715_bfr_before (
		.din(new_net_3715),
		.dout(new_net_3714)
	);

	bfr new_net_3716_bfr_before (
		.din(new_net_3716),
		.dout(new_net_3715)
	);

	bfr new_net_3717_bfr_before (
		.din(new_net_3717),
		.dout(new_net_3716)
	);

	bfr new_net_3718_bfr_before (
		.din(new_net_3718),
		.dout(new_net_3717)
	);

	bfr new_net_3719_bfr_before (
		.din(new_net_3719),
		.dout(new_net_3718)
	);

	bfr new_net_3720_bfr_before (
		.din(new_net_3720),
		.dout(new_net_3719)
	);

	bfr new_net_3721_bfr_before (
		.din(new_net_3721),
		.dout(new_net_3720)
	);

	bfr new_net_3722_bfr_before (
		.din(new_net_3722),
		.dout(new_net_3721)
	);

	bfr new_net_3723_bfr_before (
		.din(new_net_3723),
		.dout(new_net_3722)
	);

	bfr new_net_3724_bfr_before (
		.din(new_net_3724),
		.dout(new_net_3723)
	);

	bfr new_net_3725_bfr_before (
		.din(new_net_3725),
		.dout(new_net_3724)
	);

	bfr new_net_3726_bfr_before (
		.din(new_net_3726),
		.dout(new_net_3725)
	);

	bfr new_net_3727_bfr_before (
		.din(new_net_3727),
		.dout(new_net_3726)
	);

	bfr new_net_3728_bfr_before (
		.din(new_net_3728),
		.dout(new_net_3727)
	);

	bfr new_net_3729_bfr_before (
		.din(new_net_3729),
		.dout(new_net_3728)
	);

	bfr new_net_3730_bfr_before (
		.din(new_net_3730),
		.dout(new_net_3729)
	);

	bfr new_net_3731_bfr_before (
		.din(new_net_3731),
		.dout(new_net_3730)
	);

	bfr new_net_3732_bfr_before (
		.din(new_net_3732),
		.dout(new_net_3731)
	);

	bfr new_net_3733_bfr_before (
		.din(new_net_3733),
		.dout(new_net_3732)
	);

	bfr new_net_3734_bfr_before (
		.din(new_net_3734),
		.dout(new_net_3733)
	);

	bfr new_net_3735_bfr_before (
		.din(new_net_3735),
		.dout(new_net_3734)
	);

	bfr new_net_3736_bfr_before (
		.din(new_net_3736),
		.dout(new_net_3735)
	);

	bfr new_net_3737_bfr_before (
		.din(new_net_3737),
		.dout(new_net_3736)
	);

	bfr new_net_3738_bfr_before (
		.din(new_net_3738),
		.dout(new_net_3737)
	);

	bfr new_net_3739_bfr_before (
		.din(new_net_3739),
		.dout(new_net_3738)
	);

	bfr new_net_3740_bfr_before (
		.din(new_net_3740),
		.dout(new_net_3739)
	);

	bfr new_net_3741_bfr_before (
		.din(new_net_3741),
		.dout(new_net_3740)
	);

	bfr new_net_3742_bfr_before (
		.din(new_net_3742),
		.dout(new_net_3741)
	);

	bfr new_net_3743_bfr_before (
		.din(new_net_3743),
		.dout(new_net_3742)
	);

	bfr new_net_3744_bfr_before (
		.din(new_net_3744),
		.dout(new_net_3743)
	);

	bfr new_net_3745_bfr_before (
		.din(new_net_3745),
		.dout(new_net_3744)
	);

	spl3L new_net_1933_v_fanout (
		.a(new_net_1933),
		.b(new_net_912),
		.c(new_net_913),
		.d(new_net_3745)
	);

	spl2 _0929__v_fanout (
		.a(_0929_),
		.b(new_net_1343),
		.c(new_net_1344)
	);

	bfr new_net_3746_bfr_after (
		.din(_0127_),
		.dout(new_net_3746)
	);

	bfr new_net_3747_bfr_after (
		.din(new_net_3746),
		.dout(new_net_3747)
	);

	bfr new_net_3748_bfr_after (
		.din(new_net_3747),
		.dout(new_net_3748)
	);

	spl2 _0127__v_fanout (
		.a(new_net_3748),
		.b(new_net_135),
		.c(new_net_136)
	);

	bfr new_net_3749_bfr_before (
		.din(new_net_3749),
		.dout(new_net_257)
	);

	spl3L new_net_1995_v_fanout (
		.a(new_net_1995),
		.b(new_net_259),
		.c(new_net_261),
		.d(new_net_3749)
	);

	spl2 new_net_1762_v_fanout (
		.a(new_net_1762),
		.b(new_net_1470),
		.c(new_net_1475)
	);

	spl2 new_net_1904_v_fanout (
		.a(new_net_1904),
		.b(new_net_920),
		.c(new_net_1905)
	);

	spl4L new_net_1913_v_fanout (
		.a(new_net_1913),
		.b(new_net_100),
		.c(new_net_102),
		.d(new_net_98),
		.e(new_net_84)
	);

	spl2 _0710__v_fanout (
		.a(_0710_),
		.b(new_net_1335),
		.c(new_net_1336)
	);

	bfr new_net_3750_bfr_before (
		.din(new_net_3750),
		.dout(new_net_828)
	);

	spl3L new_net_1882_v_fanout (
		.a(new_net_1882),
		.b(new_net_826),
		.c(new_net_827),
		.d(new_net_3750)
	);

	bfr new_net_3751_bfr_after (
		.din(_0201_),
		.dout(new_net_3751)
	);

	spl2 _0201__v_fanout (
		.a(new_net_3751),
		.b(new_net_232),
		.c(new_net_233)
	);

	bfr new_net_3752_bfr_after (
		.din(_0147_),
		.dout(new_net_3752)
	);

	spl2 _0147__v_fanout (
		.a(new_net_3752),
		.b(new_net_430),
		.c(new_net_431)
	);

	spl2 new_net_1785_v_fanout (
		.a(new_net_1785),
		.b(new_net_1786),
		.c(new_net_1197)
	);

	spl4L new_net_1911_v_fanout (
		.a(new_net_1911),
		.b(new_net_93),
		.c(new_net_85),
		.d(new_net_94),
		.e(new_net_87)
	);

	spl4L new_net_1914_v_fanout (
		.a(new_net_1914),
		.b(new_net_90),
		.c(new_net_92),
		.d(new_net_95),
		.e(new_net_96)
	);

	spl2 _0031__v_fanout (
		.a(_0031_),
		.b(new_net_327),
		.c(new_net_328)
	);

	bfr new_net_3753_bfr_before (
		.din(new_net_3753),
		.dout(new_net_1094)
	);

	bfr new_net_3754_bfr_before (
		.din(new_net_3754),
		.dout(new_net_3753)
	);

	spl2 new_net_1831_v_fanout (
		.a(new_net_1831),
		.b(new_net_3754),
		.c(new_net_1096)
	);

	spl2 new_net_1994_v_fanout (
		.a(new_net_1994),
		.b(new_net_258),
		.c(new_net_260)
	);

	spl2 _0741__v_fanout (
		.a(_0741_),
		.b(new_net_362),
		.c(new_net_363)
	);

	bfr new_net_3755_bfr_before (
		.din(new_net_3755),
		.dout(new_net_1802)
	);

	bfr new_net_3756_bfr_before (
		.din(new_net_3756),
		.dout(new_net_3755)
	);

	spl2 new_net_1801_v_fanout (
		.a(new_net_1801),
		.b(new_net_3756),
		.c(new_net_591)
	);

	spl3L new_net_1917_v_fanout (
		.a(new_net_1917),
		.b(new_net_1915),
		.c(new_net_1912),
		.d(new_net_1911)
	);

	spl2 new_net_1949_v_fanout (
		.a(new_net_1949),
		.b(new_net_715),
		.c(new_net_716)
	);

	spl2 new_net_1908_v_fanout (
		.a(new_net_1908),
		.b(new_net_651),
		.c(new_net_652)
	);

	spl3L new_net_1934_v_fanout (
		.a(new_net_1934),
		.b(new_net_915),
		.c(new_net_914),
		.d(new_net_916)
	);

	spl2 _0951__v_fanout (
		.a(_0951_),
		.b(new_net_901),
		.c(new_net_902)
	);

	bfr new_net_3757_bfr_before (
		.din(new_net_3757),
		.dout(new_net_771)
	);

	spl2 new_net_1812_v_fanout (
		.a(new_net_1812),
		.b(new_net_772),
		.c(new_net_3757)
	);

	bfr new_net_3758_bfr_before (
		.din(new_net_3758),
		.dout(new_net_1208)
	);

	spl4L new_net_1745_v_fanout (
		.a(new_net_1745),
		.b(new_net_3758),
		.c(new_net_1233),
		.d(new_net_1744),
		.e(new_net_1217)
	);

	bfr new_net_3759_bfr_before (
		.din(new_net_3759),
		.dout(new_net_1055)
	);

	spl2 new_net_1863_v_fanout (
		.a(new_net_1863),
		.b(new_net_1054),
		.c(new_net_3759)
	);

	spl4L new_net_2004_v_fanout (
		.a(new_net_2004),
		.b(new_net_729),
		.c(new_net_728),
		.d(new_net_727),
		.e(new_net_725)
	);

	spl4L new_net_1950_v_fanout (
		.a(new_net_1950),
		.b(new_net_708),
		.c(new_net_709),
		.d(new_net_710),
		.e(new_net_717)
	);

	spl4L new_net_1910_v_fanout (
		.a(new_net_1910),
		.b(new_net_648),
		.c(new_net_649),
		.d(new_net_650),
		.e(new_net_647)
	);

	spl4L new_net_1990_v_fanout (
		.a(new_net_1990),
		.b(new_net_570),
		.c(new_net_571),
		.d(new_net_569),
		.e(new_net_568)
	);

	bfr new_net_3760_bfr_after (
		.din(_0742_),
		.dout(new_net_3760)
	);

	spl2 _0742__v_fanout (
		.a(new_net_3760),
		.b(new_net_156),
		.c(new_net_157)
	);

	spl4L new_net_1921_v_fanout (
		.a(new_net_1921),
		.b(new_net_761),
		.c(new_net_763),
		.d(new_net_764),
		.e(new_net_760)
	);

	spl4L new_net_1922_v_fanout (
		.a(new_net_1922),
		.b(new_net_765),
		.c(new_net_767),
		.d(new_net_766),
		.e(new_net_762)
	);

	spl4L new_net_1925_v_fanout (
		.a(new_net_1925),
		.b(new_net_300),
		.c(new_net_301),
		.d(new_net_297),
		.e(new_net_296)
	);

	bfr new_net_3761_bfr_before (
		.din(new_net_3761),
		.dout(new_net_1591)
	);

	bfr new_net_3762_bfr_before (
		.din(new_net_3762),
		.dout(new_net_3761)
	);

	spl2 new_net_1832_v_fanout (
		.a(new_net_1832),
		.b(new_net_3762),
		.c(new_net_1593)
	);

	spl2 new_net_1923_v_fanout (
		.a(new_net_1923),
		.b(new_net_302),
		.c(new_net_303)
	);

	spl2 new_net_1724_v_fanout (
		.a(new_net_1724),
		.b(new_net_1077),
		.c(new_net_1078)
	);

	bfr new_net_3763_bfr_after (
		.din(_0121_),
		.dout(new_net_3763)
	);

	spl2 _0121__v_fanout (
		.a(new_net_3763),
		.b(new_net_1159),
		.c(new_net_1160)
	);

	spl2 new_net_1916_v_fanout (
		.a(new_net_1916),
		.b(new_net_1913),
		.c(new_net_1914)
	);

	spl4L new_net_1951_v_fanout (
		.a(new_net_1951),
		.b(new_net_714),
		.c(new_net_712),
		.d(new_net_713),
		.e(new_net_711)
	);

	spl2 _0950__v_fanout (
		.a(_0950_),
		.b(new_net_127),
		.c(new_net_128)
	);

	spl4L new_net_1909_v_fanout (
		.a(new_net_1909),
		.b(new_net_645),
		.c(new_net_644),
		.d(new_net_646),
		.e(new_net_643)
	);

	spl2 new_net_1920_v_fanout (
		.a(new_net_1920),
		.b(new_net_768),
		.c(new_net_769)
	);

	spl2 new_net_2003_v_fanout (
		.a(new_net_2003),
		.b(new_net_733),
		.c(new_net_734)
	);

	spl4L new_net_1941_v_fanout (
		.a(new_net_1941),
		.b(new_net_518),
		.c(new_net_516),
		.d(new_net_517),
		.e(new_net_515)
	);

	spl4L new_net_1940_v_fanout (
		.a(new_net_1940),
		.b(new_net_513),
		.c(new_net_514),
		.d(new_net_512),
		.e(new_net_511)
	);

	spl4L new_net_1924_v_fanout (
		.a(new_net_1924),
		.b(new_net_295),
		.c(new_net_299),
		.d(new_net_298),
		.e(new_net_304)
	);

	spl4L new_net_2005_v_fanout (
		.a(new_net_2005),
		.b(new_net_730),
		.c(new_net_732),
		.d(new_net_731),
		.e(new_net_726)
	);

	spl4L new_net_1935_v_fanout (
		.a(new_net_1935),
		.b(new_net_910),
		.c(new_net_1933),
		.d(new_net_909),
		.e(new_net_908)
	);

	spl4L new_net_1938_v_fanout (
		.a(new_net_1938),
		.b(new_net_273),
		.c(new_net_275),
		.d(new_net_274),
		.e(new_net_272)
	);

	spl2 new_net_1936_v_fanout (
		.a(new_net_1936),
		.b(new_net_276),
		.c(new_net_277)
	);

	spl2 new_net_1939_v_fanout (
		.a(new_net_1939),
		.b(new_net_519),
		.c(new_net_520)
	);

	spl2 new_net_1728_v_fanout (
		.a(new_net_1728),
		.b(new_net_1729),
		.c(new_net_1239)
	);

	spl4L new_net_1937_v_fanout (
		.a(new_net_1937),
		.b(new_net_269),
		.c(new_net_271),
		.d(new_net_270),
		.e(new_net_268)
	);

	spl4L new_net_1991_v_fanout (
		.a(new_net_1991),
		.b(new_net_573),
		.c(new_net_574),
		.d(new_net_575),
		.e(new_net_572)
	);

	spl2 new_net_1761_v_fanout (
		.a(new_net_1761),
		.b(new_net_1465),
		.c(new_net_1762)
	);

	bfr new_net_3764_bfr_after (
		.din(_0930_),
		.dout(new_net_3764)
	);

	spl2 _0930__v_fanout (
		.a(new_net_3764),
		.b(new_net_448),
		.c(new_net_449)
	);

	spl2 new_net_1989_v_fanout (
		.a(new_net_1989),
		.b(new_net_576),
		.c(new_net_577)
	);

	spl3L _0266__v_fanout (
		.a(_0266_),
		.b(new_net_1910),
		.c(new_net_1909),
		.d(new_net_1908)
	);

	spl2 _0592__v_fanout (
		.a(_0592_),
		.b(new_net_1917),
		.c(new_net_1916)
	);

	bfr new_net_3765_bfr_after (
		.din(_0851_),
		.dout(new_net_3765)
	);

	bfr new_net_3766_bfr_after (
		.din(new_net_3765),
		.dout(new_net_3766)
	);

	bfr new_net_3767_bfr_after (
		.din(new_net_3766),
		.dout(new_net_3767)
	);

	bfr new_net_3768_bfr_after (
		.din(new_net_3767),
		.dout(new_net_3768)
	);

	bfr new_net_3769_bfr_after (
		.din(new_net_3768),
		.dout(new_net_3769)
	);

	bfr new_net_3770_bfr_after (
		.din(new_net_3769),
		.dout(new_net_3770)
	);

	bfr new_net_3771_bfr_after (
		.din(new_net_3770),
		.dout(new_net_3771)
	);

	bfr new_net_3772_bfr_after (
		.din(new_net_3771),
		.dout(new_net_3772)
	);

	bfr new_net_3773_bfr_after (
		.din(new_net_3772),
		.dout(new_net_3773)
	);

	bfr new_net_3774_bfr_before (
		.din(new_net_3774),
		.dout(new_net_1918)
	);

	bfr new_net_3775_bfr_before (
		.din(new_net_3775),
		.dout(new_net_3774)
	);

	bfr new_net_3776_bfr_before (
		.din(new_net_3776),
		.dout(new_net_3775)
	);

	spl2 _0851__v_fanout (
		.a(new_net_3773),
		.b(new_net_585),
		.c(new_net_3776)
	);

	spl4L new_net_1850_v_fanout (
		.a(new_net_1850),
		.b(new_net_1672),
		.c(new_net_1675),
		.d(new_net_1676),
		.e(new_net_1671)
	);

	spl2 new_net_1803_v_fanout (
		.a(new_net_1803),
		.b(new_net_1006),
		.c(new_net_1013)
	);

	spl2 new_net_1841_v_fanout (
		.a(new_net_1841),
		.b(new_net_1048),
		.c(new_net_1046)
	);

	spl3L _0093__v_fanout (
		.a(_0093_),
		.b(new_net_1920),
		.c(new_net_1921),
		.d(new_net_1922)
	);

	spl2 new_net_1760_v_fanout (
		.a(new_net_1760),
		.b(new_net_1467),
		.c(new_net_1761)
	);

	bfr new_net_3777_bfr_after (
		.din(_0614_),
		.dout(new_net_3777)
	);

	bfr new_net_3778_bfr_after (
		.din(new_net_3777),
		.dout(new_net_3778)
	);

	bfr new_net_3779_bfr_before (
		.din(new_net_3779),
		.dout(new_net_131)
	);

	bfr new_net_3780_bfr_before (
		.din(new_net_3780),
		.dout(new_net_3779)
	);

	spl4L _0614__v_fanout (
		.a(new_net_3778),
		.b(new_net_133),
		.c(new_net_132),
		.d(new_net_134),
		.e(new_net_3780)
	);

	spl4L new_net_1804_v_fanout (
		.a(new_net_1804),
		.b(new_net_1008),
		.c(new_net_1004),
		.d(new_net_1003),
		.e(new_net_1010)
	);

	bfr new_net_3781_bfr_before (
		.din(new_net_3781),
		.dout(G5218)
	);

	bfr new_net_3782_bfr_before (
		.din(new_net_3782),
		.dout(new_net_3781)
	);

	bfr new_net_3783_bfr_before (
		.din(new_net_3783),
		.dout(new_net_3782)
	);

	bfr new_net_3784_bfr_before (
		.din(new_net_3784),
		.dout(new_net_3783)
	);

	bfr new_net_3785_bfr_before (
		.din(new_net_3785),
		.dout(new_net_3784)
	);

	bfr new_net_3786_bfr_before (
		.din(new_net_3786),
		.dout(new_net_3785)
	);

	bfr new_net_3787_bfr_before (
		.din(new_net_3787),
		.dout(new_net_3786)
	);

	bfr new_net_3788_bfr_before (
		.din(new_net_3788),
		.dout(new_net_3787)
	);

	bfr new_net_3789_bfr_before (
		.din(new_net_3789),
		.dout(new_net_3788)
	);

	bfr new_net_3790_bfr_before (
		.din(new_net_3790),
		.dout(new_net_3789)
	);

	bfr new_net_3791_bfr_before (
		.din(new_net_3791),
		.dout(new_net_3790)
	);

	bfr new_net_3792_bfr_before (
		.din(new_net_3792),
		.dout(new_net_3791)
	);

	bfr new_net_3793_bfr_before (
		.din(new_net_3793),
		.dout(new_net_3792)
	);

	bfr new_net_3794_bfr_before (
		.din(new_net_3794),
		.dout(new_net_3793)
	);

	bfr new_net_3795_bfr_before (
		.din(new_net_3795),
		.dout(new_net_3794)
	);

	bfr new_net_3796_bfr_before (
		.din(new_net_3796),
		.dout(new_net_3795)
	);

	bfr new_net_3797_bfr_before (
		.din(new_net_3797),
		.dout(new_net_3796)
	);

	bfr new_net_3798_bfr_before (
		.din(new_net_3798),
		.dout(new_net_3797)
	);

	bfr new_net_3799_bfr_before (
		.din(new_net_3799),
		.dout(new_net_3798)
	);

	bfr new_net_3800_bfr_before (
		.din(new_net_3800),
		.dout(new_net_3799)
	);

	bfr new_net_3801_bfr_before (
		.din(new_net_3801),
		.dout(new_net_3800)
	);

	bfr new_net_3802_bfr_before (
		.din(new_net_3802),
		.dout(new_net_3801)
	);

	bfr new_net_3803_bfr_before (
		.din(new_net_3803),
		.dout(new_net_3802)
	);

	bfr new_net_3804_bfr_before (
		.din(new_net_3804),
		.dout(new_net_3803)
	);

	bfr new_net_3805_bfr_before (
		.din(new_net_3805),
		.dout(new_net_3804)
	);

	bfr new_net_3806_bfr_before (
		.din(new_net_3806),
		.dout(new_net_3805)
	);

	bfr new_net_3807_bfr_before (
		.din(new_net_3807),
		.dout(new_net_3806)
	);

	bfr new_net_3808_bfr_before (
		.din(new_net_3808),
		.dout(new_net_3807)
	);

	bfr new_net_3809_bfr_before (
		.din(new_net_3809),
		.dout(new_net_3808)
	);

	bfr new_net_3810_bfr_before (
		.din(new_net_3810),
		.dout(new_net_3809)
	);

	bfr new_net_3811_bfr_before (
		.din(new_net_3811),
		.dout(new_net_3810)
	);

	bfr new_net_3812_bfr_before (
		.din(new_net_3812),
		.dout(new_net_3811)
	);

	bfr new_net_3813_bfr_before (
		.din(new_net_3813),
		.dout(new_net_3812)
	);

	bfr new_net_3814_bfr_before (
		.din(new_net_3814),
		.dout(new_net_3813)
	);

	bfr new_net_3815_bfr_before (
		.din(new_net_3815),
		.dout(new_net_3814)
	);

	bfr new_net_3816_bfr_before (
		.din(new_net_3816),
		.dout(new_net_3815)
	);

	bfr new_net_3817_bfr_before (
		.din(new_net_3817),
		.dout(new_net_3816)
	);

	bfr new_net_3818_bfr_before (
		.din(new_net_3818),
		.dout(new_net_3817)
	);

	bfr new_net_3819_bfr_before (
		.din(new_net_3819),
		.dout(new_net_3818)
	);

	spl2 new_net_1878_v_fanout (
		.a(new_net_1878),
		.b(new_net_1337),
		.c(new_net_3819)
	);

	spl2 new_net_1883_v_fanout (
		.a(new_net_1883),
		.b(new_net_457),
		.c(new_net_459)
	);

	spl4L new_net_1884_v_fanout (
		.a(new_net_1884),
		.b(new_net_463),
		.c(new_net_464),
		.d(new_net_462),
		.e(new_net_456)
	);

	bfr new_net_3820_bfr_after (
		.din(new_net_2),
		.dout(new_net_3820)
	);

	bfr new_net_3821_bfr_after (
		.din(new_net_3820),
		.dout(new_net_3821)
	);

	bfr new_net_3822_bfr_before (
		.din(new_net_3822),
		.dout(G5203)
	);

	bfr new_net_3823_bfr_before (
		.din(new_net_3823),
		.dout(new_net_3822)
	);

	bfr new_net_3824_bfr_before (
		.din(new_net_3824),
		.dout(new_net_3823)
	);

	bfr new_net_3825_bfr_before (
		.din(new_net_3825),
		.dout(new_net_3824)
	);

	bfr new_net_3826_bfr_before (
		.din(new_net_3826),
		.dout(new_net_3825)
	);

	bfr new_net_3827_bfr_before (
		.din(new_net_3827),
		.dout(new_net_3826)
	);

	bfr new_net_3828_bfr_before (
		.din(new_net_3828),
		.dout(new_net_3827)
	);

	bfr new_net_3829_bfr_before (
		.din(new_net_3829),
		.dout(new_net_3828)
	);

	bfr new_net_3830_bfr_before (
		.din(new_net_3830),
		.dout(new_net_3829)
	);

	bfr new_net_3831_bfr_before (
		.din(new_net_3831),
		.dout(new_net_3830)
	);

	bfr new_net_3832_bfr_before (
		.din(new_net_3832),
		.dout(new_net_3831)
	);

	bfr new_net_3833_bfr_before (
		.din(new_net_3833),
		.dout(new_net_3832)
	);

	bfr new_net_3834_bfr_before (
		.din(new_net_3834),
		.dout(new_net_3833)
	);

	bfr new_net_3835_bfr_before (
		.din(new_net_3835),
		.dout(new_net_3834)
	);

	bfr new_net_3836_bfr_before (
		.din(new_net_3836),
		.dout(new_net_3835)
	);

	bfr new_net_3837_bfr_before (
		.din(new_net_3837),
		.dout(new_net_3836)
	);

	bfr new_net_3838_bfr_before (
		.din(new_net_3838),
		.dout(new_net_3837)
	);

	bfr new_net_3839_bfr_before (
		.din(new_net_3839),
		.dout(new_net_3838)
	);

	bfr new_net_3840_bfr_before (
		.din(new_net_3840),
		.dout(new_net_3839)
	);

	bfr new_net_3841_bfr_before (
		.din(new_net_3841),
		.dout(new_net_3840)
	);

	bfr new_net_3842_bfr_before (
		.din(new_net_3842),
		.dout(new_net_3841)
	);

	bfr new_net_3843_bfr_before (
		.din(new_net_3843),
		.dout(new_net_3842)
	);

	bfr new_net_3844_bfr_before (
		.din(new_net_3844),
		.dout(new_net_3843)
	);

	bfr new_net_3845_bfr_before (
		.din(new_net_3845),
		.dout(new_net_3844)
	);

	bfr new_net_3846_bfr_before (
		.din(new_net_3846),
		.dout(new_net_3845)
	);

	bfr new_net_3847_bfr_before (
		.din(new_net_3847),
		.dout(new_net_3846)
	);

	bfr new_net_3848_bfr_before (
		.din(new_net_3848),
		.dout(new_net_3847)
	);

	bfr new_net_3849_bfr_before (
		.din(new_net_3849),
		.dout(new_net_3848)
	);

	bfr new_net_3850_bfr_before (
		.din(new_net_3850),
		.dout(new_net_3849)
	);

	bfr new_net_3851_bfr_before (
		.din(new_net_3851),
		.dout(new_net_3850)
	);

	bfr new_net_3852_bfr_before (
		.din(new_net_3852),
		.dout(new_net_3851)
	);

	bfr new_net_3853_bfr_before (
		.din(new_net_3853),
		.dout(new_net_3852)
	);

	bfr new_net_3854_bfr_before (
		.din(new_net_3854),
		.dout(new_net_3853)
	);

	bfr new_net_3855_bfr_before (
		.din(new_net_3855),
		.dout(new_net_3854)
	);

	bfr new_net_3856_bfr_before (
		.din(new_net_3856),
		.dout(new_net_3855)
	);

	bfr new_net_3857_bfr_before (
		.din(new_net_3857),
		.dout(new_net_3856)
	);

	bfr new_net_3858_bfr_before (
		.din(new_net_3858),
		.dout(new_net_3857)
	);

	spl2 new_net_2_v_fanout (
		.a(new_net_3821),
		.b(new_net_3858),
		.c(new_net_1621)
	);

	spl3L new_net_1885_v_fanout (
		.a(new_net_1885),
		.b(new_net_465),
		.c(new_net_466),
		.d(new_net_458)
	);

	bfr new_net_3859_bfr_after (
		.din(_1046_),
		.dout(new_net_3859)
	);

	bfr new_net_3860_bfr_after (
		.din(new_net_3859),
		.dout(new_net_3860)
	);

	bfr new_net_3861_bfr_after (
		.din(new_net_3860),
		.dout(new_net_3861)
	);

	bfr new_net_3862_bfr_after (
		.din(new_net_3861),
		.dout(new_net_3862)
	);

	bfr new_net_3863_bfr_after (
		.din(new_net_3862),
		.dout(new_net_3863)
	);

	bfr new_net_3864_bfr_after (
		.din(new_net_3863),
		.dout(new_net_3864)
	);

	bfr new_net_3865_bfr_after (
		.din(new_net_3864),
		.dout(new_net_3865)
	);

	bfr new_net_3866_bfr_after (
		.din(new_net_3865),
		.dout(new_net_3866)
	);

	bfr new_net_3867_bfr_after (
		.din(new_net_3866),
		.dout(new_net_3867)
	);

	bfr new_net_3868_bfr_after (
		.din(new_net_3867),
		.dout(new_net_3868)
	);

	bfr new_net_3869_bfr_after (
		.din(new_net_3868),
		.dout(new_net_3869)
	);

	bfr new_net_3870_bfr_after (
		.din(new_net_3869),
		.dout(new_net_3870)
	);

	bfr new_net_3871_bfr_after (
		.din(new_net_3870),
		.dout(new_net_3871)
	);

	bfr new_net_3872_bfr_after (
		.din(new_net_3871),
		.dout(new_net_3872)
	);

	bfr new_net_3873_bfr_after (
		.din(new_net_3872),
		.dout(new_net_3873)
	);

	bfr new_net_3874_bfr_after (
		.din(new_net_3873),
		.dout(new_net_3874)
	);

	bfr new_net_3875_bfr_after (
		.din(new_net_3874),
		.dout(new_net_3875)
	);

	bfr new_net_3876_bfr_after (
		.din(new_net_3875),
		.dout(new_net_3876)
	);

	bfr new_net_3877_bfr_after (
		.din(new_net_3876),
		.dout(new_net_3877)
	);

	bfr new_net_3878_bfr_after (
		.din(new_net_3877),
		.dout(new_net_3878)
	);

	bfr new_net_3879_bfr_after (
		.din(new_net_3878),
		.dout(new_net_3879)
	);

	bfr new_net_3880_bfr_after (
		.din(new_net_3879),
		.dout(new_net_3880)
	);

	bfr new_net_3881_bfr_after (
		.din(new_net_3880),
		.dout(new_net_3881)
	);

	bfr new_net_3882_bfr_after (
		.din(new_net_3881),
		.dout(new_net_3882)
	);

	bfr new_net_3883_bfr_after (
		.din(new_net_3882),
		.dout(new_net_3883)
	);

	bfr new_net_3884_bfr_after (
		.din(new_net_3883),
		.dout(new_net_3884)
	);

	bfr new_net_3885_bfr_after (
		.din(new_net_3884),
		.dout(new_net_3885)
	);

	bfr new_net_3886_bfr_after (
		.din(new_net_3885),
		.dout(new_net_3886)
	);

	bfr new_net_3887_bfr_after (
		.din(new_net_3886),
		.dout(new_net_3887)
	);

	bfr new_net_3888_bfr_after (
		.din(new_net_3887),
		.dout(new_net_3888)
	);

	bfr new_net_3889_bfr_after (
		.din(new_net_3888),
		.dout(new_net_3889)
	);

	bfr new_net_3890_bfr_after (
		.din(new_net_3889),
		.dout(new_net_3890)
	);

	bfr new_net_3891_bfr_after (
		.din(new_net_3890),
		.dout(new_net_3891)
	);

	bfr new_net_3892_bfr_after (
		.din(new_net_3891),
		.dout(new_net_3892)
	);

	bfr new_net_3893_bfr_after (
		.din(new_net_3892),
		.dout(new_net_3893)
	);

	bfr new_net_3894_bfr_after (
		.din(new_net_3893),
		.dout(new_net_3894)
	);

	bfr new_net_3895_bfr_after (
		.din(new_net_3894),
		.dout(new_net_3895)
	);

	spl2 _1046__v_fanout (
		.a(new_net_3895),
		.b(new_net_1129),
		.c(new_net_1130)
	);

	spl2 new_net_1808_v_fanout (
		.a(new_net_1808),
		.b(new_net_1068),
		.c(new_net_1072)
	);

	spl2 new_net_1771_v_fanout (
		.a(new_net_1771),
		.b(new_net_978),
		.c(new_net_985)
	);

	bfr new_net_3896_bfr_after (
		.din(_0943_),
		.dout(new_net_3896)
	);

	bfr new_net_3897_bfr_after (
		.din(new_net_3896),
		.dout(new_net_3897)
	);

	bfr new_net_3898_bfr_before (
		.din(new_net_3898),
		.dout(new_net_1628)
	);

	spl3L _0943__v_fanout (
		.a(new_net_3897),
		.b(new_net_3898),
		.c(new_net_1630),
		.d(new_net_1629)
	);

	spl4L new_net_1873_v_fanout (
		.a(new_net_1873),
		.b(new_net_1380),
		.c(new_net_1375),
		.d(new_net_1377),
		.e(new_net_1378)
	);

	spl3L _0105__v_fanout (
		.a(_0105_),
		.b(new_net_1925),
		.c(new_net_1923),
		.d(new_net_1924)
	);

	spl4L new_net_1809_v_fanout (
		.a(new_net_1809),
		.b(new_net_1076),
		.c(new_net_1074),
		.d(new_net_1067),
		.e(new_net_1070)
	);

	bfr new_net_3899_bfr_after (
		.din(_0252_),
		.dout(new_net_3899)
	);

	bfr new_net_3900_bfr_after (
		.din(new_net_3899),
		.dout(new_net_3900)
	);

	bfr new_net_3901_bfr_after (
		.din(new_net_3900),
		.dout(new_net_3901)
	);

	bfr new_net_3902_bfr_after (
		.din(new_net_3901),
		.dout(new_net_3902)
	);

	bfr new_net_3903_bfr_after (
		.din(new_net_3902),
		.dout(new_net_3903)
	);

	bfr new_net_3904_bfr_after (
		.din(new_net_3903),
		.dout(new_net_3904)
	);

	bfr new_net_3905_bfr_after (
		.din(new_net_3904),
		.dout(new_net_3905)
	);

	bfr new_net_3906_bfr_after (
		.din(new_net_3905),
		.dout(new_net_3906)
	);

	bfr new_net_3907_bfr_after (
		.din(new_net_3906),
		.dout(new_net_3907)
	);

	bfr new_net_3908_bfr_after (
		.din(new_net_3907),
		.dout(new_net_3908)
	);

	bfr new_net_3909_bfr_after (
		.din(new_net_3908),
		.dout(new_net_3909)
	);

	bfr new_net_3910_bfr_after (
		.din(new_net_3909),
		.dout(new_net_3910)
	);

	bfr new_net_3911_bfr_after (
		.din(new_net_3910),
		.dout(new_net_3911)
	);

	bfr new_net_3912_bfr_before (
		.din(new_net_3912),
		.dout(new_net_1926)
	);

	spl2 _0252__v_fanout (
		.a(new_net_3911),
		.b(new_net_432),
		.c(new_net_3912)
	);

	bfr new_net_3913_bfr_after (
		.din(_0949_),
		.dout(new_net_3913)
	);

	bfr new_net_3914_bfr_before (
		.din(new_net_3914),
		.dout(new_net_741)
	);

	bfr new_net_3915_bfr_before (
		.din(new_net_3915),
		.dout(new_net_3914)
	);

	spl4L _0949__v_fanout (
		.a(new_net_3913),
		.b(new_net_742),
		.c(new_net_744),
		.d(new_net_743),
		.e(new_net_3915)
	);

	spl4L new_net_1846_v_fanout (
		.a(new_net_1846),
		.b(new_net_1172),
		.c(new_net_1175),
		.d(new_net_1177),
		.e(new_net_1171)
	);

	spl2 new_net_0_v_fanout (
		.a(new_net_0),
		.b(new_net_1934),
		.c(new_net_1935)
	);

	spl4L new_net_1750_v_fanout (
		.a(new_net_1750),
		.b(new_net_1527),
		.c(new_net_1514),
		.d(new_net_1521),
		.e(new_net_1531)
	);

	bfr new_net_3916_bfr_before (
		.din(new_net_3916),
		.dout(G5199)
	);

	bfr new_net_3917_bfr_before (
		.din(new_net_3917),
		.dout(new_net_3916)
	);

	bfr new_net_3918_bfr_before (
		.din(new_net_3918),
		.dout(new_net_3917)
	);

	bfr new_net_3919_bfr_before (
		.din(new_net_3919),
		.dout(new_net_3918)
	);

	bfr new_net_3920_bfr_before (
		.din(new_net_3920),
		.dout(new_net_3919)
	);

	bfr new_net_3921_bfr_before (
		.din(new_net_3921),
		.dout(new_net_3920)
	);

	bfr new_net_3922_bfr_before (
		.din(new_net_3922),
		.dout(new_net_3921)
	);

	bfr new_net_3923_bfr_before (
		.din(new_net_3923),
		.dout(new_net_3922)
	);

	bfr new_net_3924_bfr_before (
		.din(new_net_3924),
		.dout(new_net_3923)
	);

	bfr new_net_3925_bfr_before (
		.din(new_net_3925),
		.dout(new_net_3924)
	);

	bfr new_net_3926_bfr_before (
		.din(new_net_3926),
		.dout(new_net_3925)
	);

	bfr new_net_3927_bfr_before (
		.din(new_net_3927),
		.dout(new_net_3926)
	);

	bfr new_net_3928_bfr_before (
		.din(new_net_3928),
		.dout(new_net_3927)
	);

	bfr new_net_3929_bfr_before (
		.din(new_net_3929),
		.dout(new_net_3928)
	);

	bfr new_net_3930_bfr_before (
		.din(new_net_3930),
		.dout(new_net_3929)
	);

	bfr new_net_3931_bfr_before (
		.din(new_net_3931),
		.dout(new_net_3930)
	);

	bfr new_net_3932_bfr_before (
		.din(new_net_3932),
		.dout(new_net_3931)
	);

	bfr new_net_3933_bfr_before (
		.din(new_net_3933),
		.dout(new_net_3932)
	);

	bfr new_net_3934_bfr_before (
		.din(new_net_3934),
		.dout(new_net_3933)
	);

	bfr new_net_3935_bfr_before (
		.din(new_net_3935),
		.dout(new_net_3934)
	);

	bfr new_net_3936_bfr_before (
		.din(new_net_3936),
		.dout(new_net_3935)
	);

	bfr new_net_3937_bfr_before (
		.din(new_net_3937),
		.dout(new_net_3936)
	);

	bfr new_net_3938_bfr_before (
		.din(new_net_3938),
		.dout(new_net_3937)
	);

	bfr new_net_3939_bfr_before (
		.din(new_net_3939),
		.dout(new_net_3938)
	);

	bfr new_net_3940_bfr_before (
		.din(new_net_3940),
		.dout(new_net_3939)
	);

	bfr new_net_3941_bfr_before (
		.din(new_net_3941),
		.dout(new_net_3940)
	);

	bfr new_net_3942_bfr_before (
		.din(new_net_3942),
		.dout(new_net_3941)
	);

	bfr new_net_3943_bfr_before (
		.din(new_net_3943),
		.dout(new_net_3942)
	);

	bfr new_net_3944_bfr_before (
		.din(new_net_3944),
		.dout(new_net_3943)
	);

	bfr new_net_3945_bfr_before (
		.din(new_net_3945),
		.dout(new_net_3944)
	);

	bfr new_net_3946_bfr_before (
		.din(new_net_3946),
		.dout(new_net_3945)
	);

	bfr new_net_3947_bfr_before (
		.din(new_net_3947),
		.dout(new_net_3946)
	);

	bfr new_net_3948_bfr_before (
		.din(new_net_3948),
		.dout(new_net_3947)
	);

	bfr new_net_3949_bfr_before (
		.din(new_net_3949),
		.dout(new_net_3948)
	);

	bfr new_net_3950_bfr_before (
		.din(new_net_3950),
		.dout(new_net_3949)
	);

	bfr new_net_3951_bfr_before (
		.din(new_net_3951),
		.dout(new_net_3950)
	);

	bfr new_net_3952_bfr_before (
		.din(new_net_3952),
		.dout(new_net_3951)
	);

	bfr new_net_3953_bfr_before (
		.din(new_net_3953),
		.dout(new_net_3952)
	);

	bfr new_net_3954_bfr_before (
		.din(new_net_3954),
		.dout(new_net_3953)
	);

	spl2 new_net_14_v_fanout (
		.a(new_net_14),
		.b(new_net_3954),
		.c(new_net_860)
	);

	spl3L new_net_1749_v_fanout (
		.a(new_net_1749),
		.b(new_net_1522),
		.c(new_net_1515),
		.d(new_net_1520)
	);

	spl3L _0268__v_fanout (
		.a(_0268_),
		.b(new_net_1936),
		.c(new_net_1938),
		.d(new_net_1937)
	);

	bfr new_net_3955_bfr_after (
		.din(_0778_),
		.dout(new_net_3955)
	);

	bfr new_net_3956_bfr_after (
		.din(new_net_3955),
		.dout(new_net_3956)
	);

	spl4L _0778__v_fanout (
		.a(new_net_3956),
		.b(new_net_812),
		.c(new_net_813),
		.d(new_net_811),
		.e(new_net_810)
	);

	spl3L _0258__v_fanout (
		.a(_0258_),
		.b(new_net_1939),
		.c(new_net_1941),
		.d(new_net_1940)
	);

	spl4L new_net_1874_v_fanout (
		.a(new_net_1874),
		.b(new_net_1369),
		.c(new_net_1368),
		.d(new_net_1367),
		.e(new_net_1365)
	);

	bfr new_net_3957_bfr_after (
		.din(_0933_),
		.dout(new_net_3957)
	);

	bfr new_net_3958_bfr_after (
		.din(new_net_3957),
		.dout(new_net_3958)
	);

	bfr new_net_3959_bfr_before (
		.din(new_net_3959),
		.dout(new_net_1406)
	);

	bfr new_net_3960_bfr_before (
		.din(new_net_3960),
		.dout(new_net_3959)
	);

	spl2 _0933__v_fanout (
		.a(new_net_3958),
		.b(new_net_3960),
		.c(new_net_1407)
	);

	bfr new_net_3961_bfr_after (
		.din(new_net_25),
		.dout(new_net_3961)
	);

	bfr new_net_3962_bfr_after (
		.din(new_net_3961),
		.dout(new_net_3962)
	);

	bfr new_net_3963_bfr_after (
		.din(new_net_3962),
		.dout(new_net_3963)
	);

	bfr new_net_3964_bfr_after (
		.din(new_net_3963),
		.dout(new_net_3964)
	);

	bfr new_net_3965_bfr_after (
		.din(new_net_3964),
		.dout(new_net_3965)
	);

	bfr new_net_3966_bfr_after (
		.din(new_net_3965),
		.dout(new_net_3966)
	);

	bfr new_net_3967_bfr_after (
		.din(new_net_3966),
		.dout(new_net_3967)
	);

	bfr new_net_3968_bfr_after (
		.din(new_net_3967),
		.dout(new_net_3968)
	);

	bfr new_net_3969_bfr_after (
		.din(new_net_3968),
		.dout(new_net_3969)
	);

	bfr new_net_3970_bfr_after (
		.din(new_net_3969),
		.dout(new_net_3970)
	);

	bfr new_net_3971_bfr_after (
		.din(new_net_3970),
		.dout(new_net_3971)
	);

	bfr new_net_3972_bfr_after (
		.din(new_net_3971),
		.dout(new_net_3972)
	);

	bfr new_net_3973_bfr_after (
		.din(new_net_3972),
		.dout(new_net_3973)
	);

	bfr new_net_3974_bfr_after (
		.din(new_net_3973),
		.dout(new_net_3974)
	);

	bfr new_net_3975_bfr_after (
		.din(new_net_3974),
		.dout(new_net_3975)
	);

	bfr new_net_3976_bfr_after (
		.din(new_net_3975),
		.dout(new_net_3976)
	);

	bfr new_net_3977_bfr_after (
		.din(new_net_3976),
		.dout(new_net_3977)
	);

	bfr new_net_3978_bfr_after (
		.din(new_net_3977),
		.dout(new_net_3978)
	);

	bfr new_net_3979_bfr_after (
		.din(new_net_3978),
		.dout(new_net_3979)
	);

	bfr new_net_3980_bfr_after (
		.din(new_net_3979),
		.dout(new_net_3980)
	);

	bfr new_net_3981_bfr_after (
		.din(new_net_3980),
		.dout(new_net_3981)
	);

	bfr new_net_3982_bfr_after (
		.din(new_net_3981),
		.dout(new_net_3982)
	);

	bfr new_net_3983_bfr_after (
		.din(new_net_3982),
		.dout(new_net_3983)
	);

	bfr new_net_3984_bfr_after (
		.din(new_net_3983),
		.dout(new_net_3984)
	);

	bfr new_net_3985_bfr_after (
		.din(new_net_3984),
		.dout(new_net_3985)
	);

	bfr new_net_3986_bfr_after (
		.din(new_net_3985),
		.dout(new_net_3986)
	);

	bfr new_net_3987_bfr_after (
		.din(new_net_3986),
		.dout(new_net_3987)
	);

	bfr new_net_3988_bfr_after (
		.din(new_net_3987),
		.dout(new_net_3988)
	);

	bfr new_net_3989_bfr_after (
		.din(new_net_3988),
		.dout(new_net_3989)
	);

	bfr new_net_3990_bfr_after (
		.din(new_net_3989),
		.dout(new_net_3990)
	);

	bfr new_net_3991_bfr_after (
		.din(new_net_3990),
		.dout(new_net_3991)
	);

	bfr new_net_3992_bfr_after (
		.din(new_net_3991),
		.dout(new_net_3992)
	);

	bfr new_net_3993_bfr_after (
		.din(new_net_3992),
		.dout(new_net_3993)
	);

	bfr new_net_3994_bfr_after (
		.din(new_net_3993),
		.dout(new_net_3994)
	);

	bfr new_net_3995_bfr_after (
		.din(new_net_3994),
		.dout(new_net_3995)
	);

	bfr new_net_3996_bfr_after (
		.din(new_net_3995),
		.dout(new_net_3996)
	);

	bfr new_net_3997_bfr_after (
		.din(new_net_3996),
		.dout(new_net_3997)
	);

	bfr new_net_3998_bfr_after (
		.din(new_net_3997),
		.dout(new_net_3998)
	);

	bfr new_net_3999_bfr_after (
		.din(new_net_3998),
		.dout(new_net_3999)
	);

	spl4L new_net_25_v_fanout (
		.a(new_net_3999),
		.b(G5225),
		.c(G5224),
		.d(G5223),
		.e(G5222)
	);

	bfr new_net_4000_bfr_after (
		.din(_0097_),
		.dout(new_net_4000)
	);

	bfr new_net_4001_bfr_after (
		.din(new_net_4000),
		.dout(new_net_4001)
	);

	bfr new_net_4002_bfr_after (
		.din(new_net_4001),
		.dout(new_net_4002)
	);

	bfr new_net_4003_bfr_after (
		.din(new_net_4002),
		.dout(new_net_4003)
	);

	bfr new_net_4004_bfr_after (
		.din(new_net_4003),
		.dout(new_net_4004)
	);

	bfr new_net_4005_bfr_after (
		.din(new_net_4004),
		.dout(new_net_4005)
	);

	bfr new_net_4006_bfr_after (
		.din(new_net_4005),
		.dout(new_net_4006)
	);

	bfr new_net_4007_bfr_after (
		.din(new_net_4006),
		.dout(new_net_4007)
	);

	bfr new_net_4008_bfr_after (
		.din(new_net_4007),
		.dout(new_net_4008)
	);

	bfr new_net_4009_bfr_after (
		.din(new_net_4008),
		.dout(new_net_4009)
	);

	bfr new_net_4010_bfr_after (
		.din(new_net_4009),
		.dout(new_net_4010)
	);

	bfr new_net_4011_bfr_after (
		.din(new_net_4010),
		.dout(new_net_4011)
	);

	bfr new_net_4012_bfr_before (
		.din(new_net_4012),
		.dout(new_net_1942)
	);

	spl2 _0097__v_fanout (
		.a(new_net_4011),
		.b(new_net_1148),
		.c(new_net_4012)
	);

	spl3L _0256__v_fanout (
		.a(_0256_),
		.b(new_net_1949),
		.c(new_net_1950),
		.d(new_net_1951)
	);

	spl4L new_net_1847_v_fanout (
		.a(new_net_1847),
		.b(new_net_1173),
		.c(new_net_1179),
		.d(new_net_1174),
		.e(new_net_1169)
	);

	bfr new_net_4013_bfr_after (
		.din(_0800_),
		.dout(new_net_4013)
	);

	bfr new_net_4014_bfr_after (
		.din(new_net_4013),
		.dout(new_net_4014)
	);

	spl3L _0800__v_fanout (
		.a(new_net_4014),
		.b(new_net_1299),
		.c(new_net_1301),
		.d(new_net_1300)
	);

	bfr new_net_4015_bfr_after (
		.din(_0262_),
		.dout(new_net_4015)
	);

	bfr new_net_4016_bfr_after (
		.din(new_net_4015),
		.dout(new_net_4016)
	);

	bfr new_net_4017_bfr_after (
		.din(new_net_4016),
		.dout(new_net_4017)
	);

	bfr new_net_4018_bfr_after (
		.din(new_net_4017),
		.dout(new_net_4018)
	);

	bfr new_net_4019_bfr_after (
		.din(new_net_4018),
		.dout(new_net_4019)
	);

	bfr new_net_4020_bfr_after (
		.din(new_net_4019),
		.dout(new_net_4020)
	);

	bfr new_net_4021_bfr_after (
		.din(new_net_4020),
		.dout(new_net_4021)
	);

	bfr new_net_4022_bfr_after (
		.din(new_net_4021),
		.dout(new_net_4022)
	);

	bfr new_net_4023_bfr_after (
		.din(new_net_4022),
		.dout(new_net_4023)
	);

	bfr new_net_4024_bfr_after (
		.din(new_net_4023),
		.dout(new_net_4024)
	);

	bfr new_net_4025_bfr_after (
		.din(new_net_4024),
		.dout(new_net_4025)
	);

	bfr new_net_4026_bfr_after (
		.din(new_net_4025),
		.dout(new_net_4026)
	);

	bfr new_net_4027_bfr_after (
		.din(new_net_4026),
		.dout(new_net_4027)
	);

	bfr new_net_4028_bfr_before (
		.din(new_net_4028),
		.dout(new_net_1952)
	);

	spl2 _0262__v_fanout (
		.a(new_net_4027),
		.b(new_net_1357),
		.c(new_net_4028)
	);

	spl4L new_net_1826_v_fanout (
		.a(new_net_1826),
		.b(new_net_1549),
		.c(new_net_1556),
		.d(new_net_1555),
		.e(new_net_1548)
	);

	spl3L new_net_1869_v_fanout (
		.a(new_net_1869),
		.b(new_net_1656),
		.c(new_net_1658),
		.d(new_net_1663)
	);

	spl2 new_net_1836_v_fanout (
		.a(new_net_1836),
		.b(new_net_752),
		.c(new_net_755)
	);

	spl4L new_net_1843_v_fanout (
		.a(new_net_1843),
		.b(new_net_1050),
		.c(new_net_1051),
		.d(new_net_1049),
		.e(new_net_1045)
	);

	bfr new_net_4029_bfr_after (
		.din(_0099_),
		.dout(new_net_4029)
	);

	bfr new_net_4030_bfr_after (
		.din(new_net_4029),
		.dout(new_net_4030)
	);

	bfr new_net_4031_bfr_after (
		.din(new_net_4030),
		.dout(new_net_4031)
	);

	bfr new_net_4032_bfr_after (
		.din(new_net_4031),
		.dout(new_net_4032)
	);

	bfr new_net_4033_bfr_after (
		.din(new_net_4032),
		.dout(new_net_4033)
	);

	bfr new_net_4034_bfr_after (
		.din(new_net_4033),
		.dout(new_net_4034)
	);

	bfr new_net_4035_bfr_after (
		.din(new_net_4034),
		.dout(new_net_4035)
	);

	bfr new_net_4036_bfr_after (
		.din(new_net_4035),
		.dout(new_net_4036)
	);

	bfr new_net_4037_bfr_after (
		.din(new_net_4036),
		.dout(new_net_4037)
	);

	bfr new_net_4038_bfr_after (
		.din(new_net_4037),
		.dout(new_net_4038)
	);

	bfr new_net_4039_bfr_after (
		.din(new_net_4038),
		.dout(new_net_4039)
	);

	bfr new_net_4040_bfr_after (
		.din(new_net_4039),
		.dout(new_net_4040)
	);

	bfr new_net_4041_bfr_after (
		.din(new_net_4040),
		.dout(new_net_4041)
	);

	bfr new_net_4042_bfr_before (
		.din(new_net_4042),
		.dout(new_net_1959)
	);

	spl2 _0099__v_fanout (
		.a(new_net_4041),
		.b(new_net_4042),
		.c(new_net_677)
	);

	spl4L new_net_1875_v_fanout (
		.a(new_net_1875),
		.b(new_net_1373),
		.c(new_net_1376),
		.d(new_net_1370),
		.e(new_net_1366)
	);

	bfr new_net_4043_bfr_before (
		.din(new_net_4043),
		.dout(new_net_1513)
	);

	spl4L new_net_1753_v_fanout (
		.a(new_net_1753),
		.b(new_net_1518),
		.c(new_net_1524),
		.d(new_net_1517),
		.e(new_net_4043)
	);

	bfr new_net_4044_bfr_after (
		.din(_1228_),
		.dout(new_net_4044)
	);

	bfr new_net_4045_bfr_after (
		.din(new_net_4044),
		.dout(new_net_4045)
	);

	bfr new_net_4046_bfr_after (
		.din(new_net_4045),
		.dout(new_net_4046)
	);

	bfr new_net_4047_bfr_after (
		.din(new_net_4046),
		.dout(new_net_4047)
	);

	bfr new_net_4048_bfr_after (
		.din(new_net_4047),
		.dout(new_net_4048)
	);

	bfr new_net_4049_bfr_after (
		.din(new_net_4048),
		.dout(new_net_4049)
	);

	bfr new_net_4050_bfr_after (
		.din(new_net_4049),
		.dout(new_net_4050)
	);

	bfr new_net_4051_bfr_after (
		.din(new_net_4050),
		.dout(new_net_4051)
	);

	bfr new_net_4052_bfr_after (
		.din(new_net_4051),
		.dout(new_net_4052)
	);

	bfr new_net_4053_bfr_after (
		.din(new_net_4052),
		.dout(new_net_4053)
	);

	bfr new_net_4054_bfr_after (
		.din(new_net_4053),
		.dout(new_net_4054)
	);

	bfr new_net_4055_bfr_after (
		.din(new_net_4054),
		.dout(new_net_4055)
	);

	bfr new_net_4056_bfr_after (
		.din(new_net_4055),
		.dout(new_net_4056)
	);

	bfr new_net_4057_bfr_before (
		.din(new_net_4057),
		.dout(new_net_1967)
	);

	spl2 _1228__v_fanout (
		.a(new_net_4056),
		.b(new_net_801),
		.c(new_net_4057)
	);

	bfr new_net_4058_bfr_after (
		.din(_0937_),
		.dout(new_net_4058)
	);

	bfr new_net_4059_bfr_after (
		.din(new_net_4058),
		.dout(new_net_4059)
	);

	bfr new_net_4060_bfr_before (
		.din(new_net_4060),
		.dout(new_net_1060)
	);

	spl4L _0937__v_fanout (
		.a(new_net_4059),
		.b(new_net_1062),
		.c(new_net_1061),
		.d(new_net_1063),
		.e(new_net_4060)
	);

	spl3L new_net_1837_v_fanout (
		.a(new_net_1837),
		.b(new_net_749),
		.c(new_net_757),
		.d(new_net_751)
	);

	bfr new_net_4061_bfr_after (
		.din(_0250_),
		.dout(new_net_4061)
	);

	bfr new_net_4062_bfr_after (
		.din(new_net_4061),
		.dout(new_net_4062)
	);

	bfr new_net_4063_bfr_after (
		.din(new_net_4062),
		.dout(new_net_4063)
	);

	bfr new_net_4064_bfr_after (
		.din(new_net_4063),
		.dout(new_net_4064)
	);

	bfr new_net_4065_bfr_after (
		.din(new_net_4064),
		.dout(new_net_4065)
	);

	bfr new_net_4066_bfr_after (
		.din(new_net_4065),
		.dout(new_net_4066)
	);

	bfr new_net_4067_bfr_after (
		.din(new_net_4066),
		.dout(new_net_4067)
	);

	bfr new_net_4068_bfr_after (
		.din(new_net_4067),
		.dout(new_net_4068)
	);

	bfr new_net_4069_bfr_after (
		.din(new_net_4068),
		.dout(new_net_4069)
	);

	bfr new_net_4070_bfr_after (
		.din(new_net_4069),
		.dout(new_net_4070)
	);

	bfr new_net_4071_bfr_after (
		.din(new_net_4070),
		.dout(new_net_4071)
	);

	bfr new_net_4072_bfr_after (
		.din(new_net_4071),
		.dout(new_net_4072)
	);

	bfr new_net_4073_bfr_before (
		.din(new_net_4073),
		.dout(new_net_1974)
	);

	spl2 _0250__v_fanout (
		.a(new_net_4072),
		.b(new_net_384),
		.c(new_net_4073)
	);

	bfr new_net_4074_bfr_after (
		.din(_1076_),
		.dout(new_net_4074)
	);

	bfr new_net_4075_bfr_after (
		.din(new_net_4074),
		.dout(new_net_4075)
	);

	bfr new_net_4076_bfr_after (
		.din(new_net_4075),
		.dout(new_net_4076)
	);

	bfr new_net_4077_bfr_after (
		.din(new_net_4076),
		.dout(new_net_4077)
	);

	bfr new_net_4078_bfr_after (
		.din(new_net_4077),
		.dout(new_net_4078)
	);

	bfr new_net_4079_bfr_after (
		.din(new_net_4078),
		.dout(new_net_4079)
	);

	bfr new_net_4080_bfr_after (
		.din(new_net_4079),
		.dout(new_net_4080)
	);

	bfr new_net_4081_bfr_after (
		.din(new_net_4080),
		.dout(new_net_4081)
	);

	bfr new_net_4082_bfr_after (
		.din(new_net_4081),
		.dout(new_net_4082)
	);

	bfr new_net_4083_bfr_after (
		.din(new_net_4082),
		.dout(new_net_4083)
	);

	bfr new_net_4084_bfr_after (
		.din(new_net_4083),
		.dout(new_net_4084)
	);

	bfr new_net_4085_bfr_after (
		.din(new_net_4084),
		.dout(new_net_4085)
	);

	bfr new_net_4086_bfr_after (
		.din(new_net_4085),
		.dout(new_net_4086)
	);

	bfr new_net_4087_bfr_after (
		.din(new_net_4086),
		.dout(new_net_4087)
	);

	bfr new_net_4088_bfr_after (
		.din(new_net_4087),
		.dout(new_net_4088)
	);

	bfr new_net_4089_bfr_after (
		.din(new_net_4088),
		.dout(new_net_4089)
	);

	bfr new_net_4090_bfr_after (
		.din(new_net_4089),
		.dout(new_net_4090)
	);

	bfr new_net_4091_bfr_after (
		.din(new_net_4090),
		.dout(new_net_4091)
	);

	bfr new_net_4092_bfr_after (
		.din(new_net_4091),
		.dout(new_net_4092)
	);

	bfr new_net_4093_bfr_before (
		.din(new_net_4093),
		.dout(new_net_1282)
	);

	bfr new_net_4094_bfr_before (
		.din(new_net_4094),
		.dout(new_net_1284)
	);

	spl3L _1076__v_fanout (
		.a(new_net_4092),
		.b(new_net_4093),
		.c(new_net_1283),
		.d(new_net_4094)
	);

	spl4L new_net_1851_v_fanout (
		.a(new_net_1851),
		.b(new_net_1669),
		.c(new_net_1670),
		.d(new_net_1667),
		.e(new_net_1677)
	);

	bfr new_net_4095_bfr_after (
		.din(_0821_),
		.dout(new_net_4095)
	);

	bfr new_net_4096_bfr_after (
		.din(new_net_4095),
		.dout(new_net_4096)
	);

	spl4L _0821__v_fanout (
		.a(new_net_4096),
		.b(new_net_47),
		.c(new_net_49),
		.d(new_net_48),
		.e(new_net_46)
	);

	bfr new_net_4097_bfr_after (
		.din(new_net_26),
		.dout(new_net_4097)
	);

	bfr new_net_4098_bfr_after (
		.din(new_net_4097),
		.dout(new_net_4098)
	);

	bfr new_net_4099_bfr_after (
		.din(new_net_4098),
		.dout(new_net_4099)
	);

	bfr new_net_4100_bfr_after (
		.din(new_net_4099),
		.dout(new_net_4100)
	);

	bfr new_net_4101_bfr_after (
		.din(new_net_4100),
		.dout(new_net_4101)
	);

	bfr new_net_4102_bfr_after (
		.din(new_net_4101),
		.dout(new_net_4102)
	);

	bfr new_net_4103_bfr_after (
		.din(new_net_4102),
		.dout(new_net_4103)
	);

	bfr new_net_4104_bfr_after (
		.din(new_net_4103),
		.dout(new_net_4104)
	);

	bfr new_net_4105_bfr_after (
		.din(new_net_4104),
		.dout(new_net_4105)
	);

	bfr new_net_4106_bfr_after (
		.din(new_net_4105),
		.dout(new_net_4106)
	);

	bfr new_net_4107_bfr_after (
		.din(new_net_4106),
		.dout(new_net_4107)
	);

	bfr new_net_4108_bfr_after (
		.din(new_net_4107),
		.dout(new_net_4108)
	);

	bfr new_net_4109_bfr_after (
		.din(new_net_4108),
		.dout(new_net_4109)
	);

	bfr new_net_4110_bfr_after (
		.din(new_net_4109),
		.dout(new_net_4110)
	);

	bfr new_net_4111_bfr_after (
		.din(new_net_4110),
		.dout(new_net_4111)
	);

	bfr new_net_4112_bfr_after (
		.din(new_net_4111),
		.dout(new_net_4112)
	);

	bfr new_net_4113_bfr_after (
		.din(new_net_4112),
		.dout(new_net_4113)
	);

	bfr new_net_4114_bfr_after (
		.din(new_net_4113),
		.dout(new_net_4114)
	);

	bfr new_net_4115_bfr_after (
		.din(new_net_4114),
		.dout(new_net_4115)
	);

	bfr new_net_4116_bfr_after (
		.din(new_net_4115),
		.dout(new_net_4116)
	);

	bfr new_net_4117_bfr_after (
		.din(new_net_4116),
		.dout(new_net_4117)
	);

	bfr new_net_4118_bfr_after (
		.din(new_net_4117),
		.dout(new_net_4118)
	);

	bfr new_net_4119_bfr_after (
		.din(new_net_4118),
		.dout(new_net_4119)
	);

	bfr new_net_4120_bfr_after (
		.din(new_net_4119),
		.dout(new_net_4120)
	);

	bfr new_net_4121_bfr_after (
		.din(new_net_4120),
		.dout(new_net_4121)
	);

	bfr new_net_4122_bfr_after (
		.din(new_net_4121),
		.dout(new_net_4122)
	);

	bfr new_net_4123_bfr_after (
		.din(new_net_4122),
		.dout(new_net_4123)
	);

	bfr new_net_4124_bfr_after (
		.din(new_net_4123),
		.dout(new_net_4124)
	);

	bfr new_net_4125_bfr_after (
		.din(new_net_4124),
		.dout(new_net_4125)
	);

	bfr new_net_4126_bfr_after (
		.din(new_net_4125),
		.dout(new_net_4126)
	);

	bfr new_net_4127_bfr_after (
		.din(new_net_4126),
		.dout(new_net_4127)
	);

	bfr new_net_4128_bfr_after (
		.din(new_net_4127),
		.dout(new_net_4128)
	);

	bfr new_net_4129_bfr_after (
		.din(new_net_4128),
		.dout(new_net_4129)
	);

	bfr new_net_4130_bfr_after (
		.din(new_net_4129),
		.dout(new_net_4130)
	);

	bfr new_net_4131_bfr_after (
		.din(new_net_4130),
		.dout(new_net_4131)
	);

	bfr new_net_4132_bfr_after (
		.din(new_net_4131),
		.dout(new_net_4132)
	);

	bfr new_net_4133_bfr_after (
		.din(new_net_4132),
		.dout(new_net_4133)
	);

	bfr new_net_4134_bfr_after (
		.din(new_net_4133),
		.dout(new_net_4134)
	);

	bfr new_net_4135_bfr_after (
		.din(new_net_4134),
		.dout(new_net_4135)
	);

	spl2 new_net_26_v_fanout (
		.a(new_net_4135),
		.b(G5226),
		.c(G5227)
	);

	bfr new_net_4136_bfr_after (
		.din(_1047_),
		.dout(new_net_4136)
	);

	bfr new_net_4137_bfr_after (
		.din(new_net_4136),
		.dout(new_net_4137)
	);

	bfr new_net_4138_bfr_after (
		.din(new_net_4137),
		.dout(new_net_4138)
	);

	bfr new_net_4139_bfr_after (
		.din(new_net_4138),
		.dout(new_net_4139)
	);

	bfr new_net_4140_bfr_after (
		.din(new_net_4139),
		.dout(new_net_4140)
	);

	bfr new_net_4141_bfr_after (
		.din(new_net_4140),
		.dout(new_net_4141)
	);

	bfr new_net_4142_bfr_after (
		.din(new_net_4141),
		.dout(new_net_4142)
	);

	bfr new_net_4143_bfr_after (
		.din(new_net_4142),
		.dout(new_net_4143)
	);

	bfr new_net_4144_bfr_after (
		.din(new_net_4143),
		.dout(new_net_4144)
	);

	bfr new_net_4145_bfr_after (
		.din(new_net_4144),
		.dout(new_net_4145)
	);

	bfr new_net_4146_bfr_after (
		.din(new_net_4145),
		.dout(new_net_4146)
	);

	bfr new_net_4147_bfr_after (
		.din(new_net_4146),
		.dout(new_net_4147)
	);

	bfr new_net_4148_bfr_before (
		.din(new_net_4148),
		.dout(new_net_1982)
	);

	spl2 _1047__v_fanout (
		.a(new_net_4147),
		.b(new_net_1569),
		.c(new_net_4148)
	);

	bfr new_net_4149_bfr_before (
		.din(new_net_4149),
		.dout(new_net_1655)
	);

	spl4L new_net_1870_v_fanout (
		.a(new_net_1870),
		.b(new_net_1661),
		.c(new_net_1662),
		.d(new_net_1664),
		.e(new_net_4149)
	);

	spl3L _0091__v_fanout (
		.a(_0091_),
		.b(new_net_1990),
		.c(new_net_1989),
		.d(new_net_1991)
	);

	spl2 new_net_1813_v_fanout (
		.a(new_net_1813),
		.b(new_net_878),
		.c(new_net_881)
	);

	bfr new_net_4150_bfr_after (
		.din(_0897_),
		.dout(new_net_4150)
	);

	bfr new_net_4151_bfr_before (
		.din(new_net_4151),
		.dout(new_net_1992)
	);

	bfr new_net_4152_bfr_before (
		.din(new_net_4152),
		.dout(new_net_4151)
	);

	spl3L _0897__v_fanout (
		.a(new_net_4150),
		.b(new_net_4152),
		.c(new_net_346),
		.d(new_net_349)
	);

	bfr new_net_4153_bfr_after (
		.din(_0689_),
		.dout(new_net_4153)
	);

	bfr new_net_4154_bfr_after (
		.din(new_net_4153),
		.dout(new_net_4154)
	);

	spl3L _0689__v_fanout (
		.a(new_net_4154),
		.b(new_net_1594),
		.c(new_net_1595),
		.d(new_net_1596)
	);

	bfr new_net_4155_bfr_after (
		.din(_0663_),
		.dout(new_net_4155)
	);

	bfr new_net_4156_bfr_before (
		.din(new_net_4156),
		.dout(new_net_1993)
	);

	spl4L _0663__v_fanout (
		.a(new_net_4155),
		.b(new_net_1021),
		.c(new_net_1018),
		.d(new_net_4156),
		.e(new_net_1017)
	);

	bfr new_net_4157_bfr_before (
		.din(new_net_4157),
		.dout(new_net_1516)
	);

	spl4L new_net_1752_v_fanout (
		.a(new_net_1752),
		.b(new_net_1519),
		.c(new_net_4157),
		.d(new_net_1530),
		.e(new_net_1528)
	);

	bfr new_net_4158_bfr_after (
		.din(_0645_),
		.dout(new_net_4158)
	);

	bfr new_net_4159_bfr_after (
		.din(new_net_4158),
		.dout(new_net_4159)
	);

	spl4L _0645__v_fanout (
		.a(new_net_4159),
		.b(new_net_1291),
		.c(new_net_1293),
		.d(new_net_1292),
		.e(new_net_1290)
	);

	bfr new_net_4160_bfr_after (
		.din(_0740_),
		.dout(new_net_4160)
	);

	spl2 _0740__v_fanout (
		.a(new_net_4160),
		.b(new_net_1994),
		.c(new_net_1995)
	);

	bfr new_net_4161_bfr_after (
		.din(_0601_),
		.dout(new_net_4161)
	);

	bfr new_net_4162_bfr_after (
		.din(new_net_4161),
		.dout(new_net_4162)
	);

	bfr new_net_4163_bfr_after (
		.din(new_net_4162),
		.dout(new_net_4163)
	);

	spl4L _0601__v_fanout (
		.a(new_net_4163),
		.b(new_net_611),
		.c(new_net_614),
		.d(new_net_620),
		.e(new_net_1996)
	);

	spl3L _0103__v_fanout (
		.a(_0103_),
		.b(new_net_2005),
		.c(new_net_2004),
		.d(new_net_2003)
	);

	spl3L new_net_1765_v_fanout (
		.a(new_net_1765),
		.b(new_net_336),
		.c(new_net_343),
		.d(new_net_345)
	);

	spl4L new_net_1814_v_fanout (
		.a(new_net_1814),
		.b(new_net_874),
		.c(new_net_872),
		.d(new_net_879),
		.e(new_net_876)
	);

	spl2 new_net_1825_v_fanout (
		.a(new_net_1825),
		.b(new_net_1561),
		.c(new_net_1562)
	);

	spl3L new_net_1772_v_fanout (
		.a(new_net_1772),
		.b(new_net_994),
		.c(new_net_983),
		.d(new_net_993)
	);

	spl4L new_net_1842_v_fanout (
		.a(new_net_1842),
		.b(new_net_1043),
		.c(new_net_1038),
		.d(new_net_1040),
		.e(new_net_1041)
	);

	spl3L new_net_1779_v_fanout (
		.a(new_net_1779),
		.b(new_net_1246),
		.c(new_net_1249),
		.d(new_net_1245)
	);

	spl4L new_net_1751_v_fanout (
		.a(new_net_1751),
		.b(new_net_1526),
		.c(new_net_1525),
		.d(new_net_1529),
		.e(new_net_1523)
	);

	spl3L new_net_1755_v_fanout (
		.a(new_net_1755),
		.b(new_net_1752),
		.c(new_net_1749),
		.d(new_net_1750)
	);

	bfr new_net_4164_bfr_before (
		.din(new_net_4164),
		.dout(new_net_1251)
	);

	bfr new_net_4165_bfr_before (
		.din(new_net_4165),
		.dout(new_net_1252)
	);

	spl3L new_net_1782_v_fanout (
		.a(new_net_1782),
		.b(new_net_4164),
		.c(new_net_1253),
		.d(new_net_4165)
	);

	spl3L new_net_1810_v_fanout (
		.a(new_net_1810),
		.b(new_net_1069),
		.c(new_net_1073),
		.d(new_net_1075)
	);

	bfr new_net_4166_bfr_before (
		.din(new_net_4166),
		.dout(new_net_988)
	);

	spl4L new_net_1775_v_fanout (
		.a(new_net_1775),
		.b(new_net_992),
		.c(new_net_4166),
		.d(new_net_990),
		.e(new_net_1772)
	);

	spl3L new_net_1876_v_fanout (
		.a(new_net_1876),
		.b(new_net_1873),
		.c(new_net_1875),
		.d(new_net_1372)
	);

	spl4L new_net_1893_v_fanout (
		.a(new_net_1893),
		.b(new_net_1608),
		.c(new_net_1607),
		.d(new_net_1603),
		.e(new_net_1605)
	);

	spl4L new_net_1887_v_fanout (
		.a(new_net_1887),
		.b(new_net_1885),
		.c(new_net_1883),
		.d(new_net_467),
		.e(new_net_460)
	);

	bfr new_net_4167_bfr_after (
		.din(new_net_24),
		.dout(new_net_4167)
	);

	bfr new_net_4168_bfr_after (
		.din(new_net_4167),
		.dout(new_net_4168)
	);

	bfr new_net_4169_bfr_after (
		.din(new_net_4168),
		.dout(new_net_4169)
	);

	bfr new_net_4170_bfr_after (
		.din(new_net_4169),
		.dout(new_net_4170)
	);

	bfr new_net_4171_bfr_after (
		.din(new_net_4170),
		.dout(new_net_4171)
	);

	bfr new_net_4172_bfr_after (
		.din(new_net_4171),
		.dout(new_net_4172)
	);

	bfr new_net_4173_bfr_after (
		.din(new_net_4172),
		.dout(new_net_4173)
	);

	bfr new_net_4174_bfr_after (
		.din(new_net_4173),
		.dout(new_net_4174)
	);

	bfr new_net_4175_bfr_after (
		.din(new_net_4174),
		.dout(new_net_4175)
	);

	bfr new_net_4176_bfr_after (
		.din(new_net_4175),
		.dout(new_net_4176)
	);

	bfr new_net_4177_bfr_after (
		.din(new_net_4176),
		.dout(new_net_4177)
	);

	bfr new_net_4178_bfr_after (
		.din(new_net_4177),
		.dout(new_net_4178)
	);

	bfr new_net_4179_bfr_after (
		.din(new_net_4178),
		.dout(new_net_4179)
	);

	bfr new_net_4180_bfr_after (
		.din(new_net_4179),
		.dout(new_net_4180)
	);

	bfr new_net_4181_bfr_after (
		.din(new_net_4180),
		.dout(new_net_4181)
	);

	bfr new_net_4182_bfr_after (
		.din(new_net_4181),
		.dout(new_net_4182)
	);

	bfr new_net_4183_bfr_after (
		.din(new_net_4182),
		.dout(new_net_4183)
	);

	bfr new_net_4184_bfr_after (
		.din(new_net_4183),
		.dout(new_net_4184)
	);

	bfr new_net_4185_bfr_after (
		.din(new_net_4184),
		.dout(new_net_4185)
	);

	bfr new_net_4186_bfr_after (
		.din(new_net_4185),
		.dout(new_net_4186)
	);

	bfr new_net_4187_bfr_after (
		.din(new_net_4186),
		.dout(new_net_4187)
	);

	bfr new_net_4188_bfr_after (
		.din(new_net_4187),
		.dout(new_net_4188)
	);

	bfr new_net_4189_bfr_after (
		.din(new_net_4188),
		.dout(new_net_4189)
	);

	bfr new_net_4190_bfr_after (
		.din(new_net_4189),
		.dout(new_net_4190)
	);

	bfr new_net_4191_bfr_after (
		.din(new_net_4190),
		.dout(new_net_4191)
	);

	bfr new_net_4192_bfr_after (
		.din(new_net_4191),
		.dout(new_net_4192)
	);

	bfr new_net_4193_bfr_after (
		.din(new_net_4192),
		.dout(new_net_4193)
	);

	bfr new_net_4194_bfr_after (
		.din(new_net_4193),
		.dout(new_net_4194)
	);

	bfr new_net_4195_bfr_after (
		.din(new_net_4194),
		.dout(new_net_4195)
	);

	bfr new_net_4196_bfr_after (
		.din(new_net_4195),
		.dout(new_net_4196)
	);

	bfr new_net_4197_bfr_after (
		.din(new_net_4196),
		.dout(new_net_4197)
	);

	bfr new_net_4198_bfr_after (
		.din(new_net_4197),
		.dout(new_net_4198)
	);

	bfr new_net_4199_bfr_after (
		.din(new_net_4198),
		.dout(new_net_4199)
	);

	bfr new_net_4200_bfr_after (
		.din(new_net_4199),
		.dout(new_net_4200)
	);

	bfr new_net_4201_bfr_after (
		.din(new_net_4200),
		.dout(new_net_4201)
	);

	bfr new_net_4202_bfr_after (
		.din(new_net_4201),
		.dout(new_net_4202)
	);

	bfr new_net_4203_bfr_after (
		.din(new_net_4202),
		.dout(new_net_4203)
	);

	bfr new_net_4204_bfr_after (
		.din(new_net_4203),
		.dout(new_net_4204)
	);

	bfr new_net_4205_bfr_after (
		.din(new_net_4204),
		.dout(new_net_4205)
	);

	bfr new_net_4206_bfr_after (
		.din(new_net_4205),
		.dout(new_net_4206)
	);

	spl3L new_net_24_v_fanout (
		.a(new_net_4206),
		.b(G5196),
		.c(G5202),
		.d(G5201)
	);

	spl4L new_net_1872_v_fanout (
		.a(new_net_1872),
		.b(new_net_1665),
		.c(new_net_1869),
		.d(new_net_1660),
		.e(new_net_1870)
	);

	spl3L new_net_1891_v_fanout (
		.a(new_net_1891),
		.b(new_net_1609),
		.c(new_net_1610),
		.d(new_net_1611)
	);

	bfr new_net_4207_bfr_before (
		.din(new_net_4207),
		.dout(new_net_1396)
	);

	spl4L new_net_1907_v_fanout (
		.a(new_net_1907),
		.b(new_net_4207),
		.c(new_net_1394),
		.d(new_net_1395),
		.e(new_net_1393)
	);

	bfr new_net_4208_bfr_before (
		.din(new_net_4208),
		.dout(new_net_342)
	);

	spl3L new_net_1768_v_fanout (
		.a(new_net_1768),
		.b(new_net_337),
		.c(new_net_341),
		.d(new_net_4208)
	);

	spl4L new_net_1880_v_fanout (
		.a(new_net_1880),
		.b(new_net_952),
		.c(new_net_954),
		.d(new_net_953),
		.e(new_net_955)
	);

	spl2 new_net_1871_v_fanout (
		.a(new_net_1871),
		.b(new_net_1657),
		.c(new_net_1659)
	);

	bfr new_net_4209_bfr_before (
		.din(new_net_4209),
		.dout(new_net_750)
	);

	bfr new_net_4210_bfr_before (
		.din(new_net_4210),
		.dout(new_net_758)
	);

	spl4L new_net_1839_v_fanout (
		.a(new_net_1839),
		.b(new_net_4209),
		.c(new_net_4210),
		.d(new_net_759),
		.e(new_net_1836)
	);

	spl4L new_net_1888_v_fanout (
		.a(new_net_1888),
		.b(new_net_1313),
		.c(new_net_1314),
		.d(new_net_1315),
		.e(new_net_1312)
	);

	spl3L new_net_1903_v_fanout (
		.a(new_net_1903),
		.b(new_net_173),
		.c(new_net_177),
		.d(new_net_174)
	);

	spl3L new_net_1725_v_fanout (
		.a(new_net_1725),
		.b(new_net_1115),
		.c(new_net_1116),
		.d(new_net_1117)
	);

	bfr new_net_4211_bfr_before (
		.din(new_net_4211),
		.dout(new_net_986)
	);

	spl2 new_net_1773_v_fanout (
		.a(new_net_1773),
		.b(new_net_982),
		.c(new_net_4211)
	);

	bfr new_net_4212_bfr_before (
		.din(new_net_4212),
		.dout(new_net_1015)
	);

	bfr new_net_4213_bfr_before (
		.din(new_net_4213),
		.dout(new_net_1011)
	);

	spl4L new_net_1805_v_fanout (
		.a(new_net_1805),
		.b(new_net_1012),
		.c(new_net_4213),
		.d(new_net_1804),
		.e(new_net_4212)
	);

	bfr new_net_4214_bfr_before (
		.din(new_net_4214),
		.dout(new_net_1688)
	);

	bfr new_net_4215_bfr_before (
		.din(new_net_4215),
		.dout(new_net_1689)
	);

	spl4L new_net_1722_v_fanout (
		.a(new_net_1722),
		.b(new_net_4214),
		.c(new_net_4215),
		.d(new_net_1692),
		.e(new_net_1698)
	);

	spl4L new_net_1877_v_fanout (
		.a(new_net_1877),
		.b(new_net_1374),
		.c(new_net_1874),
		.d(new_net_1379),
		.e(new_net_1371)
	);

	spl2 new_net_1848_v_fanout (
		.a(new_net_1848),
		.b(new_net_1170),
		.c(new_net_1178)
	);

	bfr new_net_4216_bfr_before (
		.din(new_net_4216),
		.dout(new_net_1552)
	);

	spl4L new_net_1829_v_fanout (
		.a(new_net_1829),
		.b(new_net_1557),
		.c(new_net_1563),
		.d(new_net_4216),
		.e(new_net_1546)
	);

	spl4L new_net_1889_v_fanout (
		.a(new_net_1889),
		.b(new_net_1305),
		.c(new_net_1308),
		.d(new_net_1307),
		.e(new_net_1304)
	);

	spl3L new_net_1758_v_fanout (
		.a(new_net_1758),
		.b(new_net_839),
		.c(new_net_840),
		.d(new_net_841)
	);

	spl4L new_net_1759_v_fanout (
		.a(new_net_1759),
		.b(new_net_837),
		.c(new_net_838),
		.d(new_net_836),
		.e(new_net_835)
	);

	spl4L new_net_1764_v_fanout (
		.a(new_net_1764),
		.b(new_net_1472),
		.c(new_net_1468),
		.d(new_net_1469),
		.e(new_net_1466)
	);

	spl4L new_net_1827_v_fanout (
		.a(new_net_1827),
		.b(new_net_1553),
		.c(new_net_1826),
		.d(new_net_1551),
		.e(new_net_1560)
	);

	bfr new_net_4217_bfr_before (
		.din(new_net_4217),
		.dout(new_net_1139)
	);

	bfr new_net_4218_bfr_before (
		.din(new_net_4218),
		.dout(new_net_1144)
	);

	bfr new_net_4219_bfr_before (
		.din(new_net_4219),
		.dout(new_net_1142)
	);

	spl4L new_net_1748_v_fanout (
		.a(new_net_1748),
		.b(new_net_4218),
		.c(new_net_4219),
		.d(new_net_1143),
		.e(new_net_4217)
	);

	bfr new_net_4220_bfr_before (
		.din(new_net_4220),
		.dout(new_net_1001)
	);

	spl4L new_net_1806_v_fanout (
		.a(new_net_1806),
		.b(new_net_1005),
		.c(new_net_1002),
		.d(new_net_4220),
		.e(new_net_1803)
	);

	bfr new_net_4221_bfr_before (
		.din(new_net_4221),
		.dout(new_net_1176)
	);

	spl3L new_net_1849_v_fanout (
		.a(new_net_1849),
		.b(new_net_1846),
		.c(new_net_1847),
		.d(new_net_4221)
	);

	bfr new_net_4222_bfr_before (
		.din(new_net_4222),
		.dout(new_net_1052)
	);

	spl4L new_net_1845_v_fanout (
		.a(new_net_1845),
		.b(new_net_1039),
		.c(new_net_1841),
		.d(new_net_4222),
		.e(new_net_1843)
	);

	spl4L new_net_1747_v_fanout (
		.a(new_net_1747),
		.b(new_net_1141),
		.c(new_net_1140),
		.d(new_net_1138),
		.e(new_net_1137)
	);

	bfr new_net_4223_bfr_before (
		.din(new_net_4223),
		.dout(new_net_980)
	);

	bfr new_net_4224_bfr_before (
		.din(new_net_4224),
		.dout(new_net_989)
	);

	spl4L new_net_1776_v_fanout (
		.a(new_net_1776),
		.b(new_net_4223),
		.c(new_net_979),
		.d(new_net_4224),
		.e(new_net_987)
	);

	spl4L new_net_1890_v_fanout (
		.a(new_net_1890),
		.b(new_net_1310),
		.c(new_net_1311),
		.d(new_net_1309),
		.e(new_net_1306)
	);

	bfr new_net_4225_bfr_before (
		.din(new_net_4225),
		.dout(new_net_873)
	);

	bfr new_net_4226_bfr_before (
		.din(new_net_4226),
		.dout(new_net_880)
	);

	spl3L new_net_1815_v_fanout (
		.a(new_net_1815),
		.b(new_net_4225),
		.c(new_net_1814),
		.d(new_net_4226)
	);

	bfr new_net_4227_bfr_before (
		.din(new_net_4227),
		.dout(new_net_1014)
	);

	bfr new_net_4228_bfr_before (
		.din(new_net_4228),
		.dout(new_net_1009)
	);

	spl4L new_net_1807_v_fanout (
		.a(new_net_1807),
		.b(new_net_4227),
		.c(new_net_1016),
		.d(new_net_4228),
		.e(new_net_1007)
	);

	spl4L new_net_1853_v_fanout (
		.a(new_net_1853),
		.b(new_net_1673),
		.c(new_net_1666),
		.d(new_net_1850),
		.e(new_net_1851)
	);

	bfr new_net_4229_bfr_before (
		.din(new_net_4229),
		.dout(new_net_1250)
	);

	bfr new_net_4230_bfr_before (
		.din(new_net_4230),
		.dout(new_net_1247)
	);

	bfr new_net_4231_bfr_before (
		.din(new_net_4231),
		.dout(new_net_1244)
	);

	spl4L new_net_1781_v_fanout (
		.a(new_net_1781),
		.b(new_net_4229),
		.c(new_net_4230),
		.d(new_net_4231),
		.e(new_net_1248)
	);

	bfr new_net_4232_bfr_before (
		.din(new_net_4232),
		.dout(new_net_1558)
	);

	spl4L new_net_1830_v_fanout (
		.a(new_net_1830),
		.b(new_net_4232),
		.c(new_net_1547),
		.d(new_net_1545),
		.e(new_net_1825)
	);

	spl4L new_net_1767_v_fanout (
		.a(new_net_1767),
		.b(new_net_338),
		.c(new_net_339),
		.d(new_net_340),
		.e(new_net_335)
	);

	spl2 new_net_1754_v_fanout (
		.a(new_net_1754),
		.b(new_net_1753),
		.c(new_net_1751)
	);

	bfr new_net_4233_bfr_before (
		.din(new_net_4233),
		.dout(new_net_1694)
	);

	bfr new_net_4234_bfr_before (
		.din(new_net_4234),
		.dout(new_net_1690)
	);

	spl4L new_net_1723_v_fanout (
		.a(new_net_1723),
		.b(new_net_4233),
		.c(new_net_1693),
		.d(new_net_4234),
		.e(new_net_1691)
	);

	spl2 new_net_1879_v_fanout (
		.a(new_net_1879),
		.b(new_net_960),
		.c(new_net_961)
	);

	bfr new_net_4235_bfr_before (
		.din(new_net_4235),
		.dout(new_net_1066)
	);

	bfr new_net_4236_bfr_before (
		.din(new_net_4236),
		.dout(new_net_1071)
	);

	spl4L new_net_1811_v_fanout (
		.a(new_net_1811),
		.b(new_net_4235),
		.c(new_net_1809),
		.d(new_net_4236),
		.e(new_net_1808)
	);

	spl2 new_net_1886_v_fanout (
		.a(new_net_1886),
		.b(new_net_461),
		.c(new_net_1884)
	);

	bfr new_net_4237_bfr_before (
		.din(new_net_4237),
		.dout(new_net_875)
	);

	bfr new_net_4238_bfr_before (
		.din(new_net_4238),
		.dout(new_net_871)
	);

	bfr new_net_4239_bfr_before (
		.din(new_net_4239),
		.dout(new_net_877)
	);

	spl4L new_net_1816_v_fanout (
		.a(new_net_1816),
		.b(new_net_4237),
		.c(new_net_4238),
		.d(new_net_4239),
		.e(new_net_1813)
	);

	spl4L new_net_1881_v_fanout (
		.a(new_net_1881),
		.b(new_net_951),
		.c(new_net_957),
		.d(new_net_959),
		.e(new_net_956)
	);

	bfr new_net_4240_bfr_before (
		.din(new_net_4240),
		.dout(new_net_1042)
	);

	spl4L new_net_1844_v_fanout (
		.a(new_net_1844),
		.b(new_net_1044),
		.c(new_net_1842),
		.d(new_net_1047),
		.e(new_net_4240)
	);

	spl2 new_net_1834_v_fanout (
		.a(new_net_1834),
		.b(new_net_1634),
		.c(new_net_1638)
	);

	bfr new_net_4241_bfr_before (
		.din(new_net_4241),
		.dout(new_net_1602)
	);

	spl4L new_net_1892_v_fanout (
		.a(new_net_1892),
		.b(new_net_4241),
		.c(new_net_1606),
		.d(new_net_1604),
		.e(new_net_1612)
	);

	spl4L new_net_1828_v_fanout (
		.a(new_net_1828),
		.b(new_net_1559),
		.c(new_net_1550),
		.d(new_net_1544),
		.e(new_net_1554)
	);

	bfr new_net_4242_bfr_before (
		.din(new_net_4242),
		.dout(new_net_344)
	);

	spl2 new_net_1766_v_fanout (
		.a(new_net_1766),
		.b(new_net_4242),
		.c(new_net_1765)
	);

	bfr new_net_4243_bfr_before (
		.din(new_net_4243),
		.dout(new_net_753)
	);

	bfr new_net_4244_bfr_before (
		.din(new_net_4244),
		.dout(new_net_756)
	);

	spl4L new_net_1838_v_fanout (
		.a(new_net_1838),
		.b(new_net_4243),
		.c(new_net_4244),
		.d(new_net_1837),
		.e(new_net_754)
	);

	bfr new_net_4245_bfr_before (
		.din(new_net_4245),
		.dout(new_net_1118)
	);

	bfr new_net_4246_bfr_before (
		.din(new_net_4246),
		.dout(new_net_1108)
	);

	bfr new_net_4247_bfr_before (
		.din(new_net_4247),
		.dout(new_net_1111)
	);

	spl4L new_net_1726_v_fanout (
		.a(new_net_1726),
		.b(new_net_4246),
		.c(new_net_4247),
		.d(new_net_1109),
		.e(new_net_4245)
	);

	bfr new_net_4248_bfr_before (
		.din(new_net_4248),
		.dout(new_net_1868)
	);

	bfr new_net_4249_bfr_before (
		.din(new_net_4249),
		.dout(new_net_4248)
	);

	spl3L new_net_1867_v_fanout (
		.a(new_net_1867),
		.b(new_net_1266),
		.c(new_net_4249),
		.d(new_net_1267)
	);

	bfr new_net_4250_bfr_before (
		.din(new_net_4250),
		.dout(new_net_1032)
	);

	spl3L new_net_1833_v_fanout (
		.a(new_net_1833),
		.b(new_net_1033),
		.c(new_net_1031),
		.d(new_net_4250)
	);

	bfr new_net_4251_bfr_before (
		.din(new_net_4251),
		.dout(new_net_991)
	);

	bfr new_net_4252_bfr_before (
		.din(new_net_4252),
		.dout(new_net_984)
	);

	spl4L new_net_1774_v_fanout (
		.a(new_net_1774),
		.b(new_net_4251),
		.c(new_net_1771),
		.d(new_net_4252),
		.e(new_net_981)
	);

	spl3L new_net_1746_v_fanout (
		.a(new_net_1746),
		.b(new_net_1145),
		.c(new_net_1146),
		.d(new_net_1147)
	);

	bfr new_net_4253_bfr_before (
		.din(new_net_4253),
		.dout(new_net_1243)
	);

	spl2 new_net_1780_v_fanout (
		.a(new_net_1780),
		.b(new_net_1779),
		.c(new_net_4253)
	);

	bfr new_net_4254_bfr_before (
		.din(new_net_4254),
		.dout(new_net_1414)
	);

	bfr new_net_4255_bfr_before (
		.din(new_net_4255),
		.dout(new_net_1412)
	);

	bfr new_net_4256_bfr_before (
		.din(new_net_4256),
		.dout(new_net_1413)
	);

	spl4L new_net_1757_v_fanout (
		.a(new_net_1757),
		.b(new_net_4254),
		.c(new_net_4255),
		.d(new_net_4256),
		.e(new_net_1418)
	);

	bfr new_net_4257_bfr_before (
		.din(new_net_4257),
		.dout(new_net_1674)
	);

	spl2 new_net_1852_v_fanout (
		.a(new_net_1852),
		.b(new_net_1668),
		.c(new_net_4257)
	);

	bfr new_net_4258_bfr_before (
		.din(new_net_4258),
		.dout(G5213)
	);

	bfr new_net_4259_bfr_before (
		.din(new_net_4259),
		.dout(new_net_4258)
	);

	bfr new_net_4260_bfr_before (
		.din(new_net_4260),
		.dout(new_net_4259)
	);

	bfr new_net_4261_bfr_before (
		.din(new_net_4261),
		.dout(new_net_4260)
	);

	bfr new_net_4262_bfr_before (
		.din(new_net_4262),
		.dout(new_net_4261)
	);

	bfr new_net_4263_bfr_before (
		.din(new_net_4263),
		.dout(new_net_4262)
	);

	bfr new_net_4264_bfr_before (
		.din(new_net_4264),
		.dout(new_net_4263)
	);

	bfr new_net_4265_bfr_before (
		.din(new_net_4265),
		.dout(new_net_4264)
	);

	bfr new_net_4266_bfr_before (
		.din(new_net_4266),
		.dout(new_net_4265)
	);

	bfr new_net_4267_bfr_before (
		.din(new_net_4267),
		.dout(new_net_4266)
	);

	bfr new_net_4268_bfr_before (
		.din(new_net_4268),
		.dout(new_net_4267)
	);

	bfr new_net_4269_bfr_before (
		.din(new_net_4269),
		.dout(new_net_4268)
	);

	bfr new_net_4270_bfr_before (
		.din(new_net_4270),
		.dout(new_net_4269)
	);

	bfr new_net_4271_bfr_before (
		.din(new_net_4271),
		.dout(new_net_4270)
	);

	bfr new_net_4272_bfr_before (
		.din(new_net_4272),
		.dout(new_net_4271)
	);

	bfr new_net_4273_bfr_before (
		.din(new_net_4273),
		.dout(new_net_4272)
	);

	bfr new_net_4274_bfr_before (
		.din(new_net_4274),
		.dout(new_net_4273)
	);

	bfr new_net_4275_bfr_before (
		.din(new_net_4275),
		.dout(new_net_4274)
	);

	bfr new_net_4276_bfr_before (
		.din(new_net_4276),
		.dout(new_net_4275)
	);

	bfr new_net_4277_bfr_before (
		.din(new_net_4277),
		.dout(new_net_4276)
	);

	bfr new_net_4278_bfr_before (
		.din(new_net_4278),
		.dout(new_net_4277)
	);

	bfr new_net_4279_bfr_before (
		.din(new_net_4279),
		.dout(new_net_4278)
	);

	bfr new_net_4280_bfr_before (
		.din(new_net_4280),
		.dout(new_net_4279)
	);

	bfr new_net_4281_bfr_before (
		.din(new_net_4281),
		.dout(new_net_4280)
	);

	bfr new_net_4282_bfr_before (
		.din(new_net_4282),
		.dout(new_net_4281)
	);

	bfr new_net_4283_bfr_before (
		.din(new_net_4283),
		.dout(new_net_4282)
	);

	bfr new_net_4284_bfr_before (
		.din(new_net_4284),
		.dout(new_net_4283)
	);

	bfr new_net_4285_bfr_before (
		.din(new_net_4285),
		.dout(new_net_4284)
	);

	bfr new_net_4286_bfr_before (
		.din(new_net_4286),
		.dout(new_net_4285)
	);

	bfr new_net_4287_bfr_before (
		.din(new_net_4287),
		.dout(new_net_4286)
	);

	bfr new_net_4288_bfr_before (
		.din(new_net_4288),
		.dout(new_net_4287)
	);

	bfr new_net_4289_bfr_before (
		.din(new_net_4289),
		.dout(new_net_4288)
	);

	bfr new_net_4290_bfr_before (
		.din(new_net_4290),
		.dout(new_net_4289)
	);

	bfr new_net_4291_bfr_before (
		.din(new_net_4291),
		.dout(new_net_4290)
	);

	bfr new_net_4292_bfr_before (
		.din(new_net_4292),
		.dout(new_net_4291)
	);

	bfr new_net_4293_bfr_before (
		.din(new_net_4293),
		.dout(new_net_4292)
	);

	bfr new_net_4294_bfr_before (
		.din(new_net_4294),
		.dout(new_net_4293)
	);

	bfr new_net_4295_bfr_before (
		.din(new_net_4295),
		.dout(new_net_4294)
	);

	bfr new_net_4296_bfr_before (
		.din(new_net_4296),
		.dout(new_net_4295)
	);

	bfr new_net_4297_bfr_before (
		.din(new_net_4297),
		.dout(new_net_4296)
	);

	spl2 new_net_13_v_fanout (
		.a(new_net_13),
		.b(new_net_4297),
		.c(new_net_748)
	);

	spl3L new_net_1721_v_fanout (
		.a(new_net_1721),
		.b(new_net_1695),
		.c(new_net_1696),
		.d(new_net_1697)
	);

	spl3L new_net_1906_v_fanout (
		.a(new_net_1906),
		.b(new_net_1397),
		.c(new_net_1398),
		.d(new_net_1399)
	);

	bfr new_net_4298_bfr_before (
		.din(new_net_4298),
		.dout(new_net_1416)
	);

	bfr new_net_4299_bfr_before (
		.din(new_net_4299),
		.dout(new_net_1417)
	);

	spl3L new_net_1756_v_fanout (
		.a(new_net_1756),
		.b(new_net_4298),
		.c(new_net_1415),
		.d(new_net_4299)
	);

	bfr new_net_4300_bfr_before (
		.din(new_net_4300),
		.dout(new_net_1471)
	);

	bfr new_net_4301_bfr_before (
		.din(new_net_4301),
		.dout(new_net_1473)
	);

	bfr new_net_4302_bfr_before (
		.din(new_net_4302),
		.dout(new_net_1474)
	);

	spl4L new_net_1763_v_fanout (
		.a(new_net_1763),
		.b(new_net_4301),
		.c(new_net_4302),
		.d(new_net_1760),
		.e(new_net_4300)
	);

	bfr new_net_4303_bfr_before (
		.din(new_net_4303),
		.dout(new_net_175)
	);

	spl2 new_net_1902_v_fanout (
		.a(new_net_1902),
		.b(new_net_4303),
		.c(new_net_176)
	);

	bfr new_net_4304_bfr_before (
		.din(new_net_4304),
		.dout(new_net_1633)
	);

	bfr new_net_4305_bfr_before (
		.din(new_net_4305),
		.dout(new_net_1637)
	);

	bfr new_net_4306_bfr_before (
		.din(new_net_4306),
		.dout(new_net_1635)
	);

	spl4L new_net_1835_v_fanout (
		.a(new_net_1835),
		.b(new_net_4305),
		.c(new_net_4306),
		.d(new_net_1636),
		.e(new_net_4304)
	);

	spl4L new_net_1727_v_fanout (
		.a(new_net_1727),
		.b(new_net_1114),
		.c(new_net_1113),
		.d(new_net_1110),
		.e(new_net_1112)
	);

	bfr new_net_4307_bfr_before (
		.din(new_net_4307),
		.dout(new_net_1289)
	);

	bfr new_net_4308_bfr_before (
		.din(new_net_4308),
		.dout(new_net_4307)
	);

	bfr new_net_4309_bfr_before (
		.din(new_net_4309),
		.dout(new_net_4308)
	);

	spl2 G149_v_fanout (
		.a(G149),
		.b(new_net_1288),
		.c(new_net_4309)
	);

	bfr new_net_4310_bfr_after (
		.din(G69),
		.dout(new_net_4310)
	);

	bfr new_net_4311_bfr_after (
		.din(new_net_4310),
		.dout(new_net_4311)
	);

	bfr new_net_4312_bfr_after (
		.din(new_net_4311),
		.dout(new_net_4312)
	);

	spl2 G69_v_fanout (
		.a(new_net_4312),
		.b(new_net_1322),
		.c(new_net_1323)
	);

	bfr new_net_4313_bfr_before (
		.din(new_net_4313),
		.dout(new_net_1721)
	);

	spl3L G167_v_fanout (
		.a(G167),
		.b(new_net_1722),
		.c(new_net_4313),
		.d(new_net_1723)
	);

	bfr new_net_4314_bfr_before (
		.din(new_net_4314),
		.dout(new_net_1724)
	);

	bfr new_net_4315_bfr_before (
		.din(new_net_4315),
		.dout(new_net_4314)
	);

	bfr new_net_4316_bfr_before (
		.din(new_net_4316),
		.dout(new_net_4315)
	);

	bfr new_net_4317_bfr_before (
		.din(new_net_4317),
		.dout(new_net_4316)
	);

	spl2 G141_v_fanout (
		.a(G141),
		.b(new_net_4317),
		.c(new_net_1079)
	);

	bfr new_net_4318_bfr_before (
		.din(new_net_4318),
		.dout(new_net_1727)
	);

	bfr new_net_4319_bfr_before (
		.din(new_net_4319),
		.dout(new_net_1725)
	);

	spl3L G105_v_fanout (
		.a(G105),
		.b(new_net_4318),
		.c(new_net_4319),
		.d(new_net_1726)
	);

	bfr new_net_4320_bfr_after (
		.din(G27),
		.dout(new_net_4320)
	);

	bfr new_net_4321_bfr_after (
		.din(new_net_4320),
		.dout(new_net_4321)
	);

	bfr new_net_4322_bfr_after (
		.din(new_net_4321),
		.dout(new_net_4322)
	);

	spl2 G27_v_fanout (
		.a(new_net_4322),
		.b(new_net_790),
		.c(new_net_791)
	);

	bfr new_net_4323_bfr_after (
		.din(G21),
		.dout(new_net_4323)
	);

	bfr new_net_4324_bfr_after (
		.din(new_net_4323),
		.dout(new_net_4324)
	);

	bfr new_net_4325_bfr_after (
		.din(new_net_4324),
		.dout(new_net_4325)
	);

	bfr new_net_4326_bfr_after (
		.din(new_net_4325),
		.dout(new_net_4326)
	);

	bfr new_net_4327_bfr_after (
		.din(new_net_4326),
		.dout(new_net_4327)
	);

	bfr new_net_4328_bfr_after (
		.din(new_net_4327),
		.dout(new_net_4328)
	);

	spl2 G21_v_fanout (
		.a(new_net_4328),
		.b(new_net_331),
		.c(new_net_332)
	);

	bfr new_net_4329_bfr_after (
		.din(G5),
		.dout(new_net_4329)
	);

	bfr new_net_4330_bfr_after (
		.din(new_net_4329),
		.dout(new_net_4330)
	);

	bfr new_net_4331_bfr_after (
		.din(new_net_4330),
		.dout(new_net_4331)
	);

	spl2 G5_v_fanout (
		.a(new_net_4331),
		.b(new_net_882),
		.c(new_net_883)
	);

	bfr new_net_4332_bfr_after (
		.din(G4),
		.dout(new_net_4332)
	);

	bfr new_net_4333_bfr_after (
		.din(new_net_4332),
		.dout(new_net_4333)
	);

	bfr new_net_4334_bfr_after (
		.din(new_net_4333),
		.dout(new_net_4334)
	);

	spl2 G4_v_fanout (
		.a(new_net_4334),
		.b(new_net_525),
		.c(new_net_526)
	);

	bfr new_net_4335_bfr_before (
		.din(new_net_4335),
		.dout(new_net_996)
	);

	bfr new_net_4336_bfr_before (
		.din(new_net_4336),
		.dout(new_net_4335)
	);

	bfr new_net_4337_bfr_before (
		.din(new_net_4337),
		.dout(new_net_4336)
	);

	bfr new_net_4338_bfr_before (
		.din(new_net_4338),
		.dout(new_net_4337)
	);

	bfr new_net_4339_bfr_before (
		.din(new_net_4339),
		.dout(new_net_4338)
	);

	bfr new_net_4340_bfr_before (
		.din(new_net_4340),
		.dout(new_net_4339)
	);

	spl2 G139_v_fanout (
		.a(G139),
		.b(new_net_995),
		.c(new_net_4340)
	);

	bfr new_net_4341_bfr_before (
		.din(new_net_4341),
		.dout(new_net_1745)
	);

	bfr new_net_4342_bfr_before (
		.din(new_net_4342),
		.dout(new_net_4341)
	);

	bfr new_net_4343_bfr_before (
		.din(new_net_4343),
		.dout(new_net_4342)
	);

	bfr new_net_4344_bfr_before (
		.din(new_net_4344),
		.dout(new_net_1728)
	);

	bfr new_net_4345_bfr_before (
		.din(new_net_4345),
		.dout(new_net_4344)
	);

	bfr new_net_4346_bfr_before (
		.din(new_net_4346),
		.dout(new_net_4345)
	);

	spl4L G176_v_fanout (
		.a(G176),
		.b(new_net_1232),
		.c(new_net_4343),
		.d(new_net_4346),
		.e(new_net_1230)
	);

	bfr new_net_4347_bfr_after (
		.din(G111),
		.dout(new_net_4347)
	);

	spl3L G111_v_fanout (
		.a(new_net_4347),
		.b(new_net_1296),
		.c(new_net_1298),
		.d(new_net_1297)
	);

	bfr new_net_4348_bfr_before (
		.din(new_net_4348),
		.dout(new_net_1747)
	);

	bfr new_net_4349_bfr_before (
		.din(new_net_4349),
		.dout(new_net_1746)
	);

	spl3L G96_v_fanout (
		.a(G96),
		.b(new_net_1748),
		.c(new_net_4348),
		.d(new_net_4349)
	);

	bfr new_net_4350_bfr_after (
		.din(G71),
		.dout(new_net_4350)
	);

	bfr new_net_4351_bfr_after (
		.din(new_net_4350),
		.dout(new_net_4351)
	);

	bfr new_net_4352_bfr_after (
		.din(new_net_4351),
		.dout(new_net_4352)
	);

	spl2 G71_v_fanout (
		.a(new_net_4352),
		.b(new_net_1358),
		.c(new_net_1359)
	);

	spl2 G155_v_fanout (
		.a(G155),
		.b(new_net_1400),
		.c(new_net_1401)
	);

	spl2 G123_v_fanout (
		.a(G123),
		.b(new_net_1754),
		.c(new_net_1755)
	);

	spl2 G119_v_fanout (
		.a(G119),
		.b(new_net_1757),
		.c(new_net_1756)
	);

	bfr new_net_4353_bfr_before (
		.din(new_net_4353),
		.dout(new_net_1625)
	);

	bfr new_net_4354_bfr_before (
		.din(new_net_4354),
		.dout(new_net_4353)
	);

	spl2 G127_v_fanout (
		.a(G127),
		.b(new_net_1624),
		.c(new_net_4354)
	);

	bfr new_net_4355_bfr_after (
		.din(G82),
		.dout(new_net_4355)
	);

	bfr new_net_4356_bfr_after (
		.din(new_net_4355),
		.dout(new_net_4356)
	);

	bfr new_net_4357_bfr_after (
		.din(new_net_4356),
		.dout(new_net_4357)
	);

	spl2 G82_v_fanout (
		.a(new_net_4357),
		.b(new_net_413),
		.c(new_net_414)
	);

	bfr new_net_4358_bfr_after (
		.din(G88),
		.dout(new_net_4358)
	);

	spl2 G88_v_fanout (
		.a(new_net_4358),
		.b(new_net_1758),
		.c(new_net_1759)
	);

	bfr new_net_4359_bfr_before (
		.din(new_net_4359),
		.dout(new_net_1764)
	);

	spl2 G121_v_fanout (
		.a(G121),
		.b(new_net_1763),
		.c(new_net_4359)
	);

	bfr new_net_4360_bfr_before (
		.din(new_net_4360),
		.dout(new_net_1767)
	);

	spl3L G168_v_fanout (
		.a(G168),
		.b(new_net_1768),
		.c(new_net_1766),
		.d(new_net_4360)
	);

	bfr new_net_4361_bfr_after (
		.din(G72),
		.dout(new_net_4361)
	);

	bfr new_net_4362_bfr_after (
		.din(new_net_4361),
		.dout(new_net_4362)
	);

	bfr new_net_4363_bfr_after (
		.din(new_net_4362),
		.dout(new_net_4363)
	);

	spl2 G72_v_fanout (
		.a(new_net_4363),
		.b(new_net_1385),
		.c(new_net_1386)
	);

	bfr new_net_4364_bfr_after (
		.din(G87),
		.dout(new_net_4364)
	);

	bfr new_net_4365_bfr_after (
		.din(new_net_4364),
		.dout(new_net_4365)
	);

	bfr new_net_4366_bfr_after (
		.din(new_net_4365),
		.dout(new_net_4366)
	);

	spl2 G87_v_fanout (
		.a(new_net_4366),
		.b(new_net_816),
		.c(new_net_817)
	);

	spl2 G165_v_fanout (
		.a(G165),
		.b(new_net_1626),
		.c(new_net_1627)
	);

	bfr new_net_4367_bfr_after (
		.din(G75),
		.dout(new_net_4367)
	);

	bfr new_net_4368_bfr_after (
		.din(new_net_4367),
		.dout(new_net_4368)
	);

	bfr new_net_4369_bfr_after (
		.din(new_net_4368),
		.dout(new_net_4369)
	);

	spl2 G75_v_fanout (
		.a(new_net_4369),
		.b(new_net_1421),
		.c(new_net_1422)
	);

	bfr new_net_4370_bfr_after (
		.din(G18),
		.dout(new_net_4370)
	);

	bfr new_net_4371_bfr_after (
		.din(new_net_4370),
		.dout(new_net_4371)
	);

	bfr new_net_4372_bfr_after (
		.din(new_net_4371),
		.dout(new_net_4372)
	);

	spl2 G18_v_fanout (
		.a(new_net_4372),
		.b(new_net_1489),
		.c(new_net_1490)
	);

	bfr new_net_4373_bfr_after (
		.din(G162),
		.dout(new_net_4373)
	);

	bfr new_net_4374_bfr_after (
		.din(new_net_4373),
		.dout(new_net_4374)
	);

	bfr new_net_4375_bfr_after (
		.din(new_net_4374),
		.dout(new_net_4375)
	);

	bfr new_net_4376_bfr_after (
		.din(new_net_4375),
		.dout(new_net_4376)
	);

	bfr new_net_4377_bfr_after (
		.din(new_net_4376),
		.dout(new_net_4377)
	);

	bfr new_net_4378_bfr_after (
		.din(new_net_4377),
		.dout(new_net_4378)
	);

	bfr new_net_4379_bfr_before (
		.din(new_net_4379),
		.dout(new_net_1191)
	);

	bfr new_net_4380_bfr_before (
		.din(new_net_4380),
		.dout(new_net_4379)
	);

	spl2 G162_v_fanout (
		.a(new_net_4378),
		.b(new_net_1190),
		.c(new_net_4380)
	);

	bfr new_net_4381_bfr_before (
		.din(new_net_4381),
		.dout(new_net_1770)
	);

	bfr new_net_4382_bfr_before (
		.din(new_net_4382),
		.dout(new_net_4381)
	);

	bfr new_net_4383_bfr_before (
		.din(new_net_4383),
		.dout(new_net_4382)
	);

	bfr new_net_4384_bfr_before (
		.din(new_net_4384),
		.dout(new_net_4383)
	);

	bfr new_net_4385_bfr_before (
		.din(new_net_4385),
		.dout(new_net_1769)
	);

	bfr new_net_4386_bfr_before (
		.din(new_net_4386),
		.dout(new_net_4385)
	);

	bfr new_net_4387_bfr_before (
		.din(new_net_4387),
		.dout(new_net_4386)
	);

	bfr new_net_4388_bfr_before (
		.din(new_net_4388),
		.dout(new_net_4387)
	);

	spl4L G66_v_fanout (
		.a(G66),
		.b(new_net_1277),
		.c(new_net_1275),
		.d(new_net_4388),
		.e(new_net_4384)
	);

	bfr new_net_4389_bfr_before (
		.din(new_net_4389),
		.dout(new_net_1261)
	);

	bfr new_net_4390_bfr_before (
		.din(new_net_4390),
		.dout(new_net_4389)
	);

	spl2 G125_v_fanout (
		.a(G125),
		.b(new_net_1260),
		.c(new_net_4390)
	);

	spl4L G100_v_fanout (
		.a(G100),
		.b(new_net_1773),
		.c(new_net_1774),
		.d(new_net_1776),
		.e(new_net_1775)
	);

	bfr new_net_4391_bfr_after (
		.din(G61),
		.dout(new_net_4391)
	);

	bfr new_net_4392_bfr_after (
		.din(new_net_4391),
		.dout(new_net_4392)
	);

	bfr new_net_4393_bfr_after (
		.din(new_net_4392),
		.dout(new_net_4393)
	);

	bfr new_net_4394_bfr_after (
		.din(new_net_4393),
		.dout(new_net_4394)
	);

	bfr new_net_4395_bfr_after (
		.din(new_net_4394),
		.dout(new_net_4395)
	);

	spl2 G61_v_fanout (
		.a(new_net_4395),
		.b(new_net_1101),
		.c(new_net_1102)
	);

	bfr new_net_4396_bfr_before (
		.din(new_net_4396),
		.dout(new_net_1777)
	);

	bfr new_net_4397_bfr_before (
		.din(new_net_4397),
		.dout(new_net_4396)
	);

	bfr new_net_4398_bfr_before (
		.din(new_net_4398),
		.dout(new_net_4397)
	);

	spl2 G147_v_fanout (
		.a(G147),
		.b(new_net_4398),
		.c(new_net_1255)
	);

	bfr new_net_4399_bfr_after (
		.din(G86),
		.dout(new_net_4399)
	);

	bfr new_net_4400_bfr_after (
		.din(new_net_4399),
		.dout(new_net_4400)
	);

	bfr new_net_4401_bfr_after (
		.din(new_net_4400),
		.dout(new_net_4401)
	);

	spl2 G86_v_fanout (
		.a(new_net_4401),
		.b(new_net_808),
		.c(new_net_809)
	);

	bfr new_net_4402_bfr_after (
		.din(G85),
		.dout(new_net_4402)
	);

	bfr new_net_4403_bfr_after (
		.din(new_net_4402),
		.dout(new_net_4403)
	);

	bfr new_net_4404_bfr_after (
		.din(new_net_4403),
		.dout(new_net_4404)
	);

	spl2 G85_v_fanout (
		.a(new_net_4404),
		.b(new_net_1705),
		.c(new_net_1706)
	);

	bfr new_net_4405_bfr_after (
		.din(G73),
		.dout(new_net_4405)
	);

	bfr new_net_4406_bfr_after (
		.din(new_net_4405),
		.dout(new_net_4406)
	);

	bfr new_net_4407_bfr_after (
		.din(new_net_4406),
		.dout(new_net_4407)
	);

	spl2 G73_v_fanout (
		.a(new_net_4407),
		.b(new_net_1391),
		.c(new_net_1392)
	);

	bfr new_net_4408_bfr_after (
		.din(G39),
		.dout(new_net_4408)
	);

	bfr new_net_4409_bfr_after (
		.din(new_net_4408),
		.dout(new_net_4409)
	);

	bfr new_net_4410_bfr_after (
		.din(new_net_4409),
		.dout(new_net_4410)
	);

	spl2 G39_v_fanout (
		.a(new_net_4410),
		.b(new_net_468),
		.c(new_net_469)
	);

	bfr new_net_4411_bfr_after (
		.din(G25),
		.dout(new_net_4411)
	);

	bfr new_net_4412_bfr_after (
		.din(new_net_4411),
		.dout(new_net_4412)
	);

	bfr new_net_4413_bfr_after (
		.din(new_net_4412),
		.dout(new_net_4413)
	);

	spl2 G25_v_fanout (
		.a(new_net_4413),
		.b(new_net_593),
		.c(new_net_594)
	);

	bfr new_net_4414_bfr_before (
		.din(new_net_4414),
		.dout(new_net_1419)
	);

	bfr new_net_4415_bfr_before (
		.din(new_net_4415),
		.dout(new_net_4414)
	);

	bfr new_net_4416_bfr_before (
		.din(new_net_4416),
		.dout(new_net_4415)
	);

	bfr new_net_4417_bfr_before (
		.din(new_net_4417),
		.dout(new_net_4416)
	);

	bfr new_net_4418_bfr_before (
		.din(new_net_4418),
		.dout(new_net_4417)
	);

	bfr new_net_4419_bfr_before (
		.din(new_net_4419),
		.dout(new_net_4418)
	);

	bfr new_net_4420_bfr_before (
		.din(new_net_4420),
		.dout(new_net_4419)
	);

	bfr new_net_4421_bfr_before (
		.din(new_net_4421),
		.dout(new_net_4420)
	);

	bfr new_net_4422_bfr_before (
		.din(new_net_4422),
		.dout(new_net_4421)
	);

	bfr new_net_4423_bfr_before (
		.din(new_net_4423),
		.dout(new_net_4422)
	);

	bfr new_net_4424_bfr_before (
		.din(new_net_4424),
		.dout(new_net_4423)
	);

	bfr new_net_4425_bfr_before (
		.din(new_net_4425),
		.dout(new_net_4424)
	);

	bfr new_net_4426_bfr_before (
		.din(new_net_4426),
		.dout(new_net_4425)
	);

	bfr new_net_4427_bfr_before (
		.din(new_net_4427),
		.dout(new_net_4426)
	);

	bfr new_net_4428_bfr_before (
		.din(new_net_4428),
		.dout(new_net_4427)
	);

	bfr new_net_4429_bfr_before (
		.din(new_net_4429),
		.dout(new_net_4428)
	);

	bfr new_net_4430_bfr_before (
		.din(new_net_4430),
		.dout(new_net_4429)
	);

	bfr new_net_4431_bfr_before (
		.din(new_net_4431),
		.dout(new_net_4430)
	);

	bfr new_net_4432_bfr_before (
		.din(new_net_4432),
		.dout(new_net_4431)
	);

	bfr new_net_4433_bfr_before (
		.din(new_net_4433),
		.dout(new_net_4432)
	);

	bfr new_net_4434_bfr_before (
		.din(new_net_4434),
		.dout(new_net_4433)
	);

	bfr new_net_4435_bfr_before (
		.din(new_net_4435),
		.dout(new_net_4434)
	);

	spl2 G157_v_fanout (
		.a(G157),
		.b(new_net_4435),
		.c(new_net_1420)
	);

	spl3L G109_v_fanout (
		.a(G109),
		.b(new_net_1780),
		.c(new_net_1781),
		.d(new_net_1782)
	);

	spl2 G156_v_fanout (
		.a(G156),
		.b(new_net_1404),
		.c(new_net_1405)
	);

	bfr new_net_4436_bfr_after (
		.din(G2),
		.dout(new_net_4436)
	);

	bfr new_net_4437_bfr_after (
		.din(new_net_4436),
		.dout(new_net_4437)
	);

	bfr new_net_4438_bfr_after (
		.din(new_net_4437),
		.dout(new_net_4438)
	);

	bfr new_net_4439_bfr_after (
		.din(new_net_4438),
		.dout(new_net_4439)
	);

	bfr new_net_4440_bfr_after (
		.din(new_net_4439),
		.dout(new_net_4440)
	);

	bfr new_net_4441_bfr_after (
		.din(new_net_4440),
		.dout(new_net_4441)
	);

	bfr new_net_4442_bfr_after (
		.din(new_net_4441),
		.dout(new_net_4442)
	);

	bfr new_net_4443_bfr_after (
		.din(new_net_4442),
		.dout(new_net_4443)
	);

	bfr new_net_4444_bfr_after (
		.din(new_net_4443),
		.dout(new_net_4444)
	);

	bfr new_net_4445_bfr_before (
		.din(new_net_4445),
		.dout(new_net_1783)
	);

	bfr new_net_4446_bfr_before (
		.din(new_net_4446),
		.dout(new_net_4445)
	);

	bfr new_net_4447_bfr_before (
		.din(new_net_4447),
		.dout(new_net_4446)
	);

	spl3L G2_v_fanout (
		.a(new_net_4444),
		.b(new_net_50),
		.c(new_net_53),
		.d(new_net_4447)
	);

	bfr new_net_4448_bfr_after (
		.din(G146),
		.dout(new_net_4448)
	);

	bfr new_net_4449_bfr_after (
		.din(new_net_4448),
		.dout(new_net_4449)
	);

	bfr new_net_4450_bfr_after (
		.din(new_net_4449),
		.dout(new_net_4450)
	);

	bfr new_net_4451_bfr_before (
		.din(new_net_4451),
		.dout(new_net_1195)
	);

	spl2 G146_v_fanout (
		.a(new_net_4450),
		.b(new_net_4451),
		.c(new_net_1785)
	);

	bfr new_net_4452_bfr_after (
		.din(G41),
		.dout(new_net_4452)
	);

	bfr new_net_4453_bfr_after (
		.din(new_net_4452),
		.dout(new_net_4453)
	);

	bfr new_net_4454_bfr_after (
		.din(new_net_4453),
		.dout(new_net_4454)
	);

	spl2 G41_v_fanout (
		.a(new_net_4454),
		.b(new_net_692),
		.c(new_net_693)
	);

	bfr new_net_4455_bfr_after (
		.din(G68),
		.dout(new_net_4455)
	);

	bfr new_net_4456_bfr_after (
		.din(new_net_4455),
		.dout(new_net_4456)
	);

	bfr new_net_4457_bfr_after (
		.din(new_net_4456),
		.dout(new_net_4457)
	);

	spl2 G68_v_fanout (
		.a(new_net_4457),
		.b(new_net_1302),
		.c(new_net_1303)
	);

	spl3L G159_v_fanout (
		.a(G159),
		.b(new_net_1453),
		.c(new_net_1455),
		.d(new_net_1454)
	);

	bfr new_net_4458_bfr_before (
		.din(new_net_4458),
		.dout(new_net_1787)
	);

	bfr new_net_4459_bfr_before (
		.din(new_net_4459),
		.dout(new_net_4458)
	);

	bfr new_net_4460_bfr_before (
		.din(new_net_4460),
		.dout(new_net_4459)
	);

	bfr new_net_4461_bfr_before (
		.din(new_net_4461),
		.dout(new_net_4460)
	);

	spl2 G135_v_fanout (
		.a(G135),
		.b(new_net_900),
		.c(new_net_4461)
	);

	bfr new_net_4462_bfr_before (
		.din(new_net_4462),
		.dout(new_net_1788)
	);

	bfr new_net_4463_bfr_before (
		.din(new_net_4463),
		.dout(new_net_4462)
	);

	bfr new_net_4464_bfr_before (
		.din(new_net_4464),
		.dout(new_net_4463)
	);

	bfr new_net_4465_bfr_before (
		.din(new_net_4465),
		.dout(new_net_4464)
	);

	bfr new_net_4466_bfr_before (
		.din(new_net_4466),
		.dout(new_net_4465)
	);

	bfr new_net_4467_bfr_before (
		.din(new_net_4467),
		.dout(new_net_4466)
	);

	bfr new_net_4468_bfr_before (
		.din(new_net_4468),
		.dout(new_net_4467)
	);

	bfr new_net_4469_bfr_before (
		.din(new_net_4469),
		.dout(new_net_4468)
	);

	bfr new_net_4470_bfr_before (
		.din(new_net_4470),
		.dout(new_net_4469)
	);

	bfr new_net_4471_bfr_before (
		.din(new_net_4471),
		.dout(new_net_4470)
	);

	bfr new_net_4472_bfr_before (
		.din(new_net_4472),
		.dout(new_net_4471)
	);

	bfr new_net_4473_bfr_before (
		.din(new_net_4473),
		.dout(new_net_4472)
	);

	bfr new_net_4474_bfr_before (
		.din(new_net_4474),
		.dout(new_net_4473)
	);

	bfr new_net_4475_bfr_before (
		.din(new_net_4475),
		.dout(new_net_4474)
	);

	bfr new_net_4476_bfr_before (
		.din(new_net_4476),
		.dout(new_net_4475)
	);

	bfr new_net_4477_bfr_before (
		.din(new_net_4477),
		.dout(new_net_4476)
	);

	bfr new_net_4478_bfr_before (
		.din(new_net_4478),
		.dout(new_net_4477)
	);

	bfr new_net_4479_bfr_before (
		.din(new_net_4479),
		.dout(new_net_4478)
	);

	bfr new_net_4480_bfr_before (
		.din(new_net_4480),
		.dout(new_net_4479)
	);

	bfr new_net_4481_bfr_before (
		.din(new_net_4481),
		.dout(new_net_4480)
	);

	bfr new_net_4482_bfr_before (
		.din(new_net_4482),
		.dout(new_net_4481)
	);

	bfr new_net_4483_bfr_before (
		.din(new_net_4483),
		.dout(new_net_4482)
	);

	bfr new_net_4484_bfr_before (
		.din(new_net_4484),
		.dout(new_net_4483)
	);

	bfr new_net_4485_bfr_before (
		.din(new_net_4485),
		.dout(new_net_4484)
	);

	bfr new_net_4486_bfr_before (
		.din(new_net_4486),
		.dout(new_net_4485)
	);

	bfr new_net_4487_bfr_before (
		.din(new_net_4487),
		.dout(new_net_4486)
	);

	bfr new_net_4488_bfr_before (
		.din(new_net_4488),
		.dout(new_net_4487)
	);

	bfr new_net_4489_bfr_before (
		.din(new_net_4489),
		.dout(new_net_4488)
	);

	bfr new_net_4490_bfr_before (
		.din(new_net_4490),
		.dout(new_net_4489)
	);

	bfr new_net_4491_bfr_before (
		.din(new_net_4491),
		.dout(new_net_4490)
	);

	bfr new_net_4492_bfr_before (
		.din(new_net_4492),
		.dout(new_net_4491)
	);

	bfr new_net_4493_bfr_before (
		.din(new_net_4493),
		.dout(new_net_4492)
	);

	bfr new_net_4494_bfr_before (
		.din(new_net_4494),
		.dout(new_net_4493)
	);

	bfr new_net_4495_bfr_before (
		.din(new_net_4495),
		.dout(new_net_4494)
	);

	bfr new_net_4496_bfr_before (
		.din(new_net_4496),
		.dout(new_net_4495)
	);

	bfr new_net_4497_bfr_before (
		.din(new_net_4497),
		.dout(new_net_4496)
	);

	bfr new_net_4498_bfr_before (
		.din(new_net_4498),
		.dout(new_net_4497)
	);

	bfr new_net_4499_bfr_before (
		.din(new_net_4499),
		.dout(new_net_4498)
	);

	bfr new_net_4500_bfr_before (
		.din(new_net_4500),
		.dout(new_net_4499)
	);

	bfr new_net_4501_bfr_before (
		.din(new_net_4501),
		.dout(new_net_4500)
	);

	spl2 G152_v_fanout (
		.a(G152),
		.b(new_net_1340),
		.c(new_net_4501)
	);

	bfr new_net_4502_bfr_before (
		.din(new_net_4502),
		.dout(new_net_1789)
	);

	bfr new_net_4503_bfr_before (
		.din(new_net_4503),
		.dout(new_net_4502)
	);

	bfr new_net_4504_bfr_before (
		.din(new_net_4504),
		.dout(new_net_4503)
	);

	bfr new_net_4505_bfr_before (
		.din(new_net_4505),
		.dout(new_net_4504)
	);

	bfr new_net_4506_bfr_before (
		.din(new_net_4506),
		.dout(new_net_4505)
	);

	bfr new_net_4507_bfr_before (
		.din(new_net_4507),
		.dout(new_net_4506)
	);

	bfr new_net_4508_bfr_before (
		.din(new_net_4508),
		.dout(new_net_4507)
	);

	bfr new_net_4509_bfr_before (
		.din(new_net_4509),
		.dout(new_net_4508)
	);

	bfr new_net_4510_bfr_before (
		.din(new_net_4510),
		.dout(new_net_4509)
	);

	bfr new_net_4511_bfr_before (
		.din(new_net_4511),
		.dout(new_net_4510)
	);

	bfr new_net_4512_bfr_before (
		.din(new_net_4512),
		.dout(new_net_4511)
	);

	bfr new_net_4513_bfr_before (
		.din(new_net_4513),
		.dout(new_net_4512)
	);

	bfr new_net_4514_bfr_before (
		.din(new_net_4514),
		.dout(new_net_4513)
	);

	spl3L G174_v_fanout (
		.a(G174),
		.b(new_net_929),
		.c(new_net_947),
		.d(new_net_4514)
	);

	bfr new_net_4515_bfr_before (
		.din(new_net_4515),
		.dout(new_net_1801)
	);

	bfr new_net_4516_bfr_before (
		.din(new_net_4516),
		.dout(new_net_4515)
	);

	bfr new_net_4517_bfr_before (
		.din(new_net_4517),
		.dout(new_net_4516)
	);

	bfr new_net_4518_bfr_before (
		.din(new_net_4518),
		.dout(new_net_4517)
	);

	spl2 G170_v_fanout (
		.a(G170),
		.b(new_net_4518),
		.c(new_net_590)
	);

	bfr new_net_4519_bfr_after (
		.din(G77),
		.dout(new_net_4519)
	);

	bfr new_net_4520_bfr_after (
		.din(new_net_4519),
		.dout(new_net_4520)
	);

	bfr new_net_4521_bfr_after (
		.din(new_net_4520),
		.dout(new_net_4521)
	);

	spl2 G77_v_fanout (
		.a(new_net_4521),
		.b(new_net_1437),
		.c(new_net_1438)
	);

	bfr new_net_4522_bfr_after (
		.din(G76),
		.dout(new_net_4522)
	);

	bfr new_net_4523_bfr_after (
		.din(new_net_4522),
		.dout(new_net_4523)
	);

	bfr new_net_4524_bfr_after (
		.din(new_net_4523),
		.dout(new_net_4524)
	);

	spl2 G76_v_fanout (
		.a(new_net_4524),
		.b(new_net_1425),
		.c(new_net_1426)
	);

	spl3L G101_v_fanout (
		.a(G101),
		.b(new_net_1805),
		.c(new_net_1806),
		.d(new_net_1807)
	);

	bfr new_net_4525_bfr_after (
		.din(G40),
		.dout(new_net_4525)
	);

	bfr new_net_4526_bfr_after (
		.din(new_net_4525),
		.dout(new_net_4526)
	);

	bfr new_net_4527_bfr_after (
		.din(new_net_4526),
		.dout(new_net_4527)
	);

	spl2 G40_v_fanout (
		.a(new_net_4527),
		.b(new_net_696),
		.c(new_net_697)
	);

	spl2 G11_v_fanout (
		.a(G11),
		.b(new_net_1271),
		.c(new_net_1272)
	);

	spl2 G153_v_fanout (
		.a(G153),
		.b(new_net_208),
		.c(new_net_209)
	);

	bfr new_net_4528_bfr_after (
		.din(G171),
		.dout(new_net_4528)
	);

	bfr new_net_4529_bfr_after (
		.din(new_net_4528),
		.dout(new_net_4529)
	);

	bfr new_net_4530_bfr_after (
		.din(new_net_4529),
		.dout(new_net_4530)
	);

	bfr new_net_4531_bfr_after (
		.din(new_net_4530),
		.dout(new_net_4531)
	);

	bfr new_net_4532_bfr_after (
		.din(new_net_4531),
		.dout(new_net_4532)
	);

	bfr new_net_4533_bfr_after (
		.din(new_net_4532),
		.dout(new_net_4533)
	);

	bfr new_net_4534_bfr_after (
		.din(new_net_4533),
		.dout(new_net_4534)
	);

	bfr new_net_4535_bfr_before (
		.din(new_net_4535),
		.dout(new_net_129)
	);

	bfr new_net_4536_bfr_before (
		.din(new_net_4536),
		.dout(new_net_4535)
	);

	bfr new_net_4537_bfr_before (
		.din(new_net_4537),
		.dout(new_net_4536)
	);

	bfr new_net_4538_bfr_before (
		.din(new_net_4538),
		.dout(new_net_4537)
	);

	bfr new_net_4539_bfr_before (
		.din(new_net_4539),
		.dout(new_net_4538)
	);

	bfr new_net_4540_bfr_before (
		.din(new_net_4540),
		.dout(new_net_4539)
	);

	spl2 G171_v_fanout (
		.a(new_net_4534),
		.b(new_net_4540),
		.c(new_net_130)
	);

	bfr new_net_4541_bfr_after (
		.din(G22),
		.dout(new_net_4541)
	);

	bfr new_net_4542_bfr_after (
		.din(new_net_4541),
		.dout(new_net_4542)
	);

	bfr new_net_4543_bfr_after (
		.din(new_net_4542),
		.dout(new_net_4543)
	);

	spl2 G22_v_fanout (
		.a(new_net_4543),
		.b(new_net_352),
		.c(new_net_353)
	);

	bfr new_net_4544_bfr_before (
		.din(new_net_4544),
		.dout(new_net_1810)
	);

	spl2 G103_v_fanout (
		.a(G103),
		.b(new_net_1811),
		.c(new_net_4544)
	);

	bfr new_net_4545_bfr_before (
		.din(new_net_4545),
		.dout(new_net_1812)
	);

	bfr new_net_4546_bfr_before (
		.din(new_net_4546),
		.dout(new_net_4545)
	);

	bfr new_net_4547_bfr_before (
		.din(new_net_4547),
		.dout(new_net_4546)
	);

	spl2 G143_v_fanout (
		.a(G143),
		.b(new_net_770),
		.c(new_net_4547)
	);

	bfr new_net_4548_bfr_after (
		.din(G14),
		.dout(new_net_4548)
	);

	bfr new_net_4549_bfr_after (
		.din(new_net_4548),
		.dout(new_net_4549)
	);

	bfr new_net_4550_bfr_after (
		.din(new_net_4549),
		.dout(new_net_4550)
	);

	spl2 G14_v_fanout (
		.a(new_net_4550),
		.b(new_net_1022),
		.c(new_net_1023)
	);

	spl2 G90_v_fanout (
		.a(G90),
		.b(new_net_1815),
		.c(new_net_1816)
	);

	bfr new_net_4551_bfr_before (
		.din(new_net_4551),
		.dout(new_net_1708)
	);

	bfr new_net_4552_bfr_before (
		.din(new_net_4552),
		.dout(new_net_4551)
	);

	spl2 G129_v_fanout (
		.a(G129),
		.b(new_net_1707),
		.c(new_net_4552)
	);

	bfr new_net_4553_bfr_after (
		.din(G26),
		.dout(new_net_4553)
	);

	bfr new_net_4554_bfr_after (
		.din(new_net_4553),
		.dout(new_net_4554)
	);

	bfr new_net_4555_bfr_after (
		.din(new_net_4554),
		.dout(new_net_4555)
	);

	spl2 G26_v_fanout (
		.a(new_net_4555),
		.b(new_net_450),
		.c(new_net_451)
	);

	bfr new_net_4556_bfr_before (
		.din(new_net_4556),
		.dout(new_net_1817)
	);

	bfr new_net_4557_bfr_before (
		.din(new_net_4557),
		.dout(new_net_4556)
	);

	bfr new_net_4558_bfr_before (
		.din(new_net_4558),
		.dout(new_net_4557)
	);

	bfr new_net_4559_bfr_before (
		.din(new_net_4559),
		.dout(new_net_4558)
	);

	bfr new_net_4560_bfr_before (
		.din(new_net_4560),
		.dout(new_net_4559)
	);

	bfr new_net_4561_bfr_before (
		.din(new_net_4561),
		.dout(new_net_4560)
	);

	bfr new_net_4562_bfr_before (
		.din(new_net_4562),
		.dout(new_net_4561)
	);

	bfr new_net_4563_bfr_before (
		.din(new_net_4563),
		.dout(new_net_4562)
	);

	bfr new_net_4564_bfr_before (
		.din(new_net_4564),
		.dout(new_net_4563)
	);

	bfr new_net_4565_bfr_before (
		.din(new_net_4565),
		.dout(new_net_4564)
	);

	bfr new_net_4566_bfr_before (
		.din(new_net_4566),
		.dout(new_net_4565)
	);

	bfr new_net_4567_bfr_before (
		.din(new_net_4567),
		.dout(new_net_4566)
	);

	bfr new_net_4568_bfr_before (
		.din(new_net_4568),
		.dout(new_net_4567)
	);

	bfr new_net_4569_bfr_before (
		.din(new_net_4569),
		.dout(new_net_4568)
	);

	bfr new_net_4570_bfr_before (
		.din(new_net_4570),
		.dout(new_net_4569)
	);

	bfr new_net_4571_bfr_before (
		.din(new_net_4571),
		.dout(new_net_4570)
	);

	bfr new_net_4572_bfr_before (
		.din(new_net_4572),
		.dout(new_net_4571)
	);

	spl4L G158_v_fanout (
		.a(G158),
		.b(new_net_664),
		.c(new_net_665),
		.d(new_net_4572),
		.e(new_net_662)
	);

	spl4L G124_v_fanout (
		.a(G124),
		.b(new_net_1829),
		.c(new_net_1828),
		.d(new_net_1830),
		.e(new_net_1827)
	);

	bfr new_net_4573_bfr_after (
		.din(G70),
		.dout(new_net_4573)
	);

	bfr new_net_4574_bfr_after (
		.din(new_net_4573),
		.dout(new_net_4574)
	);

	bfr new_net_4575_bfr_after (
		.din(new_net_4574),
		.dout(new_net_4575)
	);

	spl2 G70_v_fanout (
		.a(new_net_4575),
		.b(new_net_745),
		.c(new_net_746)
	);

	bfr new_net_4576_bfr_after (
		.din(G15),
		.dout(new_net_4576)
	);

	bfr new_net_4577_bfr_after (
		.din(new_net_4576),
		.dout(new_net_4577)
	);

	bfr new_net_4578_bfr_after (
		.din(new_net_4577),
		.dout(new_net_4578)
	);

	spl2 G15_v_fanout (
		.a(new_net_4578),
		.b(new_net_1458),
		.c(new_net_1459)
	);

	bfr new_net_4579_bfr_after (
		.din(G80),
		.dout(new_net_4579)
	);

	bfr new_net_4580_bfr_after (
		.din(new_net_4579),
		.dout(new_net_4580)
	);

	bfr new_net_4581_bfr_after (
		.din(new_net_4580),
		.dout(new_net_4581)
	);

	spl2 G80_v_fanout (
		.a(new_net_4581),
		.b(new_net_1542),
		.c(new_net_1543)
	);

	bfr new_net_4582_bfr_after (
		.din(G24),
		.dout(new_net_4582)
	);

	bfr new_net_4583_bfr_after (
		.din(new_net_4582),
		.dout(new_net_4583)
	);

	bfr new_net_4584_bfr_after (
		.din(new_net_4583),
		.dout(new_net_4584)
	);

	spl2 G24_v_fanout (
		.a(new_net_4584),
		.b(new_net_403),
		.c(new_net_404)
	);

	spl3L G161_v_fanout (
		.a(G161),
		.b(new_net_1532),
		.c(new_net_1534),
		.d(new_net_1533)
	);

	bfr new_net_4585_bfr_after (
		.din(G81),
		.dout(new_net_4585)
	);

	bfr new_net_4586_bfr_after (
		.din(new_net_4585),
		.dout(new_net_4586)
	);

	bfr new_net_4587_bfr_after (
		.din(new_net_4586),
		.dout(new_net_4587)
	);

	spl2 G81_v_fanout (
		.a(new_net_4587),
		.b(new_net_1583),
		.c(new_net_1584)
	);

	bfr new_net_4588_bfr_before (
		.din(new_net_4588),
		.dout(new_net_906)
	);

	bfr new_net_4589_bfr_before (
		.din(new_net_4589),
		.dout(new_net_4588)
	);

	bfr new_net_4590_bfr_before (
		.din(new_net_4590),
		.dout(new_net_4589)
	);

	bfr new_net_4591_bfr_before (
		.din(new_net_4591),
		.dout(new_net_4590)
	);

	spl2 G54_v_fanout (
		.a(G54),
		.b(new_net_4591),
		.c(new_net_907)
	);

	bfr new_net_4592_bfr_before (
		.din(new_net_4592),
		.dout(new_net_852)
	);

	bfr new_net_4593_bfr_before (
		.din(new_net_4593),
		.dout(new_net_4592)
	);

	spl3L G132_v_fanout (
		.a(G132),
		.b(new_net_851),
		.c(new_net_4593),
		.d(new_net_853)
	);

	bfr new_net_4594_bfr_before (
		.din(new_net_4594),
		.dout(new_net_1831)
	);

	bfr new_net_4595_bfr_before (
		.din(new_net_4595),
		.dout(new_net_4594)
	);

	bfr new_net_4596_bfr_before (
		.din(new_net_4596),
		.dout(new_net_4595)
	);

	spl2 G142_v_fanout (
		.a(G142),
		.b(new_net_4596),
		.c(new_net_1095)
	);

	bfr new_net_4597_bfr_before (
		.din(new_net_4597),
		.dout(new_net_1832)
	);

	bfr new_net_4598_bfr_before (
		.din(new_net_4598),
		.dout(new_net_4597)
	);

	bfr new_net_4599_bfr_before (
		.din(new_net_4599),
		.dout(new_net_4598)
	);

	spl2 G150_v_fanout (
		.a(G150),
		.b(new_net_1592),
		.c(new_net_4599)
	);

	bfr new_net_4600_bfr_after (
		.din(G78),
		.dout(new_net_4600)
	);

	bfr new_net_4601_bfr_after (
		.din(new_net_4600),
		.dout(new_net_4601)
	);

	bfr new_net_4602_bfr_after (
		.din(new_net_4601),
		.dout(new_net_4602)
	);

	spl2 G78_v_fanout (
		.a(new_net_4602),
		.b(new_net_1478),
		.c(new_net_1479)
	);

	bfr new_net_4603_bfr_before (
		.din(new_net_4603),
		.dout(new_net_848)
	);

	bfr new_net_4604_bfr_before (
		.din(new_net_4604),
		.dout(new_net_4603)
	);

	spl2 G131_v_fanout (
		.a(G131),
		.b(new_net_847),
		.c(new_net_4604)
	);

	spl3L G130_v_fanout (
		.a(G130),
		.b(new_net_1833),
		.c(new_net_1030),
		.d(new_net_1034)
	);

	spl2 G113_v_fanout (
		.a(G113),
		.b(new_net_1834),
		.c(new_net_1835)
	);

	spl2 G92_v_fanout (
		.a(G92),
		.b(new_net_1839),
		.c(new_net_1838)
	);

	bfr new_net_4605_bfr_before (
		.din(new_net_4605),
		.dout(new_net_1840)
	);

	bfr new_net_4606_bfr_before (
		.din(new_net_4606),
		.dout(new_net_4605)
	);

	bfr new_net_4607_bfr_before (
		.din(new_net_4607),
		.dout(new_net_4606)
	);

	bfr new_net_4608_bfr_before (
		.din(new_net_4608),
		.dout(new_net_4607)
	);

	bfr new_net_4609_bfr_before (
		.din(new_net_4609),
		.dout(new_net_4608)
	);

	spl2 G145_v_fanout (
		.a(G145),
		.b(new_net_4609),
		.c(new_net_905)
	);

	bfr new_net_4610_bfr_after (
		.din(G23),
		.dout(new_net_4610)
	);

	bfr new_net_4611_bfr_after (
		.din(new_net_4610),
		.dout(new_net_4611)
	);

	bfr new_net_4612_bfr_after (
		.din(new_net_4611),
		.dout(new_net_4612)
	);

	spl2 G23_v_fanout (
		.a(new_net_4612),
		.b(new_net_374),
		.c(new_net_375)
	);

	bfr new_net_4613_bfr_after (
		.din(G3),
		.dout(new_net_4613)
	);

	bfr new_net_4614_bfr_after (
		.din(new_net_4613),
		.dout(new_net_4614)
	);

	bfr new_net_4615_bfr_after (
		.din(new_net_4614),
		.dout(new_net_4615)
	);

	spl2 G3_v_fanout (
		.a(new_net_4615),
		.b(new_net_505),
		.c(new_net_506)
	);

	spl2 G102_v_fanout (
		.a(G102),
		.b(new_net_1845),
		.c(new_net_1844)
	);

	bfr new_net_4616_bfr_before (
		.din(new_net_4616),
		.dout(new_net_1848)
	);

	spl2 G107_v_fanout (
		.a(G107),
		.b(new_net_4616),
		.c(new_net_1849)
	);

	bfr new_net_4617_bfr_after (
		.din(G17),
		.dout(new_net_4617)
	);

	bfr new_net_4618_bfr_after (
		.din(new_net_4617),
		.dout(new_net_4618)
	);

	bfr new_net_4619_bfr_after (
		.din(new_net_4618),
		.dout(new_net_4619)
	);

	spl2 G17_v_fanout (
		.a(new_net_4619),
		.b(new_net_523),
		.c(new_net_524)
	);

	spl2 G166_v_fanout (
		.a(G166),
		.b(new_net_1852),
		.c(new_net_1853)
	);

	bfr new_net_4620_bfr_before (
		.din(new_net_4620),
		.dout(new_net_1854)
	);

	bfr new_net_4621_bfr_before (
		.din(new_net_4621),
		.dout(new_net_4620)
	);

	bfr new_net_4622_bfr_before (
		.din(new_net_4622),
		.dout(new_net_4621)
	);

	bfr new_net_4623_bfr_before (
		.din(new_net_4623),
		.dout(new_net_4622)
	);

	bfr new_net_4624_bfr_before (
		.din(new_net_4624),
		.dout(new_net_4623)
	);

	bfr new_net_4625_bfr_before (
		.din(new_net_4625),
		.dout(new_net_4624)
	);

	bfr new_net_4626_bfr_before (
		.din(new_net_4626),
		.dout(new_net_4625)
	);

	bfr new_net_4627_bfr_before (
		.din(new_net_4627),
		.dout(new_net_4626)
	);

	bfr new_net_4628_bfr_before (
		.din(new_net_4628),
		.dout(new_net_4627)
	);

	bfr new_net_4629_bfr_before (
		.din(new_net_4629),
		.dout(new_net_4628)
	);

	bfr new_net_4630_bfr_before (
		.din(new_net_4630),
		.dout(new_net_4629)
	);

	bfr new_net_4631_bfr_before (
		.din(new_net_4631),
		.dout(new_net_4630)
	);

	bfr new_net_4632_bfr_before (
		.din(new_net_4632),
		.dout(new_net_4631)
	);

	bfr new_net_4633_bfr_before (
		.din(new_net_4633),
		.dout(new_net_4632)
	);

	bfr new_net_4634_bfr_before (
		.din(new_net_4634),
		.dout(new_net_4633)
	);

	bfr new_net_4635_bfr_before (
		.din(new_net_4635),
		.dout(new_net_4634)
	);

	bfr new_net_4636_bfr_before (
		.din(new_net_4636),
		.dout(new_net_4635)
	);

	bfr new_net_4637_bfr_before (
		.din(new_net_4637),
		.dout(new_net_4636)
	);

	bfr new_net_4638_bfr_before (
		.din(new_net_4638),
		.dout(new_net_4637)
	);

	bfr new_net_4639_bfr_before (
		.din(new_net_4639),
		.dout(new_net_4638)
	);

	spl2 G64_v_fanout (
		.a(G64),
		.b(new_net_4639),
		.c(new_net_122)
	);

	bfr new_net_4640_bfr_before (
		.din(new_net_4640),
		.dout(new_net_1863)
	);

	bfr new_net_4641_bfr_before (
		.din(new_net_4641),
		.dout(new_net_4640)
	);

	spl2 G140_v_fanout (
		.a(G140),
		.b(new_net_1053),
		.c(new_net_4641)
	);

	bfr new_net_4642_bfr_before (
		.din(new_net_4642),
		.dout(new_net_1864)
	);

	bfr new_net_4643_bfr_before (
		.din(new_net_4643),
		.dout(new_net_4642)
	);

	bfr new_net_4644_bfr_before (
		.din(new_net_4644),
		.dout(new_net_4643)
	);

	bfr new_net_4645_bfr_before (
		.din(new_net_4645),
		.dout(new_net_4644)
	);

	bfr new_net_4646_bfr_before (
		.din(new_net_4646),
		.dout(new_net_4645)
	);

	bfr new_net_4647_bfr_before (
		.din(new_net_4647),
		.dout(new_net_4646)
	);

	bfr new_net_4648_bfr_before (
		.din(new_net_4648),
		.dout(new_net_4647)
	);

	bfr new_net_4649_bfr_before (
		.din(new_net_4649),
		.dout(new_net_4648)
	);

	bfr new_net_4650_bfr_before (
		.din(new_net_4650),
		.dout(new_net_4649)
	);

	bfr new_net_4651_bfr_before (
		.din(new_net_4651),
		.dout(new_net_4650)
	);

	bfr new_net_4652_bfr_before (
		.din(new_net_4652),
		.dout(new_net_4651)
	);

	bfr new_net_4653_bfr_before (
		.din(new_net_4653),
		.dout(new_net_4652)
	);

	bfr new_net_4654_bfr_before (
		.din(new_net_4654),
		.dout(new_net_4653)
	);

	bfr new_net_4655_bfr_before (
		.din(new_net_4655),
		.dout(new_net_4654)
	);

	bfr new_net_4656_bfr_before (
		.din(new_net_4656),
		.dout(new_net_4655)
	);

	bfr new_net_4657_bfr_before (
		.din(new_net_4657),
		.dout(new_net_4656)
	);

	bfr new_net_4658_bfr_before (
		.din(new_net_4658),
		.dout(new_net_4657)
	);

	bfr new_net_4659_bfr_before (
		.din(new_net_4659),
		.dout(new_net_4658)
	);

	bfr new_net_4660_bfr_before (
		.din(new_net_4660),
		.dout(new_net_4659)
	);

	bfr new_net_4661_bfr_before (
		.din(new_net_4661),
		.dout(new_net_4660)
	);

	bfr new_net_4662_bfr_before (
		.din(new_net_4662),
		.dout(new_net_4661)
	);

	bfr new_net_4663_bfr_before (
		.din(new_net_4663),
		.dout(new_net_4662)
	);

	bfr new_net_4664_bfr_before (
		.din(new_net_4664),
		.dout(new_net_4663)
	);

	bfr new_net_4665_bfr_before (
		.din(new_net_4665),
		.dout(new_net_4664)
	);

	bfr new_net_4666_bfr_before (
		.din(new_net_4666),
		.dout(new_net_4665)
	);

	bfr new_net_4667_bfr_before (
		.din(new_net_4667),
		.dout(new_net_4666)
	);

	bfr new_net_4668_bfr_before (
		.din(new_net_4668),
		.dout(new_net_4667)
	);

	bfr new_net_4669_bfr_before (
		.din(new_net_4669),
		.dout(new_net_4668)
	);

	bfr new_net_4670_bfr_before (
		.din(new_net_4670),
		.dout(new_net_4669)
	);

	spl4L G173_v_fanout (
		.a(G173),
		.b(new_net_149),
		.c(new_net_147),
		.d(new_net_4670),
		.e(new_net_146)
	);

	bfr new_net_4671_bfr_before (
		.din(new_net_4671),
		.dout(new_net_1269)
	);

	bfr new_net_4672_bfr_before (
		.din(new_net_4672),
		.dout(new_net_1270)
	);

	spl3L G148_v_fanout (
		.a(G148),
		.b(new_net_4671),
		.c(new_net_4672),
		.d(new_net_1867)
	);

	bfr new_net_4673_bfr_before (
		.din(new_net_4673),
		.dout(new_net_1871)
	);

	spl2 G128_v_fanout (
		.a(G128),
		.b(new_net_1872),
		.c(new_net_4673)
	);

	spl2 G98_v_fanout (
		.a(G98),
		.b(new_net_1877),
		.c(new_net_1876)
	);

	bfr new_net_4674_bfr_after (
		.din(G36),
		.dout(new_net_4674)
	);

	bfr new_net_4675_bfr_after (
		.din(new_net_4674),
		.dout(new_net_4675)
	);

	bfr new_net_4676_bfr_after (
		.din(new_net_4675),
		.dout(new_net_4676)
	);

	spl2 G36_v_fanout (
		.a(new_net_4676),
		.b(new_net_165),
		.c(new_net_166)
	);

	bfr new_net_4677_bfr_after (
		.din(G6),
		.dout(new_net_4677)
	);

	bfr new_net_4678_bfr_after (
		.din(new_net_4677),
		.dout(new_net_4678)
	);

	bfr new_net_4679_bfr_after (
		.din(new_net_4678),
		.dout(new_net_4679)
	);

	spl2 G6_v_fanout (
		.a(new_net_4679),
		.b(new_net_1064),
		.c(new_net_1065)
	);

	bfr new_net_4680_bfr_before (
		.din(new_net_4680),
		.dout(new_net_1878)
	);

	spl2 G114_v_fanout (
		.a(G114),
		.b(new_net_4680),
		.c(new_net_1338)
	);

	bfr new_net_4681_bfr_before (
		.din(new_net_4681),
		.dout(new_net_958)
	);

	spl4L G94_v_fanout (
		.a(G94),
		.b(new_net_1880),
		.c(new_net_1879),
		.d(new_net_1881),
		.e(new_net_4681)
	);

	bfr new_net_4682_bfr_before (
		.din(new_net_4682),
		.dout(new_net_1882)
	);

	bfr new_net_4683_bfr_before (
		.din(new_net_4683),
		.dout(new_net_4682)
	);

	bfr new_net_4684_bfr_before (
		.din(new_net_4684),
		.dout(new_net_4683)
	);

	spl2 G144_v_fanout (
		.a(G144),
		.b(new_net_4684),
		.c(new_net_825)
	);

	spl2 G169_v_fanout (
		.a(G169),
		.b(new_net_1886),
		.c(new_net_1887)
	);

	bfr new_net_4685_bfr_after (
		.din(G83),
		.dout(new_net_4685)
	);

	bfr new_net_4686_bfr_after (
		.din(new_net_4685),
		.dout(new_net_4686)
	);

	bfr new_net_4687_bfr_after (
		.din(new_net_4686),
		.dout(new_net_4687)
	);

	spl2 G83_v_fanout (
		.a(new_net_4687),
		.b(new_net_1622),
		.c(new_net_1623)
	);

	spl3L G163_v_fanout (
		.a(G163),
		.b(new_net_1888),
		.c(new_net_1889),
		.d(new_net_1890)
	);

	spl3L G126_v_fanout (
		.a(G126),
		.b(new_net_1893),
		.c(new_net_1891),
		.d(new_net_1892)
	);

	bfr new_net_4688_bfr_after (
		.din(G79),
		.dout(new_net_4688)
	);

	bfr new_net_4689_bfr_after (
		.din(new_net_4688),
		.dout(new_net_4689)
	);

	bfr new_net_4690_bfr_after (
		.din(new_net_4689),
		.dout(new_net_4690)
	);

	spl2 G79_v_fanout (
		.a(new_net_4690),
		.b(new_net_1717),
		.c(new_net_1718)
	);

	bfr new_net_4691_bfr_before (
		.din(new_net_4691),
		.dout(new_net_1894)
	);

	bfr new_net_4692_bfr_before (
		.din(new_net_4692),
		.dout(new_net_4691)
	);

	bfr new_net_4693_bfr_before (
		.din(new_net_4693),
		.dout(new_net_4692)
	);

	bfr new_net_4694_bfr_before (
		.din(new_net_4694),
		.dout(new_net_4693)
	);

	bfr new_net_4695_bfr_before (
		.din(new_net_4695),
		.dout(new_net_4694)
	);

	bfr new_net_4696_bfr_before (
		.din(new_net_4696),
		.dout(new_net_4695)
	);

	bfr new_net_4697_bfr_before (
		.din(new_net_4697),
		.dout(new_net_4696)
	);

	bfr new_net_4698_bfr_before (
		.din(new_net_4698),
		.dout(new_net_4697)
	);

	bfr new_net_4699_bfr_before (
		.din(new_net_4699),
		.dout(new_net_4698)
	);

	bfr new_net_4700_bfr_before (
		.din(new_net_4700),
		.dout(new_net_4699)
	);

	bfr new_net_4701_bfr_before (
		.din(new_net_4701),
		.dout(new_net_4700)
	);

	bfr new_net_4702_bfr_before (
		.din(new_net_4702),
		.dout(new_net_4701)
	);

	bfr new_net_4703_bfr_before (
		.din(new_net_4703),
		.dout(new_net_4702)
	);

	bfr new_net_4704_bfr_before (
		.din(new_net_4704),
		.dout(new_net_4703)
	);

	bfr new_net_4705_bfr_before (
		.din(new_net_4705),
		.dout(new_net_4704)
	);

	bfr new_net_4706_bfr_before (
		.din(new_net_4706),
		.dout(new_net_4705)
	);

	bfr new_net_4707_bfr_before (
		.din(new_net_4707),
		.dout(new_net_4706)
	);

	spl4L G160_v_fanout (
		.a(G160),
		.b(new_net_1495),
		.c(new_net_1494),
		.d(new_net_4707),
		.e(new_net_1493)
	);

	bfr new_net_4708_bfr_before (
		.din(new_net_4708),
		.dout(new_net_1901)
	);

	bfr new_net_4709_bfr_before (
		.din(new_net_4709),
		.dout(new_net_4708)
	);

	bfr new_net_4710_bfr_before (
		.din(new_net_4710),
		.dout(new_net_4709)
	);

	bfr new_net_4711_bfr_before (
		.din(new_net_4711),
		.dout(new_net_4710)
	);

	spl2 G138_v_fanout (
		.a(G138),
		.b(new_net_4711),
		.c(new_net_963)
	);

	spl3L G175_v_fanout (
		.a(G175),
		.b(new_net_1087),
		.c(new_net_1088),
		.d(new_net_1089)
	);

	bfr new_net_4712_bfr_after (
		.din(G84),
		.dout(new_net_4712)
	);

	bfr new_net_4713_bfr_after (
		.din(new_net_4712),
		.dout(new_net_4713)
	);

	bfr new_net_4714_bfr_after (
		.din(new_net_4713),
		.dout(new_net_4714)
	);

	spl2 G84_v_fanout (
		.a(new_net_4714),
		.b(new_net_1653),
		.c(new_net_1654)
	);

	bfr new_net_4715_bfr_after (
		.din(G74),
		.dout(new_net_4715)
	);

	bfr new_net_4716_bfr_after (
		.din(new_net_4715),
		.dout(new_net_4716)
	);

	bfr new_net_4717_bfr_after (
		.din(new_net_4716),
		.dout(new_net_4717)
	);

	spl2 G74_v_fanout (
		.a(new_net_4717),
		.b(new_net_1135),
		.c(new_net_1136)
	);

	spl4L G177_v_fanout (
		.a(G177),
		.b(new_net_221),
		.c(new_net_223),
		.d(new_net_222),
		.e(new_net_220)
	);

	spl2 G115_v_fanout (
		.a(G115),
		.b(new_net_1902),
		.c(new_net_1903)
	);

	bfr new_net_4718_bfr_after (
		.din(G16),
		.dout(new_net_4718)
	);

	bfr new_net_4719_bfr_after (
		.din(new_net_4718),
		.dout(new_net_4719)
	);

	bfr new_net_4720_bfr_after (
		.din(new_net_4719),
		.dout(new_net_4720)
	);

	spl2 G16_v_fanout (
		.a(new_net_4720),
		.b(new_net_1476),
		.c(new_net_1477)
	);

	spl3L G172_v_fanout (
		.a(G172),
		.b(new_net_141),
		.c(new_net_142),
		.d(new_net_143)
	);

	spl2 G99_v_fanout (
		.a(G99),
		.b(new_net_1439),
		.c(new_net_1440)
	);

	bfr new_net_4721_bfr_before (
		.din(new_net_4721),
		.dout(G5216)
	);

	bfr new_net_4722_bfr_before (
		.din(new_net_4722),
		.dout(new_net_4721)
	);

	bfr new_net_4723_bfr_before (
		.din(new_net_4723),
		.dout(new_net_4722)
	);

	bfr new_net_4724_bfr_before (
		.din(new_net_4724),
		.dout(new_net_4723)
	);

	bfr new_net_4725_bfr_before (
		.din(new_net_4725),
		.dout(new_net_4724)
	);

	bfr new_net_4726_bfr_before (
		.din(new_net_4726),
		.dout(new_net_4725)
	);

	bfr new_net_4727_bfr_before (
		.din(new_net_4727),
		.dout(new_net_4726)
	);

	bfr new_net_4728_bfr_before (
		.din(new_net_4728),
		.dout(new_net_4727)
	);

	bfr new_net_4729_bfr_before (
		.din(new_net_4729),
		.dout(new_net_4728)
	);

	bfr new_net_4730_bfr_before (
		.din(new_net_4730),
		.dout(new_net_4729)
	);

	bfr new_net_4731_bfr_before (
		.din(new_net_4731),
		.dout(new_net_4730)
	);

	bfr new_net_4732_bfr_before (
		.din(new_net_4732),
		.dout(new_net_4731)
	);

	bfr new_net_4733_bfr_before (
		.din(new_net_4733),
		.dout(new_net_4732)
	);

	bfr new_net_4734_bfr_before (
		.din(new_net_4734),
		.dout(new_net_4733)
	);

	bfr new_net_4735_bfr_before (
		.din(new_net_4735),
		.dout(new_net_4734)
	);

	bfr new_net_4736_bfr_before (
		.din(new_net_4736),
		.dout(new_net_4735)
	);

	bfr new_net_4737_bfr_before (
		.din(new_net_4737),
		.dout(new_net_4736)
	);

	bfr new_net_4738_bfr_before (
		.din(new_net_4738),
		.dout(new_net_4737)
	);

	bfr new_net_4739_bfr_before (
		.din(new_net_4739),
		.dout(new_net_4738)
	);

	bfr new_net_4740_bfr_before (
		.din(new_net_4740),
		.dout(new_net_4739)
	);

	bfr new_net_4741_bfr_before (
		.din(new_net_4741),
		.dout(new_net_4740)
	);

	bfr new_net_4742_bfr_before (
		.din(new_net_4742),
		.dout(new_net_4741)
	);

	bfr new_net_4743_bfr_before (
		.din(new_net_4743),
		.dout(new_net_4742)
	);

	bfr new_net_4744_bfr_before (
		.din(new_net_4744),
		.dout(new_net_4743)
	);

	bfr new_net_4745_bfr_before (
		.din(new_net_4745),
		.dout(new_net_4744)
	);

	bfr new_net_4746_bfr_before (
		.din(new_net_4746),
		.dout(new_net_4745)
	);

	bfr new_net_4747_bfr_before (
		.din(new_net_4747),
		.dout(new_net_4746)
	);

	bfr new_net_4748_bfr_before (
		.din(new_net_4748),
		.dout(new_net_4747)
	);

	bfr new_net_4749_bfr_before (
		.din(new_net_4749),
		.dout(new_net_4748)
	);

	bfr new_net_4750_bfr_before (
		.din(new_net_4750),
		.dout(new_net_4749)
	);

	bfr new_net_4751_bfr_before (
		.din(new_net_4751),
		.dout(new_net_4750)
	);

	bfr new_net_4752_bfr_before (
		.din(new_net_4752),
		.dout(new_net_4751)
	);

	bfr new_net_4753_bfr_before (
		.din(new_net_4753),
		.dout(new_net_4752)
	);

	bfr new_net_4754_bfr_before (
		.din(new_net_4754),
		.dout(new_net_4753)
	);

	bfr new_net_4755_bfr_before (
		.din(new_net_4755),
		.dout(new_net_4754)
	);

	bfr new_net_4756_bfr_before (
		.din(new_net_4756),
		.dout(new_net_4755)
	);

	bfr new_net_4757_bfr_before (
		.din(new_net_4757),
		.dout(new_net_4756)
	);

	bfr new_net_4758_bfr_before (
		.din(new_net_4758),
		.dout(new_net_4757)
	);

	bfr new_net_4759_bfr_before (
		.din(new_net_4759),
		.dout(new_net_4758)
	);

	bfr new_net_4760_bfr_before (
		.din(new_net_4760),
		.dout(new_net_4759)
	);

	bfr new_net_4761_bfr_before (
		.din(new_net_4761),
		.dout(new_net_4760)
	);

	spl3L G1_v_fanout (
		.a(G1),
		.b(new_net_55),
		.c(new_net_4761),
		.d(new_net_57)
	);

	bfr new_net_4762_bfr_before (
		.din(new_net_4762),
		.dout(new_net_1904)
	);

	bfr new_net_4763_bfr_before (
		.din(new_net_4763),
		.dout(new_net_4762)
	);

	bfr new_net_4764_bfr_before (
		.din(new_net_4764),
		.dout(new_net_4763)
	);

	spl2 G137_v_fanout (
		.a(G137),
		.b(new_net_4764),
		.c(new_net_918)
	);

	bfr new_net_4765_bfr_after (
		.din(G42),
		.dout(new_net_4765)
	);

	bfr new_net_4766_bfr_after (
		.din(new_net_4765),
		.dout(new_net_4766)
	);

	bfr new_net_4767_bfr_after (
		.din(new_net_4766),
		.dout(new_net_4767)
	);

	spl2 G42_v_fanout (
		.a(new_net_4767),
		.b(new_net_794),
		.c(new_net_795)
	);

	spl2 G117_v_fanout (
		.a(G117),
		.b(new_net_1907),
		.c(new_net_1906)
	);

	bfr new_net_4768_bfr_after (
		.din(_0632_),
		.dout(new_net_4768)
	);

	bfr new_net_4769_bfr_after (
		.din(new_net_4768),
		.dout(new_net_4769)
	);

	bfr new_net_4770_bfr_after (
		.din(new_net_4769),
		.dout(new_net_4770)
	);

	bfr new_net_4771_bfr_after (
		.din(new_net_4770),
		.dout(new_net_4771)
	);

	bfr new_net_4772_bfr_after (
		.din(new_net_4771),
		.dout(new_net_4772)
	);

	bfr new_net_2125_bfr_after (
		.din(new_net_4772),
		.dout(new_net_2125)
	);

	bfr new_net_2146_bfr_after (
		.din(_0734_),
		.dout(new_net_2146)
	);

	bfr new_net_4773_bfr_after (
		.din(_0834_),
		.dout(new_net_4773)
	);

	bfr new_net_4774_bfr_after (
		.din(new_net_4773),
		.dout(new_net_4774)
	);

	bfr new_net_4775_bfr_after (
		.din(new_net_4774),
		.dout(new_net_4775)
	);

	bfr new_net_4776_bfr_after (
		.din(new_net_4775),
		.dout(new_net_4776)
	);

	bfr new_net_4777_bfr_after (
		.din(new_net_4776),
		.dout(new_net_4777)
	);

	bfr new_net_4778_bfr_after (
		.din(new_net_4777),
		.dout(new_net_4778)
	);

	bfr new_net_4779_bfr_after (
		.din(new_net_4778),
		.dout(new_net_4779)
	);

	bfr new_net_4780_bfr_after (
		.din(new_net_4779),
		.dout(new_net_4780)
	);

	bfr new_net_4781_bfr_after (
		.din(new_net_4780),
		.dout(new_net_4781)
	);

	bfr new_net_4782_bfr_after (
		.din(new_net_4781),
		.dout(new_net_4782)
	);

	bfr new_net_4783_bfr_after (
		.din(new_net_4782),
		.dout(new_net_4783)
	);

	bfr new_net_4784_bfr_after (
		.din(new_net_4783),
		.dout(new_net_4784)
	);

	bfr new_net_4785_bfr_after (
		.din(new_net_4784),
		.dout(new_net_4785)
	);

	bfr new_net_2167_bfr_after (
		.din(new_net_4785),
		.dout(new_net_2167)
	);

	bfr new_net_4786_bfr_after (
		.din(G95),
		.dout(new_net_4786)
	);

	bfr new_net_2188_bfr_after (
		.din(new_net_4786),
		.dout(new_net_2188)
	);

	bfr new_net_4787_bfr_after (
		.din(_0356_),
		.dout(new_net_4787)
	);

	bfr new_net_4788_bfr_after (
		.din(new_net_4787),
		.dout(new_net_4788)
	);

	bfr new_net_4789_bfr_after (
		.din(new_net_4788),
		.dout(new_net_4789)
	);

	bfr new_net_4790_bfr_after (
		.din(new_net_4789),
		.dout(new_net_4790)
	);

	bfr new_net_4791_bfr_after (
		.din(new_net_4790),
		.dout(new_net_4791)
	);

	bfr new_net_4792_bfr_after (
		.din(new_net_4791),
		.dout(new_net_4792)
	);

	bfr new_net_4793_bfr_after (
		.din(new_net_4792),
		.dout(new_net_4793)
	);

	bfr new_net_4794_bfr_after (
		.din(new_net_4793),
		.dout(new_net_4794)
	);

	bfr new_net_4795_bfr_after (
		.din(new_net_4794),
		.dout(new_net_4795)
	);

	bfr new_net_4796_bfr_after (
		.din(new_net_4795),
		.dout(new_net_4796)
	);

	bfr new_net_4797_bfr_after (
		.din(new_net_4796),
		.dout(new_net_4797)
	);

	bfr new_net_4798_bfr_after (
		.din(new_net_4797),
		.dout(new_net_4798)
	);

	bfr new_net_4799_bfr_after (
		.din(new_net_4798),
		.dout(new_net_4799)
	);

	bfr new_net_4800_bfr_after (
		.din(new_net_4799),
		.dout(new_net_4800)
	);

	bfr new_net_4801_bfr_after (
		.din(new_net_4800),
		.dout(new_net_4801)
	);

	bfr new_net_4802_bfr_after (
		.din(new_net_4801),
		.dout(new_net_4802)
	);

	bfr new_net_4803_bfr_after (
		.din(new_net_4802),
		.dout(new_net_4803)
	);

	bfr new_net_4804_bfr_after (
		.din(new_net_4803),
		.dout(new_net_4804)
	);

	bfr new_net_2293_bfr_after (
		.din(new_net_4804),
		.dout(new_net_2293)
	);

	bfr new_net_4805_bfr_after (
		.din(new_net_2429),
		.dout(new_net_4805)
	);

	bfr new_net_4806_bfr_after (
		.din(new_net_4805),
		.dout(new_net_4806)
	);

	bfr new_net_4807_bfr_after (
		.din(new_net_4806),
		.dout(new_net_4807)
	);

	bfr new_net_4808_bfr_after (
		.din(new_net_4807),
		.dout(new_net_4808)
	);

	bfr new_net_4809_bfr_after (
		.din(new_net_4808),
		.dout(new_net_4809)
	);

	bfr new_net_4810_bfr_after (
		.din(new_net_4809),
		.dout(new_net_4810)
	);

	bfr new_net_4811_bfr_after (
		.din(new_net_4810),
		.dout(new_net_4811)
	);

	bfr new_net_4812_bfr_after (
		.din(new_net_4811),
		.dout(new_net_4812)
	);

	bfr new_net_4813_bfr_after (
		.din(new_net_4812),
		.dout(new_net_4813)
	);

	bfr new_net_4814_bfr_after (
		.din(new_net_4813),
		.dout(new_net_4814)
	);

	bfr new_net_4815_bfr_after (
		.din(new_net_4814),
		.dout(new_net_4815)
	);

	bfr new_net_4816_bfr_after (
		.din(new_net_4815),
		.dout(new_net_4816)
	);

	bfr new_net_4817_bfr_after (
		.din(new_net_4816),
		.dout(new_net_4817)
	);

	bfr new_net_4818_bfr_after (
		.din(new_net_4817),
		.dout(new_net_4818)
	);

	bfr new_net_4819_bfr_after (
		.din(new_net_4818),
		.dout(new_net_4819)
	);

	bfr new_net_4820_bfr_after (
		.din(new_net_4819),
		.dout(new_net_4820)
	);

	bfr new_net_4821_bfr_after (
		.din(new_net_4820),
		.dout(new_net_4821)
	);

	bfr new_net_4822_bfr_after (
		.din(new_net_4821),
		.dout(new_net_4822)
	);

	bfr new_net_4823_bfr_after (
		.din(new_net_4822),
		.dout(new_net_4823)
	);

	bfr new_net_4824_bfr_after (
		.din(new_net_4823),
		.dout(new_net_4824)
	);

	bfr new_net_4825_bfr_after (
		.din(new_net_4824),
		.dout(new_net_4825)
	);

	bfr new_net_4826_bfr_after (
		.din(new_net_4825),
		.dout(new_net_4826)
	);

	bfr new_net_4827_bfr_after (
		.din(new_net_4826),
		.dout(new_net_4827)
	);

	bfr new_net_4828_bfr_after (
		.din(new_net_4827),
		.dout(new_net_4828)
	);

	bfr new_net_4829_bfr_after (
		.din(new_net_4828),
		.dout(new_net_4829)
	);

	bfr new_net_4830_bfr_after (
		.din(new_net_4829),
		.dout(new_net_4830)
	);

	bfr new_net_4831_bfr_after (
		.din(new_net_4830),
		.dout(new_net_4831)
	);

	bfr new_net_4832_bfr_after (
		.din(new_net_4831),
		.dout(new_net_4832)
	);

	bfr new_net_4833_bfr_after (
		.din(new_net_4832),
		.dout(new_net_4833)
	);

	bfr new_net_4834_bfr_after (
		.din(new_net_4833),
		.dout(new_net_4834)
	);

	bfr new_net_4835_bfr_after (
		.din(new_net_4834),
		.dout(new_net_4835)
	);

	bfr new_net_4836_bfr_after (
		.din(new_net_4835),
		.dout(new_net_4836)
	);

	bfr new_net_4837_bfr_after (
		.din(new_net_4836),
		.dout(new_net_4837)
	);

	bfr new_net_4838_bfr_after (
		.din(new_net_4837),
		.dout(new_net_4838)
	);

	bfr new_net_4839_bfr_after (
		.din(new_net_4838),
		.dout(new_net_4839)
	);

	bfr new_net_4840_bfr_after (
		.din(new_net_4839),
		.dout(new_net_4840)
	);

	bfr new_net_4841_bfr_after (
		.din(new_net_4840),
		.dout(new_net_4841)
	);

	bfr new_net_4842_bfr_after (
		.din(new_net_4841),
		.dout(new_net_4842)
	);

	bfr new_net_4843_bfr_after (
		.din(new_net_4842),
		.dout(new_net_4843)
	);

	bfr G5200_bfr_after (
		.din(new_net_4843),
		.dout(G5200)
	);

	bfr new_net_2209_bfr_after (
		.din(_1105_),
		.dout(new_net_2209)
	);

	bfr new_net_4844_bfr_after (
		.din(_0444_),
		.dout(new_net_4844)
	);

	bfr new_net_4845_bfr_after (
		.din(new_net_4844),
		.dout(new_net_4845)
	);

	bfr new_net_4846_bfr_after (
		.din(new_net_4845),
		.dout(new_net_4846)
	);

	bfr new_net_4847_bfr_after (
		.din(new_net_4846),
		.dout(new_net_4847)
	);

	bfr new_net_4848_bfr_after (
		.din(new_net_4847),
		.dout(new_net_4848)
	);

	bfr new_net_4849_bfr_after (
		.din(new_net_4848),
		.dout(new_net_4849)
	);

	bfr new_net_4850_bfr_after (
		.din(new_net_4849),
		.dout(new_net_4850)
	);

	bfr new_net_4851_bfr_after (
		.din(new_net_4850),
		.dout(new_net_4851)
	);

	bfr new_net_4852_bfr_after (
		.din(new_net_4851),
		.dout(new_net_4852)
	);

	bfr new_net_4853_bfr_after (
		.din(new_net_4852),
		.dout(new_net_4853)
	);

	bfr new_net_4854_bfr_after (
		.din(new_net_4853),
		.dout(new_net_4854)
	);

	bfr new_net_4855_bfr_after (
		.din(new_net_4854),
		.dout(new_net_4855)
	);

	bfr new_net_4856_bfr_after (
		.din(new_net_4855),
		.dout(new_net_4856)
	);

	bfr new_net_4857_bfr_after (
		.din(new_net_4856),
		.dout(new_net_4857)
	);

	bfr new_net_4858_bfr_after (
		.din(new_net_4857),
		.dout(new_net_4858)
	);

	bfr new_net_4859_bfr_after (
		.din(new_net_4858),
		.dout(new_net_4859)
	);

	bfr new_net_2314_bfr_after (
		.din(new_net_4859),
		.dout(new_net_2314)
	);

	bfr new_net_2230_bfr_after (
		.din(G37),
		.dout(new_net_2230)
	);

	bfr new_net_4860_bfr_after (
		.din(G28),
		.dout(new_net_4860)
	);

	bfr new_net_2251_bfr_after (
		.din(new_net_4860),
		.dout(new_net_2251)
	);

	bfr new_net_4861_bfr_after (
		.din(new_net_2467),
		.dout(new_net_4861)
	);

	bfr new_net_4862_bfr_after (
		.din(new_net_4861),
		.dout(new_net_4862)
	);

	bfr new_net_4863_bfr_after (
		.din(new_net_4862),
		.dout(new_net_4863)
	);

	bfr new_net_4864_bfr_after (
		.din(new_net_4863),
		.dout(new_net_4864)
	);

	bfr new_net_4865_bfr_after (
		.din(new_net_4864),
		.dout(new_net_4865)
	);

	bfr new_net_4866_bfr_after (
		.din(new_net_4865),
		.dout(new_net_4866)
	);

	bfr new_net_4867_bfr_after (
		.din(new_net_4866),
		.dout(new_net_4867)
	);

	bfr new_net_4868_bfr_after (
		.din(new_net_4867),
		.dout(new_net_4868)
	);

	bfr new_net_4869_bfr_after (
		.din(new_net_4868),
		.dout(new_net_4869)
	);

	bfr new_net_4870_bfr_after (
		.din(new_net_4869),
		.dout(new_net_4870)
	);

	bfr new_net_4871_bfr_after (
		.din(new_net_4870),
		.dout(new_net_4871)
	);

	bfr G5272_bfr_after (
		.din(new_net_4871),
		.dout(G5272)
	);

	bfr new_net_4872_bfr_after (
		.din(new_net_2443),
		.dout(new_net_4872)
	);

	bfr new_net_4873_bfr_after (
		.din(new_net_4872),
		.dout(new_net_4873)
	);

	bfr new_net_4874_bfr_after (
		.din(new_net_4873),
		.dout(new_net_4874)
	);

	bfr new_net_4875_bfr_after (
		.din(new_net_4874),
		.dout(new_net_4875)
	);

	bfr new_net_4876_bfr_after (
		.din(new_net_4875),
		.dout(new_net_4876)
	);

	bfr new_net_4877_bfr_after (
		.din(new_net_4876),
		.dout(new_net_4877)
	);

	bfr new_net_4878_bfr_after (
		.din(new_net_4877),
		.dout(new_net_4878)
	);

	bfr new_net_4879_bfr_after (
		.din(new_net_4878),
		.dout(new_net_4879)
	);

	bfr new_net_4880_bfr_after (
		.din(new_net_4879),
		.dout(new_net_4880)
	);

	bfr new_net_4881_bfr_after (
		.din(new_net_4880),
		.dout(new_net_4881)
	);

	bfr new_net_4882_bfr_after (
		.din(new_net_4881),
		.dout(new_net_4882)
	);

	bfr new_net_4883_bfr_after (
		.din(new_net_4882),
		.dout(new_net_4883)
	);

	bfr new_net_4884_bfr_after (
		.din(new_net_4883),
		.dout(new_net_4884)
	);

	bfr new_net_4885_bfr_after (
		.din(new_net_4884),
		.dout(new_net_4885)
	);

	bfr new_net_4886_bfr_after (
		.din(new_net_4885),
		.dout(new_net_4886)
	);

	bfr new_net_4887_bfr_after (
		.din(new_net_4886),
		.dout(new_net_4887)
	);

	bfr new_net_4888_bfr_after (
		.din(new_net_4887),
		.dout(new_net_4888)
	);

	bfr new_net_4889_bfr_after (
		.din(new_net_4888),
		.dout(new_net_4889)
	);

	bfr new_net_4890_bfr_after (
		.din(new_net_4889),
		.dout(new_net_4890)
	);

	bfr new_net_4891_bfr_after (
		.din(new_net_4890),
		.dout(new_net_4891)
	);

	bfr new_net_4892_bfr_after (
		.din(new_net_4891),
		.dout(new_net_4892)
	);

	bfr new_net_4893_bfr_after (
		.din(new_net_4892),
		.dout(new_net_4893)
	);

	bfr new_net_4894_bfr_after (
		.din(new_net_4893),
		.dout(new_net_4894)
	);

	bfr new_net_4895_bfr_after (
		.din(new_net_4894),
		.dout(new_net_4895)
	);

	bfr new_net_4896_bfr_after (
		.din(new_net_4895),
		.dout(new_net_4896)
	);

	bfr new_net_4897_bfr_after (
		.din(new_net_4896),
		.dout(new_net_4897)
	);

	bfr new_net_4898_bfr_after (
		.din(new_net_4897),
		.dout(new_net_4898)
	);

	bfr new_net_4899_bfr_after (
		.din(new_net_4898),
		.dout(new_net_4899)
	);

	bfr new_net_4900_bfr_after (
		.din(new_net_4899),
		.dout(new_net_4900)
	);

	bfr new_net_4901_bfr_after (
		.din(new_net_4900),
		.dout(new_net_4901)
	);

	bfr new_net_4902_bfr_after (
		.din(new_net_4901),
		.dout(new_net_4902)
	);

	bfr new_net_4903_bfr_after (
		.din(new_net_4902),
		.dout(new_net_4903)
	);

	bfr new_net_4904_bfr_after (
		.din(new_net_4903),
		.dout(new_net_4904)
	);

	bfr G5245_bfr_after (
		.din(new_net_4904),
		.dout(G5245)
	);

	bfr new_net_4905_bfr_after (
		.din(new_net_2455),
		.dout(new_net_4905)
	);

	bfr new_net_4906_bfr_after (
		.din(new_net_4905),
		.dout(new_net_4906)
	);

	bfr new_net_4907_bfr_after (
		.din(new_net_4906),
		.dout(new_net_4907)
	);

	bfr new_net_4908_bfr_after (
		.din(new_net_4907),
		.dout(new_net_4908)
	);

	bfr new_net_4909_bfr_after (
		.din(new_net_4908),
		.dout(new_net_4909)
	);

	bfr new_net_4910_bfr_after (
		.din(new_net_4909),
		.dout(new_net_4910)
	);

	bfr G5287_bfr_after (
		.din(new_net_4910),
		.dout(G5287)
	);

	bfr new_net_4911_bfr_after (
		.din(new_net_2479),
		.dout(new_net_4911)
	);

	bfr new_net_4912_bfr_after (
		.din(new_net_4911),
		.dout(new_net_4912)
	);

	bfr new_net_4913_bfr_after (
		.din(new_net_4912),
		.dout(new_net_4913)
	);

	bfr G5299_bfr_after (
		.din(new_net_4913),
		.dout(G5299)
	);

	bfr new_net_4914_bfr_after (
		.din(new_net_2491),
		.dout(new_net_4914)
	);

	bfr new_net_4915_bfr_after (
		.din(new_net_4914),
		.dout(new_net_4915)
	);

	bfr new_net_4916_bfr_after (
		.din(new_net_4915),
		.dout(new_net_4916)
	);

	bfr new_net_4917_bfr_after (
		.din(new_net_4916),
		.dout(new_net_4917)
	);

	bfr new_net_4918_bfr_after (
		.din(new_net_4917),
		.dout(new_net_4918)
	);

	bfr G5306_bfr_after (
		.din(new_net_4918),
		.dout(G5306)
	);

	bfr new_net_4919_bfr_after (
		.din(new_net_2503),
		.dout(new_net_4919)
	);

	bfr new_net_4920_bfr_after (
		.din(new_net_4919),
		.dout(new_net_4920)
	);

	bfr new_net_4921_bfr_after (
		.din(new_net_4920),
		.dout(new_net_4921)
	);

	bfr new_net_4922_bfr_after (
		.din(new_net_4921),
		.dout(new_net_4922)
	);

	bfr new_net_4923_bfr_after (
		.din(new_net_4922),
		.dout(new_net_4923)
	);

	bfr new_net_4924_bfr_after (
		.din(new_net_4923),
		.dout(new_net_4924)
	);

	bfr new_net_4925_bfr_after (
		.din(new_net_4924),
		.dout(new_net_4925)
	);

	bfr new_net_4926_bfr_after (
		.din(new_net_4925),
		.dout(new_net_4926)
	);

	bfr new_net_4927_bfr_after (
		.din(new_net_4926),
		.dout(new_net_4927)
	);

	bfr new_net_4928_bfr_after (
		.din(new_net_4927),
		.dout(new_net_4928)
	);

	bfr new_net_4929_bfr_after (
		.din(new_net_4928),
		.dout(new_net_4929)
	);

	bfr new_net_4930_bfr_after (
		.din(new_net_4929),
		.dout(new_net_4930)
	);

	bfr new_net_4931_bfr_after (
		.din(new_net_4930),
		.dout(new_net_4931)
	);

	bfr new_net_4932_bfr_after (
		.din(new_net_4931),
		.dout(new_net_4932)
	);

	bfr new_net_4933_bfr_after (
		.din(new_net_4932),
		.dout(new_net_4933)
	);

	bfr new_net_4934_bfr_after (
		.din(new_net_4933),
		.dout(new_net_4934)
	);

	bfr new_net_4935_bfr_after (
		.din(new_net_4934),
		.dout(new_net_4935)
	);

	bfr new_net_4936_bfr_after (
		.din(new_net_4935),
		.dout(new_net_4936)
	);

	bfr new_net_4937_bfr_after (
		.din(new_net_4936),
		.dout(new_net_4937)
	);

	bfr new_net_4938_bfr_after (
		.din(new_net_4937),
		.dout(new_net_4938)
	);

	bfr new_net_4939_bfr_after (
		.din(new_net_4938),
		.dout(new_net_4939)
	);

	bfr new_net_4940_bfr_after (
		.din(new_net_4939),
		.dout(new_net_4940)
	);

	bfr new_net_4941_bfr_after (
		.din(new_net_4940),
		.dout(new_net_4941)
	);

	bfr new_net_4942_bfr_after (
		.din(new_net_4941),
		.dout(new_net_4942)
	);

	bfr new_net_4943_bfr_after (
		.din(new_net_4942),
		.dout(new_net_4943)
	);

	bfr new_net_4944_bfr_after (
		.din(new_net_4943),
		.dout(new_net_4944)
	);

	bfr new_net_4945_bfr_after (
		.din(new_net_4944),
		.dout(new_net_4945)
	);

	bfr new_net_4946_bfr_after (
		.din(new_net_4945),
		.dout(new_net_4946)
	);

	bfr new_net_4947_bfr_after (
		.din(new_net_4946),
		.dout(new_net_4947)
	);

	bfr new_net_4948_bfr_after (
		.din(new_net_4947),
		.dout(new_net_4948)
	);

	bfr new_net_4949_bfr_after (
		.din(new_net_4948),
		.dout(new_net_4949)
	);

	bfr new_net_4950_bfr_after (
		.din(new_net_4949),
		.dout(new_net_4950)
	);

	bfr new_net_4951_bfr_after (
		.din(new_net_4950),
		.dout(new_net_4951)
	);

	bfr new_net_4952_bfr_after (
		.din(new_net_4951),
		.dout(new_net_4952)
	);

	bfr G5233_bfr_after (
		.din(new_net_4952),
		.dout(G5233)
	);

	bfr new_net_4953_bfr_after (
		.din(_0732_),
		.dout(new_net_4953)
	);

	bfr new_net_4954_bfr_after (
		.din(new_net_4953),
		.dout(new_net_4954)
	);

	bfr new_net_4955_bfr_after (
		.din(new_net_4954),
		.dout(new_net_4955)
	);

	bfr new_net_4956_bfr_after (
		.din(new_net_4955),
		.dout(new_net_4956)
	);

	bfr new_net_4957_bfr_after (
		.din(new_net_4956),
		.dout(new_net_4957)
	);

	bfr new_net_4958_bfr_after (
		.din(new_net_4957),
		.dout(new_net_4958)
	);

	bfr new_net_4959_bfr_after (
		.din(new_net_4958),
		.dout(new_net_4959)
	);

	bfr new_net_4960_bfr_after (
		.din(new_net_4959),
		.dout(new_net_4960)
	);

	bfr new_net_4961_bfr_after (
		.din(new_net_4960),
		.dout(new_net_4961)
	);

	bfr new_net_4962_bfr_after (
		.din(new_net_4961),
		.dout(new_net_4962)
	);

	bfr new_net_4963_bfr_after (
		.din(new_net_4962),
		.dout(new_net_4963)
	);

	bfr new_net_4964_bfr_after (
		.din(new_net_4963),
		.dout(new_net_4964)
	);

	bfr new_net_4965_bfr_after (
		.din(new_net_4964),
		.dout(new_net_4965)
	);

	bfr new_net_4966_bfr_after (
		.din(new_net_4965),
		.dout(new_net_4966)
	);

	bfr new_net_4967_bfr_after (
		.din(new_net_4966),
		.dout(new_net_4967)
	);

	bfr new_net_4968_bfr_after (
		.din(new_net_4967),
		.dout(new_net_4968)
	);

	bfr new_net_4969_bfr_after (
		.din(new_net_4968),
		.dout(new_net_4969)
	);

	bfr new_net_4970_bfr_after (
		.din(new_net_4969),
		.dout(new_net_4970)
	);

	bfr new_net_2155_bfr_after (
		.din(new_net_4970),
		.dout(new_net_2155)
	);

	bfr new_net_4971_bfr_after (
		.din(_0271_),
		.dout(new_net_4971)
	);

	bfr new_net_4972_bfr_after (
		.din(new_net_4971),
		.dout(new_net_4972)
	);

	bfr new_net_2267_bfr_after (
		.din(new_net_4972),
		.dout(new_net_2267)
	);

	bfr new_net_4973_bfr_after (
		.din(_0512_),
		.dout(new_net_4973)
	);

	bfr new_net_4974_bfr_after (
		.din(new_net_4973),
		.dout(new_net_4974)
	);

	bfr new_net_4975_bfr_after (
		.din(new_net_4974),
		.dout(new_net_4975)
	);

	bfr new_net_4976_bfr_after (
		.din(new_net_4975),
		.dout(new_net_4976)
	);

	bfr new_net_4977_bfr_after (
		.din(new_net_4976),
		.dout(new_net_4977)
	);

	bfr new_net_4978_bfr_after (
		.din(new_net_4977),
		.dout(new_net_4978)
	);

	bfr new_net_4979_bfr_after (
		.din(new_net_4978),
		.dout(new_net_4979)
	);

	bfr new_net_4980_bfr_after (
		.din(new_net_4979),
		.dout(new_net_4980)
	);

	bfr new_net_4981_bfr_after (
		.din(new_net_4980),
		.dout(new_net_4981)
	);

	bfr new_net_4982_bfr_after (
		.din(new_net_4981),
		.dout(new_net_4982)
	);

	bfr new_net_4983_bfr_after (
		.din(new_net_4982),
		.dout(new_net_4983)
	);

	bfr new_net_4984_bfr_after (
		.din(new_net_4983),
		.dout(new_net_4984)
	);

	bfr new_net_4985_bfr_after (
		.din(new_net_4984),
		.dout(new_net_4985)
	);

	bfr new_net_4986_bfr_after (
		.din(new_net_4985),
		.dout(new_net_4986)
	);

	bfr new_net_4987_bfr_after (
		.din(new_net_4986),
		.dout(new_net_4987)
	);

	bfr new_net_4988_bfr_after (
		.din(new_net_4987),
		.dout(new_net_4988)
	);

	bfr new_net_4989_bfr_after (
		.din(new_net_4988),
		.dout(new_net_4989)
	);

	bfr new_net_4990_bfr_after (
		.din(new_net_4989),
		.dout(new_net_4990)
	);

	bfr new_net_4991_bfr_after (
		.din(new_net_4990),
		.dout(new_net_4991)
	);

	bfr new_net_4992_bfr_after (
		.din(new_net_4991),
		.dout(new_net_4992)
	);

	bfr new_net_4993_bfr_after (
		.din(new_net_4992),
		.dout(new_net_4993)
	);

	bfr new_net_4994_bfr_after (
		.din(new_net_4993),
		.dout(new_net_4994)
	);

	bfr new_net_4995_bfr_after (
		.din(new_net_4994),
		.dout(new_net_4995)
	);

	bfr new_net_4996_bfr_after (
		.din(new_net_4995),
		.dout(new_net_4996)
	);

	bfr new_net_4997_bfr_after (
		.din(new_net_4996),
		.dout(new_net_4997)
	);

	bfr new_net_4998_bfr_after (
		.din(new_net_4997),
		.dout(new_net_4998)
	);

	bfr new_net_4999_bfr_after (
		.din(new_net_4998),
		.dout(new_net_4999)
	);

	bfr new_net_5000_bfr_after (
		.din(new_net_4999),
		.dout(new_net_5000)
	);

	bfr new_net_5001_bfr_after (
		.din(new_net_5000),
		.dout(new_net_5001)
	);

	bfr new_net_5002_bfr_after (
		.din(new_net_5001),
		.dout(new_net_5002)
	);

	bfr new_net_5003_bfr_after (
		.din(new_net_5002),
		.dout(new_net_5003)
	);

	bfr new_net_2330_bfr_after (
		.din(new_net_5003),
		.dout(new_net_2330)
	);

	bfr new_net_5004_bfr_after (
		.din(new_net_2449),
		.dout(new_net_5004)
	);

	bfr new_net_5005_bfr_after (
		.din(new_net_5004),
		.dout(new_net_5005)
	);

	bfr G5305_bfr_after (
		.din(new_net_5005),
		.dout(G5305)
	);

	bfr new_net_5006_bfr_after (
		.din(new_net_2473),
		.dout(new_net_5006)
	);

	bfr new_net_5007_bfr_after (
		.din(new_net_5006),
		.dout(new_net_5007)
	);

	bfr new_net_5008_bfr_after (
		.din(new_net_5007),
		.dout(new_net_5008)
	);

	bfr new_net_5009_bfr_after (
		.din(new_net_5008),
		.dout(new_net_5009)
	);

	bfr new_net_5010_bfr_after (
		.din(new_net_5009),
		.dout(new_net_5010)
	);

	bfr new_net_5011_bfr_after (
		.din(new_net_5010),
		.dout(new_net_5011)
	);

	bfr new_net_5012_bfr_after (
		.din(new_net_5011),
		.dout(new_net_5012)
	);

	bfr new_net_5013_bfr_after (
		.din(new_net_5012),
		.dout(new_net_5013)
	);

	bfr new_net_5014_bfr_after (
		.din(new_net_5013),
		.dout(new_net_5014)
	);

	bfr new_net_5015_bfr_after (
		.din(new_net_5014),
		.dout(new_net_5015)
	);

	bfr G5271_bfr_after (
		.din(new_net_5015),
		.dout(G5271)
	);

	bfr new_net_5016_bfr_after (
		.din(G116),
		.dout(new_net_5016)
	);

	bfr new_net_5017_bfr_after (
		.din(new_net_5016),
		.dout(new_net_5017)
	);

	bfr new_net_2107_bfr_after (
		.din(new_net_5017),
		.dout(new_net_2107)
	);

	bfr new_net_5018_bfr_after (
		.din(_0606_),
		.dout(new_net_5018)
	);

	bfr new_net_5019_bfr_after (
		.din(new_net_5018),
		.dout(new_net_5019)
	);

	bfr new_net_5020_bfr_after (
		.din(new_net_5019),
		.dout(new_net_5020)
	);

	bfr new_net_2120_bfr_after (
		.din(new_net_5020),
		.dout(new_net_2120)
	);

	bfr new_net_5021_bfr_after (
		.din(G50),
		.dout(new_net_5021)
	);

	bfr new_net_5022_bfr_after (
		.din(new_net_5021),
		.dout(new_net_5022)
	);

	bfr new_net_5023_bfr_after (
		.din(new_net_5022),
		.dout(new_net_5023)
	);

	bfr new_net_5024_bfr_after (
		.din(new_net_5023),
		.dout(new_net_5024)
	);

	bfr new_net_2141_bfr_after (
		.din(new_net_5024),
		.dout(new_net_2141)
	);

	bfr new_net_5025_bfr_after (
		.din(_0832_),
		.dout(new_net_5025)
	);

	bfr new_net_5026_bfr_after (
		.din(new_net_5025),
		.dout(new_net_5026)
	);

	bfr new_net_5027_bfr_after (
		.din(new_net_5026),
		.dout(new_net_5027)
	);

	bfr new_net_5028_bfr_after (
		.din(new_net_5027),
		.dout(new_net_5028)
	);

	bfr new_net_5029_bfr_after (
		.din(new_net_5028),
		.dout(new_net_5029)
	);

	bfr new_net_5030_bfr_after (
		.din(new_net_5029),
		.dout(new_net_5030)
	);

	bfr new_net_5031_bfr_after (
		.din(new_net_5030),
		.dout(new_net_5031)
	);

	bfr new_net_5032_bfr_after (
		.din(new_net_5031),
		.dout(new_net_5032)
	);

	bfr new_net_5033_bfr_after (
		.din(new_net_5032),
		.dout(new_net_5033)
	);

	bfr new_net_5034_bfr_after (
		.din(new_net_5033),
		.dout(new_net_5034)
	);

	bfr new_net_5035_bfr_after (
		.din(new_net_5034),
		.dout(new_net_5035)
	);

	bfr new_net_5036_bfr_after (
		.din(new_net_5035),
		.dout(new_net_5036)
	);

	bfr new_net_2162_bfr_after (
		.din(new_net_5036),
		.dout(new_net_2162)
	);

	bfr new_net_5037_bfr_after (
		.din(G89),
		.dout(new_net_5037)
	);

	bfr new_net_2183_bfr_after (
		.din(new_net_5037),
		.dout(new_net_2183)
	);

	bfr new_net_2288_bfr_after (
		.din(_0338_),
		.dout(new_net_2288)
	);

	bfr new_net_5038_bfr_after (
		.din(new_net_2427),
		.dout(new_net_5038)
	);

	bfr new_net_5039_bfr_after (
		.din(new_net_5038),
		.dout(new_net_5039)
	);

	bfr new_net_5040_bfr_after (
		.din(new_net_5039),
		.dout(new_net_5040)
	);

	bfr new_net_5041_bfr_after (
		.din(new_net_5040),
		.dout(new_net_5041)
	);

	bfr new_net_5042_bfr_after (
		.din(new_net_5041),
		.dout(new_net_5042)
	);

	bfr new_net_5043_bfr_after (
		.din(new_net_5042),
		.dout(new_net_5043)
	);

	bfr new_net_5044_bfr_after (
		.din(new_net_5043),
		.dout(new_net_5044)
	);

	bfr new_net_5045_bfr_after (
		.din(new_net_5044),
		.dout(new_net_5045)
	);

	bfr new_net_5046_bfr_after (
		.din(new_net_5045),
		.dout(new_net_5046)
	);

	bfr new_net_5047_bfr_after (
		.din(new_net_5046),
		.dout(new_net_5047)
	);

	bfr new_net_5048_bfr_after (
		.din(new_net_5047),
		.dout(new_net_5048)
	);

	bfr new_net_5049_bfr_after (
		.din(new_net_5048),
		.dout(new_net_5049)
	);

	bfr new_net_5050_bfr_after (
		.din(new_net_5049),
		.dout(new_net_5050)
	);

	bfr new_net_5051_bfr_after (
		.din(new_net_5050),
		.dout(new_net_5051)
	);

	bfr new_net_5052_bfr_after (
		.din(new_net_5051),
		.dout(new_net_5052)
	);

	bfr new_net_5053_bfr_after (
		.din(new_net_5052),
		.dout(new_net_5053)
	);

	bfr new_net_5054_bfr_after (
		.din(new_net_5053),
		.dout(new_net_5054)
	);

	bfr new_net_5055_bfr_after (
		.din(new_net_5054),
		.dout(new_net_5055)
	);

	bfr G5265_bfr_after (
		.din(new_net_5055),
		.dout(G5265)
	);

	bfr new_net_2241_bfr_after (
		.din(G63),
		.dout(new_net_2241)
	);

	bfr new_net_5056_bfr_after (
		.din(_0490_),
		.dout(new_net_5056)
	);

	bfr new_net_5057_bfr_after (
		.din(new_net_5056),
		.dout(new_net_5057)
	);

	bfr new_net_5058_bfr_after (
		.din(new_net_5057),
		.dout(new_net_5058)
	);

	bfr new_net_5059_bfr_after (
		.din(new_net_5058),
		.dout(new_net_5059)
	);

	bfr new_net_5060_bfr_after (
		.din(new_net_5059),
		.dout(new_net_5060)
	);

	bfr new_net_5061_bfr_after (
		.din(new_net_5060),
		.dout(new_net_5061)
	);

	bfr new_net_5062_bfr_after (
		.din(new_net_5061),
		.dout(new_net_5062)
	);

	bfr new_net_5063_bfr_after (
		.din(new_net_5062),
		.dout(new_net_5063)
	);

	bfr new_net_5064_bfr_after (
		.din(new_net_5063),
		.dout(new_net_5064)
	);

	bfr new_net_5065_bfr_after (
		.din(new_net_5064),
		.dout(new_net_5065)
	);

	bfr new_net_5066_bfr_after (
		.din(new_net_5065),
		.dout(new_net_5066)
	);

	bfr new_net_5067_bfr_after (
		.din(new_net_5066),
		.dout(new_net_5067)
	);

	bfr new_net_5068_bfr_after (
		.din(new_net_5067),
		.dout(new_net_5068)
	);

	bfr new_net_5069_bfr_after (
		.din(new_net_5068),
		.dout(new_net_5069)
	);

	bfr new_net_5070_bfr_after (
		.din(new_net_5069),
		.dout(new_net_5070)
	);

	bfr new_net_5071_bfr_after (
		.din(new_net_5070),
		.dout(new_net_5071)
	);

	bfr new_net_5072_bfr_after (
		.din(new_net_5071),
		.dout(new_net_5072)
	);

	bfr new_net_5073_bfr_after (
		.din(new_net_5072),
		.dout(new_net_5073)
	);

	bfr new_net_5074_bfr_after (
		.din(new_net_5073),
		.dout(new_net_5074)
	);

	bfr new_net_5075_bfr_after (
		.din(new_net_5074),
		.dout(new_net_5075)
	);

	bfr new_net_5076_bfr_after (
		.din(new_net_5075),
		.dout(new_net_5076)
	);

	bfr new_net_5077_bfr_after (
		.din(new_net_5076),
		.dout(new_net_5077)
	);

	bfr new_net_5078_bfr_after (
		.din(new_net_5077),
		.dout(new_net_5078)
	);

	bfr new_net_5079_bfr_after (
		.din(new_net_5078),
		.dout(new_net_5079)
	);

	bfr new_net_5080_bfr_after (
		.din(new_net_5079),
		.dout(new_net_5080)
	);

	bfr new_net_5081_bfr_after (
		.din(new_net_5080),
		.dout(new_net_5081)
	);

	bfr new_net_5082_bfr_after (
		.din(new_net_5081),
		.dout(new_net_5082)
	);

	bfr new_net_5083_bfr_after (
		.din(new_net_5082),
		.dout(new_net_5083)
	);

	bfr new_net_5084_bfr_after (
		.din(new_net_5083),
		.dout(new_net_5084)
	);

	bfr new_net_5085_bfr_after (
		.din(new_net_5084),
		.dout(new_net_5085)
	);

	bfr new_net_2325_bfr_after (
		.din(new_net_5085),
		.dout(new_net_2325)
	);

	bfr new_net_2262_bfr_after (
		.din(_0245_),
		.dout(new_net_2262)
	);

	bfr new_net_5086_bfr_after (
		.din(_0700_),
		.dout(new_net_5086)
	);

	bfr new_net_5087_bfr_after (
		.din(new_net_5086),
		.dout(new_net_5087)
	);

	bfr new_net_5088_bfr_after (
		.din(new_net_5087),
		.dout(new_net_5088)
	);

	bfr new_net_5089_bfr_after (
		.din(new_net_5088),
		.dout(new_net_5089)
	);

	bfr new_net_5090_bfr_after (
		.din(new_net_5089),
		.dout(new_net_5090)
	);

	bfr new_net_5091_bfr_after (
		.din(new_net_5090),
		.dout(new_net_5091)
	);

	bfr new_net_5092_bfr_after (
		.din(new_net_5091),
		.dout(new_net_5092)
	);

	bfr new_net_5093_bfr_after (
		.din(new_net_5092),
		.dout(new_net_5093)
	);

	bfr new_net_5094_bfr_after (
		.din(new_net_5093),
		.dout(new_net_5094)
	);

	bfr new_net_5095_bfr_after (
		.din(new_net_5094),
		.dout(new_net_5095)
	);

	bfr new_net_5096_bfr_after (
		.din(new_net_5095),
		.dout(new_net_5096)
	);

	bfr new_net_5097_bfr_after (
		.din(new_net_5096),
		.dout(new_net_5097)
	);

	bfr new_net_2136_bfr_after (
		.din(new_net_5097),
		.dout(new_net_2136)
	);

	bfr new_net_5098_bfr_after (
		.din(_0794_),
		.dout(new_net_5098)
	);

	bfr new_net_2157_bfr_after (
		.din(new_net_5098),
		.dout(new_net_2157)
	);

	bfr new_net_5099_bfr_after (
		.din(_0889_),
		.dout(new_net_5099)
	);

	bfr new_net_5100_bfr_after (
		.din(new_net_5099),
		.dout(new_net_5100)
	);

	bfr new_net_5101_bfr_after (
		.din(new_net_5100),
		.dout(new_net_5101)
	);

	bfr new_net_5102_bfr_after (
		.din(new_net_5101),
		.dout(new_net_5102)
	);

	bfr new_net_5103_bfr_after (
		.din(new_net_5102),
		.dout(new_net_5103)
	);

	bfr new_net_5104_bfr_after (
		.din(new_net_5103),
		.dout(new_net_5104)
	);

	bfr new_net_5105_bfr_after (
		.din(new_net_5104),
		.dout(new_net_5105)
	);

	bfr new_net_5106_bfr_after (
		.din(new_net_5105),
		.dout(new_net_5106)
	);

	bfr new_net_5107_bfr_after (
		.din(new_net_5106),
		.dout(new_net_5107)
	);

	bfr new_net_5108_bfr_after (
		.din(new_net_5107),
		.dout(new_net_5108)
	);

	bfr new_net_5109_bfr_after (
		.din(new_net_5108),
		.dout(new_net_5109)
	);

	bfr new_net_5110_bfr_after (
		.din(new_net_5109),
		.dout(new_net_5110)
	);

	bfr new_net_5111_bfr_after (
		.din(new_net_5110),
		.dout(new_net_5111)
	);

	bfr new_net_5112_bfr_after (
		.din(new_net_5111),
		.dout(new_net_5112)
	);

	bfr new_net_5113_bfr_after (
		.din(new_net_5112),
		.dout(new_net_5113)
	);

	bfr new_net_5114_bfr_after (
		.din(new_net_5113),
		.dout(new_net_5114)
	);

	bfr new_net_5115_bfr_after (
		.din(new_net_5114),
		.dout(new_net_5115)
	);

	bfr new_net_5116_bfr_after (
		.din(new_net_5115),
		.dout(new_net_5116)
	);

	bfr new_net_5117_bfr_after (
		.din(new_net_5116),
		.dout(new_net_5117)
	);

	bfr new_net_5118_bfr_after (
		.din(new_net_5117),
		.dout(new_net_5118)
	);

	bfr new_net_5119_bfr_after (
		.din(new_net_5118),
		.dout(new_net_5119)
	);

	bfr new_net_5120_bfr_after (
		.din(new_net_5119),
		.dout(new_net_5120)
	);

	bfr new_net_5121_bfr_after (
		.din(new_net_5120),
		.dout(new_net_5121)
	);

	bfr new_net_5122_bfr_after (
		.din(new_net_5121),
		.dout(new_net_5122)
	);

	bfr new_net_2178_bfr_after (
		.din(new_net_5122),
		.dout(new_net_2178)
	);

	bfr new_net_5123_bfr_after (
		.din(G13),
		.dout(new_net_5123)
	);

	bfr new_net_2115_bfr_after (
		.din(new_net_5123),
		.dout(new_net_2115)
	);

	bfr new_net_5124_bfr_after (
		.din(G44),
		.dout(new_net_5124)
	);

	bfr new_net_5125_bfr_after (
		.din(new_net_5124),
		.dout(new_net_5125)
	);

	bfr new_net_5126_bfr_after (
		.din(new_net_5125),
		.dout(new_net_5126)
	);

	bfr new_net_5127_bfr_after (
		.din(new_net_5126),
		.dout(new_net_5127)
	);

	bfr new_net_2199_bfr_after (
		.din(new_net_5127),
		.dout(new_net_2199)
	);

	bfr new_net_5128_bfr_after (
		.din(_0317_),
		.dout(new_net_5128)
	);

	bfr new_net_5129_bfr_after (
		.din(new_net_5128),
		.dout(new_net_5129)
	);

	bfr new_net_2283_bfr_after (
		.din(new_net_5129),
		.dout(new_net_2283)
	);

	bfr new_net_5130_bfr_after (
		.din(_0570_),
		.dout(new_net_5130)
	);

	bfr new_net_5131_bfr_after (
		.din(new_net_5130),
		.dout(new_net_5131)
	);

	bfr new_net_5132_bfr_after (
		.din(new_net_5131),
		.dout(new_net_5132)
	);

	bfr new_net_5133_bfr_after (
		.din(new_net_5132),
		.dout(new_net_5133)
	);

	bfr new_net_5134_bfr_after (
		.din(new_net_5133),
		.dout(new_net_5134)
	);

	bfr new_net_5135_bfr_after (
		.din(new_net_5134),
		.dout(new_net_5135)
	);

	bfr new_net_5136_bfr_after (
		.din(new_net_5135),
		.dout(new_net_5136)
	);

	bfr new_net_5137_bfr_after (
		.din(new_net_5136),
		.dout(new_net_5137)
	);

	bfr new_net_5138_bfr_after (
		.din(new_net_5137),
		.dout(new_net_5138)
	);

	bfr new_net_5139_bfr_after (
		.din(new_net_5138),
		.dout(new_net_5139)
	);

	bfr new_net_5140_bfr_after (
		.din(new_net_5139),
		.dout(new_net_5140)
	);

	bfr new_net_5141_bfr_after (
		.din(new_net_5140),
		.dout(new_net_5141)
	);

	bfr new_net_5142_bfr_after (
		.din(new_net_5141),
		.dout(new_net_5142)
	);

	bfr new_net_5143_bfr_after (
		.din(new_net_5142),
		.dout(new_net_5143)
	);

	bfr new_net_5144_bfr_after (
		.din(new_net_5143),
		.dout(new_net_5144)
	);

	bfr new_net_5145_bfr_after (
		.din(new_net_5144),
		.dout(new_net_5145)
	);

	bfr new_net_5146_bfr_after (
		.din(new_net_5145),
		.dout(new_net_5146)
	);

	bfr new_net_5147_bfr_after (
		.din(new_net_5146),
		.dout(new_net_5147)
	);

	bfr new_net_5148_bfr_after (
		.din(new_net_5147),
		.dout(new_net_5148)
	);

	bfr new_net_5149_bfr_after (
		.din(new_net_5148),
		.dout(new_net_5149)
	);

	bfr new_net_5150_bfr_after (
		.din(new_net_5149),
		.dout(new_net_5150)
	);

	bfr new_net_5151_bfr_after (
		.din(new_net_5150),
		.dout(new_net_5151)
	);

	bfr new_net_5152_bfr_after (
		.din(new_net_5151),
		.dout(new_net_5152)
	);

	bfr new_net_5153_bfr_after (
		.din(new_net_5152),
		.dout(new_net_5153)
	);

	bfr new_net_5154_bfr_after (
		.din(new_net_5153),
		.dout(new_net_5154)
	);

	bfr new_net_5155_bfr_after (
		.din(new_net_5154),
		.dout(new_net_5155)
	);

	bfr new_net_5156_bfr_after (
		.din(new_net_5155),
		.dout(new_net_5156)
	);

	bfr new_net_5157_bfr_after (
		.din(new_net_5156),
		.dout(new_net_5157)
	);

	bfr new_net_5158_bfr_after (
		.din(new_net_5157),
		.dout(new_net_5158)
	);

	bfr new_net_5159_bfr_after (
		.din(new_net_5158),
		.dout(new_net_5159)
	);

	bfr new_net_5160_bfr_after (
		.din(new_net_5159),
		.dout(new_net_5160)
	);

	bfr new_net_5161_bfr_after (
		.din(new_net_5160),
		.dout(new_net_5161)
	);

	bfr new_net_2346_bfr_after (
		.din(new_net_5161),
		.dout(new_net_2346)
	);

	bfr new_net_5162_bfr_after (
		.din(new_net_2437),
		.dout(new_net_5162)
	);

	bfr new_net_5163_bfr_after (
		.din(new_net_5162),
		.dout(new_net_5163)
	);

	bfr new_net_5164_bfr_after (
		.din(new_net_5163),
		.dout(new_net_5164)
	);

	bfr new_net_5165_bfr_after (
		.din(new_net_5164),
		.dout(new_net_5165)
	);

	bfr new_net_5166_bfr_after (
		.din(new_net_5165),
		.dout(new_net_5166)
	);

	bfr new_net_5167_bfr_after (
		.din(new_net_5166),
		.dout(new_net_5167)
	);

	bfr new_net_5168_bfr_after (
		.din(new_net_5167),
		.dout(new_net_5168)
	);

	bfr new_net_5169_bfr_after (
		.din(new_net_5168),
		.dout(new_net_5169)
	);

	bfr new_net_5170_bfr_after (
		.din(new_net_5169),
		.dout(new_net_5170)
	);

	bfr new_net_5171_bfr_after (
		.din(new_net_5170),
		.dout(new_net_5171)
	);

	bfr G5267_bfr_after (
		.din(new_net_5171),
		.dout(G5267)
	);

	bfr G5315_bfr_after (
		.din(new_net_2357),
		.dout(G5315)
	);

	bfr new_net_5172_bfr_after (
		.din(new_net_2369),
		.dout(new_net_5172)
	);

	bfr new_net_5173_bfr_after (
		.din(new_net_5172),
		.dout(new_net_5173)
	);

	bfr new_net_5174_bfr_after (
		.din(new_net_5173),
		.dout(new_net_5174)
	);

	bfr new_net_5175_bfr_after (
		.din(new_net_5174),
		.dout(new_net_5175)
	);

	bfr new_net_5176_bfr_after (
		.din(new_net_5175),
		.dout(new_net_5176)
	);

	bfr new_net_5177_bfr_after (
		.din(new_net_5176),
		.dout(new_net_5177)
	);

	bfr new_net_5178_bfr_after (
		.din(new_net_5177),
		.dout(new_net_5178)
	);

	bfr new_net_5179_bfr_after (
		.din(new_net_5178),
		.dout(new_net_5179)
	);

	bfr new_net_5180_bfr_after (
		.din(new_net_5179),
		.dout(new_net_5180)
	);

	bfr new_net_5181_bfr_after (
		.din(new_net_5180),
		.dout(new_net_5181)
	);

	bfr new_net_5182_bfr_after (
		.din(new_net_5181),
		.dout(new_net_5182)
	);

	bfr new_net_5183_bfr_after (
		.din(new_net_5182),
		.dout(new_net_5183)
	);

	bfr new_net_5184_bfr_after (
		.din(new_net_5183),
		.dout(new_net_5184)
	);

	bfr new_net_5185_bfr_after (
		.din(new_net_5184),
		.dout(new_net_5185)
	);

	bfr new_net_5186_bfr_after (
		.din(new_net_5185),
		.dout(new_net_5186)
	);

	bfr G5270_bfr_after (
		.din(new_net_5186),
		.dout(G5270)
	);

	bfr new_net_5187_bfr_after (
		.din(new_net_2381),
		.dout(new_net_5187)
	);

	bfr G5303_bfr_after (
		.din(new_net_5187),
		.dout(G5303)
	);

	bfr new_net_5188_bfr_after (
		.din(new_net_2393),
		.dout(new_net_5188)
	);

	bfr new_net_5189_bfr_after (
		.din(new_net_5188),
		.dout(new_net_5189)
	);

	bfr new_net_5190_bfr_after (
		.din(new_net_5189),
		.dout(new_net_5190)
	);

	bfr new_net_5191_bfr_after (
		.din(new_net_5190),
		.dout(new_net_5191)
	);

	bfr new_net_5192_bfr_after (
		.din(new_net_5191),
		.dout(new_net_5192)
	);

	bfr new_net_5193_bfr_after (
		.din(new_net_5192),
		.dout(new_net_5193)
	);

	bfr new_net_5194_bfr_after (
		.din(new_net_5193),
		.dout(new_net_5194)
	);

	bfr new_net_5195_bfr_after (
		.din(new_net_5194),
		.dout(new_net_5195)
	);

	bfr new_net_5196_bfr_after (
		.din(new_net_5195),
		.dout(new_net_5196)
	);

	bfr new_net_5197_bfr_after (
		.din(new_net_5196),
		.dout(new_net_5197)
	);

	bfr new_net_5198_bfr_after (
		.din(new_net_5197),
		.dout(new_net_5198)
	);

	bfr new_net_5199_bfr_after (
		.din(new_net_5198),
		.dout(new_net_5199)
	);

	bfr new_net_5200_bfr_after (
		.din(new_net_5199),
		.dout(new_net_5200)
	);

	bfr new_net_5201_bfr_after (
		.din(new_net_5200),
		.dout(new_net_5201)
	);

	bfr new_net_5202_bfr_after (
		.din(new_net_5201),
		.dout(new_net_5202)
	);

	bfr new_net_5203_bfr_after (
		.din(new_net_5202),
		.dout(new_net_5203)
	);

	bfr new_net_5204_bfr_after (
		.din(new_net_5203),
		.dout(new_net_5204)
	);

	bfr new_net_5205_bfr_after (
		.din(new_net_5204),
		.dout(new_net_5205)
	);

	bfr new_net_5206_bfr_after (
		.din(new_net_5205),
		.dout(new_net_5206)
	);

	bfr new_net_5207_bfr_after (
		.din(new_net_5206),
		.dout(new_net_5207)
	);

	bfr new_net_5208_bfr_after (
		.din(new_net_5207),
		.dout(new_net_5208)
	);

	bfr new_net_5209_bfr_after (
		.din(new_net_5208),
		.dout(new_net_5209)
	);

	bfr new_net_5210_bfr_after (
		.din(new_net_5209),
		.dout(new_net_5210)
	);

	bfr new_net_5211_bfr_after (
		.din(new_net_5210),
		.dout(new_net_5211)
	);

	bfr new_net_5212_bfr_after (
		.din(new_net_5211),
		.dout(new_net_5212)
	);

	bfr new_net_5213_bfr_after (
		.din(new_net_5212),
		.dout(new_net_5213)
	);

	bfr new_net_5214_bfr_after (
		.din(new_net_5213),
		.dout(new_net_5214)
	);

	bfr new_net_5215_bfr_after (
		.din(new_net_5214),
		.dout(new_net_5215)
	);

	bfr new_net_5216_bfr_after (
		.din(new_net_5215),
		.dout(new_net_5216)
	);

	bfr new_net_5217_bfr_after (
		.din(new_net_5216),
		.dout(new_net_5217)
	);

	bfr new_net_5218_bfr_after (
		.din(new_net_5217),
		.dout(new_net_5218)
	);

	bfr new_net_5219_bfr_after (
		.din(new_net_5218),
		.dout(new_net_5219)
	);

	bfr new_net_5220_bfr_after (
		.din(new_net_5219),
		.dout(new_net_5220)
	);

	bfr new_net_5221_bfr_after (
		.din(new_net_5220),
		.dout(new_net_5221)
	);

	bfr new_net_5222_bfr_after (
		.din(new_net_5221),
		.dout(new_net_5222)
	);

	bfr new_net_5223_bfr_after (
		.din(new_net_5222),
		.dout(new_net_5223)
	);

	bfr new_net_5224_bfr_after (
		.din(new_net_5223),
		.dout(new_net_5224)
	);

	bfr new_net_5225_bfr_after (
		.din(new_net_5224),
		.dout(new_net_5225)
	);

	bfr new_net_5226_bfr_after (
		.din(new_net_5225),
		.dout(new_net_5226)
	);

	bfr G5211_bfr_after (
		.din(new_net_5226),
		.dout(G5211)
	);

	bfr new_net_5227_bfr_after (
		.din(new_net_2405),
		.dout(new_net_5227)
	);

	bfr new_net_5228_bfr_after (
		.din(new_net_5227),
		.dout(new_net_5228)
	);

	bfr new_net_5229_bfr_after (
		.din(new_net_5228),
		.dout(new_net_5229)
	);

	bfr G5300_bfr_after (
		.din(new_net_5229),
		.dout(G5300)
	);

	bfr new_net_5230_bfr_after (
		.din(_0926_),
		.dout(new_net_5230)
	);

	bfr new_net_5231_bfr_after (
		.din(new_net_5230),
		.dout(new_net_5231)
	);

	bfr new_net_5232_bfr_after (
		.din(new_net_5231),
		.dout(new_net_5232)
	);

	bfr new_net_5233_bfr_after (
		.din(new_net_5232),
		.dout(new_net_5233)
	);

	bfr new_net_5234_bfr_after (
		.din(new_net_5233),
		.dout(new_net_5234)
	);

	bfr new_net_5235_bfr_after (
		.din(new_net_5234),
		.dout(new_net_5235)
	);

	bfr new_net_5236_bfr_after (
		.din(new_net_5235),
		.dout(new_net_5236)
	);

	bfr new_net_5237_bfr_after (
		.din(new_net_5236),
		.dout(new_net_5237)
	);

	bfr new_net_5238_bfr_after (
		.din(new_net_5237),
		.dout(new_net_5238)
	);

	bfr new_net_5239_bfr_after (
		.din(new_net_5238),
		.dout(new_net_5239)
	);

	bfr new_net_5240_bfr_after (
		.din(new_net_5239),
		.dout(new_net_5240)
	);

	bfr new_net_5241_bfr_after (
		.din(new_net_5240),
		.dout(new_net_5241)
	);

	bfr new_net_5242_bfr_after (
		.din(new_net_5241),
		.dout(new_net_5242)
	);

	bfr new_net_5243_bfr_after (
		.din(new_net_5242),
		.dout(new_net_5243)
	);

	bfr new_net_5244_bfr_after (
		.din(new_net_5243),
		.dout(new_net_5244)
	);

	bfr new_net_5245_bfr_after (
		.din(new_net_5244),
		.dout(new_net_5245)
	);

	bfr new_net_2180_bfr_after (
		.din(new_net_5245),
		.dout(new_net_2180)
	);

	bfr new_net_2117_bfr_after (
		.din(_0591_),
		.dout(new_net_2117)
	);

	bfr new_net_5246_bfr_after (
		.din(new_net_2403),
		.dout(new_net_5246)
	);

	bfr new_net_5247_bfr_after (
		.din(new_net_5246),
		.dout(new_net_5247)
	);

	bfr new_net_5248_bfr_after (
		.din(new_net_5247),
		.dout(new_net_5248)
	);

	bfr new_net_5249_bfr_after (
		.din(new_net_5248),
		.dout(new_net_5249)
	);

	bfr new_net_5250_bfr_after (
		.din(new_net_5249),
		.dout(new_net_5250)
	);

	bfr new_net_5251_bfr_after (
		.din(new_net_5250),
		.dout(new_net_5251)
	);

	bfr new_net_5252_bfr_after (
		.din(new_net_5251),
		.dout(new_net_5252)
	);

	bfr new_net_5253_bfr_after (
		.din(new_net_5252),
		.dout(new_net_5253)
	);

	bfr new_net_5254_bfr_after (
		.din(new_net_5253),
		.dout(new_net_5254)
	);

	bfr new_net_5255_bfr_after (
		.din(new_net_5254),
		.dout(new_net_5255)
	);

	bfr new_net_5256_bfr_after (
		.din(new_net_5255),
		.dout(new_net_5256)
	);

	bfr new_net_5257_bfr_after (
		.din(new_net_5256),
		.dout(new_net_5257)
	);

	bfr new_net_5258_bfr_after (
		.din(new_net_5257),
		.dout(new_net_5258)
	);

	bfr new_net_5259_bfr_after (
		.din(new_net_5258),
		.dout(new_net_5259)
	);

	bfr new_net_5260_bfr_after (
		.din(new_net_5259),
		.dout(new_net_5260)
	);

	bfr new_net_5261_bfr_after (
		.din(new_net_5260),
		.dout(new_net_5261)
	);

	bfr new_net_5262_bfr_after (
		.din(new_net_5261),
		.dout(new_net_5262)
	);

	bfr new_net_5263_bfr_after (
		.din(new_net_5262),
		.dout(new_net_5263)
	);

	bfr new_net_5264_bfr_after (
		.din(new_net_5263),
		.dout(new_net_5264)
	);

	bfr new_net_5265_bfr_after (
		.din(new_net_5264),
		.dout(new_net_5265)
	);

	bfr new_net_5266_bfr_after (
		.din(new_net_5265),
		.dout(new_net_5266)
	);

	bfr new_net_5267_bfr_after (
		.din(new_net_5266),
		.dout(new_net_5267)
	);

	bfr new_net_5268_bfr_after (
		.din(new_net_5267),
		.dout(new_net_5268)
	);

	bfr new_net_5269_bfr_after (
		.din(new_net_5268),
		.dout(new_net_5269)
	);

	bfr new_net_5270_bfr_after (
		.din(new_net_5269),
		.dout(new_net_5270)
	);

	bfr new_net_5271_bfr_after (
		.din(new_net_5270),
		.dout(new_net_5271)
	);

	bfr new_net_5272_bfr_after (
		.din(new_net_5271),
		.dout(new_net_5272)
	);

	bfr new_net_5273_bfr_after (
		.din(new_net_5272),
		.dout(new_net_5273)
	);

	bfr new_net_5274_bfr_after (
		.din(new_net_5273),
		.dout(new_net_5274)
	);

	bfr new_net_5275_bfr_after (
		.din(new_net_5274),
		.dout(new_net_5275)
	);

	bfr new_net_5276_bfr_after (
		.din(new_net_5275),
		.dout(new_net_5276)
	);

	bfr new_net_5277_bfr_after (
		.din(new_net_5276),
		.dout(new_net_5277)
	);

	bfr new_net_5278_bfr_after (
		.din(new_net_5277),
		.dout(new_net_5278)
	);

	bfr new_net_5279_bfr_after (
		.din(new_net_5278),
		.dout(new_net_5279)
	);

	bfr new_net_5280_bfr_after (
		.din(new_net_5279),
		.dout(new_net_5280)
	);

	bfr new_net_5281_bfr_after (
		.din(new_net_5280),
		.dout(new_net_5281)
	);

	bfr new_net_5282_bfr_after (
		.din(new_net_5281),
		.dout(new_net_5282)
	);

	bfr new_net_5283_bfr_after (
		.din(new_net_5282),
		.dout(new_net_5283)
	);

	bfr new_net_5284_bfr_after (
		.din(new_net_5283),
		.dout(new_net_5284)
	);

	bfr G5207_bfr_after (
		.din(new_net_5284),
		.dout(G5207)
	);

	bfr new_net_5285_bfr_after (
		.din(_0870_),
		.dout(new_net_5285)
	);

	bfr new_net_5286_bfr_after (
		.din(new_net_5285),
		.dout(new_net_5286)
	);

	bfr new_net_5287_bfr_after (
		.din(new_net_5286),
		.dout(new_net_5287)
	);

	bfr new_net_5288_bfr_after (
		.din(new_net_5287),
		.dout(new_net_5288)
	);

	bfr new_net_5289_bfr_after (
		.din(new_net_5288),
		.dout(new_net_5289)
	);

	bfr new_net_5290_bfr_after (
		.din(new_net_5289),
		.dout(new_net_5290)
	);

	bfr new_net_5291_bfr_after (
		.din(new_net_5290),
		.dout(new_net_5291)
	);

	bfr new_net_5292_bfr_after (
		.din(new_net_5291),
		.dout(new_net_5292)
	);

	bfr new_net_5293_bfr_after (
		.din(new_net_5292),
		.dout(new_net_5293)
	);

	bfr new_net_5294_bfr_after (
		.din(new_net_5293),
		.dout(new_net_5294)
	);

	bfr new_net_5295_bfr_after (
		.din(new_net_5294),
		.dout(new_net_5295)
	);

	bfr new_net_5296_bfr_after (
		.din(new_net_5295),
		.dout(new_net_5296)
	);

	bfr new_net_2173_bfr_after (
		.din(new_net_5296),
		.dout(new_net_2173)
	);

	bfr new_net_2236_bfr_after (
		.din(G134),
		.dout(new_net_2236)
	);

	bfr new_net_5297_bfr_after (
		.din(_0463_),
		.dout(new_net_5297)
	);

	bfr new_net_2320_bfr_after (
		.din(new_net_5297),
		.dout(new_net_2320)
	);

	bfr new_net_5298_bfr_after (
		.din(new_net_2375),
		.dout(new_net_5298)
	);

	bfr new_net_5299_bfr_after (
		.din(new_net_5298),
		.dout(new_net_5299)
	);

	bfr new_net_5300_bfr_after (
		.din(new_net_5299),
		.dout(new_net_5300)
	);

	bfr new_net_5301_bfr_after (
		.din(new_net_5300),
		.dout(new_net_5301)
	);

	bfr new_net_5302_bfr_after (
		.din(new_net_5301),
		.dout(new_net_5302)
	);

	bfr new_net_5303_bfr_after (
		.din(new_net_5302),
		.dout(new_net_5303)
	);

	bfr new_net_5304_bfr_after (
		.din(new_net_5303),
		.dout(new_net_5304)
	);

	bfr new_net_5305_bfr_after (
		.din(new_net_5304),
		.dout(new_net_5305)
	);

	bfr new_net_5306_bfr_after (
		.din(new_net_5305),
		.dout(new_net_5306)
	);

	bfr new_net_5307_bfr_after (
		.din(new_net_5306),
		.dout(new_net_5307)
	);

	bfr new_net_5308_bfr_after (
		.din(new_net_5307),
		.dout(new_net_5308)
	);

	bfr new_net_5309_bfr_after (
		.din(new_net_5308),
		.dout(new_net_5309)
	);

	bfr new_net_5310_bfr_after (
		.din(new_net_5309),
		.dout(new_net_5310)
	);

	bfr new_net_5311_bfr_after (
		.din(new_net_5310),
		.dout(new_net_5311)
	);

	bfr new_net_5312_bfr_after (
		.din(new_net_5311),
		.dout(new_net_5312)
	);

	bfr new_net_5313_bfr_after (
		.din(new_net_5312),
		.dout(new_net_5313)
	);

	bfr new_net_5314_bfr_after (
		.din(new_net_5313),
		.dout(new_net_5314)
	);

	bfr new_net_5315_bfr_after (
		.din(new_net_5314),
		.dout(new_net_5315)
	);

	bfr new_net_5316_bfr_after (
		.din(new_net_5315),
		.dout(new_net_5316)
	);

	bfr new_net_5317_bfr_after (
		.din(new_net_5316),
		.dout(new_net_5317)
	);

	bfr new_net_5318_bfr_after (
		.din(new_net_5317),
		.dout(new_net_5318)
	);

	bfr new_net_5319_bfr_after (
		.din(new_net_5318),
		.dout(new_net_5319)
	);

	bfr new_net_5320_bfr_after (
		.din(new_net_5319),
		.dout(new_net_5320)
	);

	bfr new_net_5321_bfr_after (
		.din(new_net_5320),
		.dout(new_net_5321)
	);

	bfr new_net_5322_bfr_after (
		.din(new_net_5321),
		.dout(new_net_5322)
	);

	bfr new_net_5323_bfr_after (
		.din(new_net_5322),
		.dout(new_net_5323)
	);

	bfr new_net_5324_bfr_after (
		.din(new_net_5323),
		.dout(new_net_5324)
	);

	bfr new_net_5325_bfr_after (
		.din(new_net_5324),
		.dout(new_net_5325)
	);

	bfr new_net_5326_bfr_after (
		.din(new_net_5325),
		.dout(new_net_5326)
	);

	bfr new_net_5327_bfr_after (
		.din(new_net_5326),
		.dout(new_net_5327)
	);

	bfr new_net_5328_bfr_after (
		.din(new_net_5327),
		.dout(new_net_5328)
	);

	bfr new_net_5329_bfr_after (
		.din(new_net_5328),
		.dout(new_net_5329)
	);

	bfr new_net_5330_bfr_after (
		.din(new_net_5329),
		.dout(new_net_5330)
	);

	bfr new_net_5331_bfr_after (
		.din(new_net_5330),
		.dout(new_net_5331)
	);

	bfr new_net_5332_bfr_after (
		.din(new_net_5331),
		.dout(new_net_5332)
	);

	bfr new_net_5333_bfr_after (
		.din(new_net_5332),
		.dout(new_net_5333)
	);

	bfr new_net_5334_bfr_after (
		.din(new_net_5333),
		.dout(new_net_5334)
	);

	bfr new_net_5335_bfr_after (
		.din(new_net_5334),
		.dout(new_net_5335)
	);

	bfr new_net_5336_bfr_after (
		.din(new_net_5335),
		.dout(new_net_5336)
	);

	bfr G5209_bfr_after (
		.din(new_net_5336),
		.dout(G5209)
	);

	bfr new_net_5337_bfr_after (
		.din(_0228_),
		.dout(new_net_5337)
	);

	bfr new_net_2257_bfr_after (
		.din(new_net_5337),
		.dout(new_net_2257)
	);

	bfr new_net_5338_bfr_after (
		.din(new_net_2351),
		.dout(new_net_5338)
	);

	bfr new_net_5339_bfr_after (
		.din(new_net_5338),
		.dout(new_net_5339)
	);

	bfr new_net_5340_bfr_after (
		.din(new_net_5339),
		.dout(new_net_5340)
	);

	bfr new_net_5341_bfr_after (
		.din(new_net_5340),
		.dout(new_net_5341)
	);

	bfr new_net_5342_bfr_after (
		.din(new_net_5341),
		.dout(new_net_5342)
	);

	bfr new_net_5343_bfr_after (
		.din(new_net_5342),
		.dout(new_net_5343)
	);

	bfr new_net_5344_bfr_after (
		.din(new_net_5343),
		.dout(new_net_5344)
	);

	bfr new_net_5345_bfr_after (
		.din(new_net_5344),
		.dout(new_net_5345)
	);

	bfr new_net_5346_bfr_after (
		.din(new_net_5345),
		.dout(new_net_5346)
	);

	bfr new_net_5347_bfr_after (
		.din(new_net_5346),
		.dout(new_net_5347)
	);

	bfr new_net_5348_bfr_after (
		.din(new_net_5347),
		.dout(new_net_5348)
	);

	bfr new_net_5349_bfr_after (
		.din(new_net_5348),
		.dout(new_net_5349)
	);

	bfr new_net_5350_bfr_after (
		.din(new_net_5349),
		.dout(new_net_5350)
	);

	bfr new_net_5351_bfr_after (
		.din(new_net_5350),
		.dout(new_net_5351)
	);

	bfr new_net_5352_bfr_after (
		.din(new_net_5351),
		.dout(new_net_5352)
	);

	bfr new_net_5353_bfr_after (
		.din(new_net_5352),
		.dout(new_net_5353)
	);

	bfr new_net_5354_bfr_after (
		.din(new_net_5353),
		.dout(new_net_5354)
	);

	bfr new_net_5355_bfr_after (
		.din(new_net_5354),
		.dout(new_net_5355)
	);

	bfr new_net_5356_bfr_after (
		.din(new_net_5355),
		.dout(new_net_5356)
	);

	bfr new_net_5357_bfr_after (
		.din(new_net_5356),
		.dout(new_net_5357)
	);

	bfr new_net_5358_bfr_after (
		.din(new_net_5357),
		.dout(new_net_5358)
	);

	bfr new_net_5359_bfr_after (
		.din(new_net_5358),
		.dout(new_net_5359)
	);

	bfr new_net_5360_bfr_after (
		.din(new_net_5359),
		.dout(new_net_5360)
	);

	bfr new_net_5361_bfr_after (
		.din(new_net_5360),
		.dout(new_net_5361)
	);

	bfr new_net_5362_bfr_after (
		.din(new_net_5361),
		.dout(new_net_5362)
	);

	bfr new_net_5363_bfr_after (
		.din(new_net_5362),
		.dout(new_net_5363)
	);

	bfr new_net_5364_bfr_after (
		.din(new_net_5363),
		.dout(new_net_5364)
	);

	bfr new_net_5365_bfr_after (
		.din(new_net_5364),
		.dout(new_net_5365)
	);

	bfr new_net_5366_bfr_after (
		.din(new_net_5365),
		.dout(new_net_5366)
	);

	bfr new_net_5367_bfr_after (
		.din(new_net_5366),
		.dout(new_net_5367)
	);

	bfr new_net_5368_bfr_after (
		.din(new_net_5367),
		.dout(new_net_5368)
	);

	bfr new_net_5369_bfr_after (
		.din(new_net_5368),
		.dout(new_net_5369)
	);

	bfr new_net_5370_bfr_after (
		.din(new_net_5369),
		.dout(new_net_5370)
	);

	bfr new_net_5371_bfr_after (
		.din(new_net_5370),
		.dout(new_net_5371)
	);

	bfr new_net_5372_bfr_after (
		.din(new_net_5371),
		.dout(new_net_5372)
	);

	bfr new_net_5373_bfr_after (
		.din(new_net_5372),
		.dout(new_net_5373)
	);

	bfr G5220_bfr_after (
		.din(new_net_5373),
		.dout(G5220)
	);

	bfr new_net_5374_bfr_after (
		.din(new_net_2399),
		.dout(new_net_5374)
	);

	bfr new_net_5375_bfr_after (
		.din(new_net_5374),
		.dout(new_net_5375)
	);

	bfr new_net_5376_bfr_after (
		.din(new_net_5375),
		.dout(new_net_5376)
	);

	bfr new_net_5377_bfr_after (
		.din(new_net_5376),
		.dout(new_net_5377)
	);

	bfr new_net_5378_bfr_after (
		.din(new_net_5377),
		.dout(new_net_5378)
	);

	bfr new_net_5379_bfr_after (
		.din(new_net_5378),
		.dout(new_net_5379)
	);

	bfr new_net_5380_bfr_after (
		.din(new_net_5379),
		.dout(new_net_5380)
	);

	bfr new_net_5381_bfr_after (
		.din(new_net_5380),
		.dout(new_net_5381)
	);

	bfr new_net_5382_bfr_after (
		.din(new_net_5381),
		.dout(new_net_5382)
	);

	bfr new_net_5383_bfr_after (
		.din(new_net_5382),
		.dout(new_net_5383)
	);

	bfr new_net_5384_bfr_after (
		.din(new_net_5383),
		.dout(new_net_5384)
	);

	bfr new_net_5385_bfr_after (
		.din(new_net_5384),
		.dout(new_net_5385)
	);

	bfr new_net_5386_bfr_after (
		.din(new_net_5385),
		.dout(new_net_5386)
	);

	bfr new_net_5387_bfr_after (
		.din(new_net_5386),
		.dout(new_net_5387)
	);

	bfr new_net_5388_bfr_after (
		.din(new_net_5387),
		.dout(new_net_5388)
	);

	bfr new_net_5389_bfr_after (
		.din(new_net_5388),
		.dout(new_net_5389)
	);

	bfr new_net_5390_bfr_after (
		.din(new_net_5389),
		.dout(new_net_5390)
	);

	bfr new_net_5391_bfr_after (
		.din(new_net_5390),
		.dout(new_net_5391)
	);

	bfr new_net_5392_bfr_after (
		.din(new_net_5391),
		.dout(new_net_5392)
	);

	bfr new_net_5393_bfr_after (
		.din(new_net_5392),
		.dout(new_net_5393)
	);

	bfr new_net_5394_bfr_after (
		.din(new_net_5393),
		.dout(new_net_5394)
	);

	bfr new_net_5395_bfr_after (
		.din(new_net_5394),
		.dout(new_net_5395)
	);

	bfr new_net_5396_bfr_after (
		.din(new_net_5395),
		.dout(new_net_5396)
	);

	bfr new_net_5397_bfr_after (
		.din(new_net_5396),
		.dout(new_net_5397)
	);

	bfr new_net_5398_bfr_after (
		.din(new_net_5397),
		.dout(new_net_5398)
	);

	bfr new_net_5399_bfr_after (
		.din(new_net_5398),
		.dout(new_net_5399)
	);

	bfr new_net_5400_bfr_after (
		.din(new_net_5399),
		.dout(new_net_5400)
	);

	bfr new_net_5401_bfr_after (
		.din(new_net_5400),
		.dout(new_net_5401)
	);

	bfr new_net_5402_bfr_after (
		.din(new_net_5401),
		.dout(new_net_5402)
	);

	bfr new_net_5403_bfr_after (
		.din(new_net_5402),
		.dout(new_net_5403)
	);

	bfr new_net_5404_bfr_after (
		.din(new_net_5403),
		.dout(new_net_5404)
	);

	bfr new_net_5405_bfr_after (
		.din(new_net_5404),
		.dout(new_net_5405)
	);

	bfr new_net_5406_bfr_after (
		.din(new_net_5405),
		.dout(new_net_5406)
	);

	bfr new_net_5407_bfr_after (
		.din(new_net_5406),
		.dout(new_net_5407)
	);

	bfr G5232_bfr_after (
		.din(new_net_5407),
		.dout(G5232)
	);

	bfr new_net_2110_bfr_after (
		.din(G12),
		.dout(new_net_2110)
	);

	bfr new_net_5408_bfr_after (
		.din(_0656_),
		.dout(new_net_5408)
	);

	bfr new_net_5409_bfr_after (
		.din(new_net_5408),
		.dout(new_net_5409)
	);

	bfr new_net_5410_bfr_after (
		.din(new_net_5409),
		.dout(new_net_5410)
	);

	bfr new_net_5411_bfr_after (
		.din(new_net_5410),
		.dout(new_net_5411)
	);

	bfr new_net_2131_bfr_after (
		.din(new_net_5411),
		.dout(new_net_2131)
	);

	bfr new_net_5412_bfr_after (
		.din(_1006_),
		.dout(new_net_5412)
	);

	bfr new_net_5413_bfr_after (
		.din(new_net_5412),
		.dout(new_net_5413)
	);

	bfr new_net_5414_bfr_after (
		.din(new_net_5413),
		.dout(new_net_5414)
	);

	bfr new_net_5415_bfr_after (
		.din(new_net_5414),
		.dout(new_net_5415)
	);

	bfr new_net_5416_bfr_after (
		.din(new_net_5415),
		.dout(new_net_5416)
	);

	bfr new_net_5417_bfr_after (
		.din(new_net_5416),
		.dout(new_net_5417)
	);

	bfr new_net_5418_bfr_after (
		.din(new_net_5417),
		.dout(new_net_5418)
	);

	bfr new_net_5419_bfr_after (
		.din(new_net_5418),
		.dout(new_net_5419)
	);

	bfr new_net_5420_bfr_after (
		.din(new_net_5419),
		.dout(new_net_5420)
	);

	bfr new_net_5421_bfr_after (
		.din(new_net_5420),
		.dout(new_net_5421)
	);

	bfr new_net_5422_bfr_after (
		.din(new_net_5421),
		.dout(new_net_5422)
	);

	bfr new_net_5423_bfr_after (
		.din(new_net_5422),
		.dout(new_net_5423)
	);

	bfr new_net_5424_bfr_after (
		.din(new_net_5423),
		.dout(new_net_5424)
	);

	bfr new_net_5425_bfr_after (
		.din(new_net_5424),
		.dout(new_net_5425)
	);

	bfr new_net_5426_bfr_after (
		.din(new_net_5425),
		.dout(new_net_5426)
	);

	bfr new_net_5427_bfr_after (
		.din(new_net_5426),
		.dout(new_net_5427)
	);

	bfr new_net_5428_bfr_after (
		.din(new_net_5427),
		.dout(new_net_5428)
	);

	bfr new_net_5429_bfr_after (
		.din(new_net_5428),
		.dout(new_net_5429)
	);

	bfr new_net_5430_bfr_after (
		.din(new_net_5429),
		.dout(new_net_5430)
	);

	bfr new_net_5431_bfr_after (
		.din(new_net_5430),
		.dout(new_net_5431)
	);

	bfr new_net_2194_bfr_after (
		.din(new_net_5431),
		.dout(new_net_2194)
	);

	bfr new_net_5432_bfr_after (
		.din(_0295_),
		.dout(new_net_5432)
	);

	bfr new_net_5433_bfr_after (
		.din(new_net_5432),
		.dout(new_net_5433)
	);

	bfr new_net_2278_bfr_after (
		.din(new_net_5433),
		.dout(new_net_2278)
	);

	bfr new_net_5434_bfr_after (
		.din(G51),
		.dout(new_net_5434)
	);

	bfr new_net_5435_bfr_after (
		.din(new_net_5434),
		.dout(new_net_5435)
	);

	bfr new_net_5436_bfr_after (
		.din(new_net_5435),
		.dout(new_net_5436)
	);

	bfr new_net_5437_bfr_after (
		.din(new_net_5436),
		.dout(new_net_5437)
	);

	bfr new_net_2341_bfr_after (
		.din(new_net_5437),
		.dout(new_net_2341)
	);

	bfr new_net_2212_bfr_after (
		.din(_1117_),
		.dout(new_net_2212)
	);

	bfr new_net_5438_bfr_after (
		.din(new_net_2465),
		.dout(new_net_5438)
	);

	bfr new_net_5439_bfr_after (
		.din(new_net_5438),
		.dout(new_net_5439)
	);

	bfr new_net_5440_bfr_after (
		.din(new_net_5439),
		.dout(new_net_5440)
	);

	bfr new_net_5441_bfr_after (
		.din(new_net_5440),
		.dout(new_net_5441)
	);

	bfr new_net_5442_bfr_after (
		.din(new_net_5441),
		.dout(new_net_5442)
	);

	bfr new_net_5443_bfr_after (
		.din(new_net_5442),
		.dout(new_net_5443)
	);

	bfr new_net_5444_bfr_after (
		.din(new_net_5443),
		.dout(new_net_5444)
	);

	bfr new_net_5445_bfr_after (
		.din(new_net_5444),
		.dout(new_net_5445)
	);

	bfr new_net_5446_bfr_after (
		.din(new_net_5445),
		.dout(new_net_5446)
	);

	bfr new_net_5447_bfr_after (
		.din(new_net_5446),
		.dout(new_net_5447)
	);

	bfr new_net_5448_bfr_after (
		.din(new_net_5447),
		.dout(new_net_5448)
	);

	bfr new_net_5449_bfr_after (
		.din(new_net_5448),
		.dout(new_net_5449)
	);

	bfr new_net_5450_bfr_after (
		.din(new_net_5449),
		.dout(new_net_5450)
	);

	bfr new_net_5451_bfr_after (
		.din(new_net_5450),
		.dout(new_net_5451)
	);

	bfr new_net_5452_bfr_after (
		.din(new_net_5451),
		.dout(new_net_5452)
	);

	bfr new_net_5453_bfr_after (
		.din(new_net_5452),
		.dout(new_net_5453)
	);

	bfr new_net_5454_bfr_after (
		.din(new_net_5453),
		.dout(new_net_5454)
	);

	bfr new_net_5455_bfr_after (
		.din(new_net_5454),
		.dout(new_net_5455)
	);

	bfr new_net_5456_bfr_after (
		.din(new_net_5455),
		.dout(new_net_5456)
	);

	bfr new_net_5457_bfr_after (
		.din(new_net_5456),
		.dout(new_net_5457)
	);

	bfr new_net_5458_bfr_after (
		.din(new_net_5457),
		.dout(new_net_5458)
	);

	bfr new_net_5459_bfr_after (
		.din(new_net_5458),
		.dout(new_net_5459)
	);

	bfr new_net_5460_bfr_after (
		.din(new_net_5459),
		.dout(new_net_5460)
	);

	bfr new_net_5461_bfr_after (
		.din(new_net_5460),
		.dout(new_net_5461)
	);

	bfr new_net_5462_bfr_after (
		.din(new_net_5461),
		.dout(new_net_5462)
	);

	bfr new_net_5463_bfr_after (
		.din(new_net_5462),
		.dout(new_net_5463)
	);

	bfr new_net_5464_bfr_after (
		.din(new_net_5463),
		.dout(new_net_5464)
	);

	bfr new_net_5465_bfr_after (
		.din(new_net_5464),
		.dout(new_net_5465)
	);

	bfr new_net_5466_bfr_after (
		.din(new_net_5465),
		.dout(new_net_5466)
	);

	bfr new_net_5467_bfr_after (
		.din(new_net_5466),
		.dout(new_net_5467)
	);

	bfr new_net_5468_bfr_after (
		.din(new_net_5467),
		.dout(new_net_5468)
	);

	bfr new_net_5469_bfr_after (
		.din(new_net_5468),
		.dout(new_net_5469)
	);

	bfr new_net_5470_bfr_after (
		.din(new_net_5469),
		.dout(new_net_5470)
	);

	bfr new_net_5471_bfr_after (
		.din(new_net_5470),
		.dout(new_net_5471)
	);

	bfr new_net_5472_bfr_after (
		.din(new_net_5471),
		.dout(new_net_5472)
	);

	bfr new_net_5473_bfr_after (
		.din(new_net_5472),
		.dout(new_net_5473)
	);

	bfr new_net_5474_bfr_after (
		.din(new_net_5473),
		.dout(new_net_5474)
	);

	bfr new_net_5475_bfr_after (
		.din(new_net_5474),
		.dout(new_net_5475)
	);

	bfr new_net_5476_bfr_after (
		.din(new_net_5475),
		.dout(new_net_5476)
	);

	bfr G5204_bfr_after (
		.din(new_net_5476),
		.dout(G5204)
	);

	bfr new_net_2109_bfr_after (
		.din(G164),
		.dout(new_net_2109)
	);

	bfr new_net_2210_bfr_after (
		.din(_1109_),
		.dout(new_net_2210)
	);

	bfr new_net_5477_bfr_after (
		.din(_0086_),
		.dout(new_net_5477)
	);

	bfr new_net_5478_bfr_after (
		.din(new_net_5477),
		.dout(new_net_5478)
	);

	bfr new_net_5479_bfr_after (
		.din(new_net_5478),
		.dout(new_net_5479)
	);

	bfr new_net_5480_bfr_after (
		.din(new_net_5479),
		.dout(new_net_5480)
	);

	bfr new_net_5481_bfr_after (
		.din(new_net_5480),
		.dout(new_net_5481)
	);

	bfr new_net_5482_bfr_after (
		.din(new_net_5481),
		.dout(new_net_5482)
	);

	bfr new_net_5483_bfr_after (
		.din(new_net_5482),
		.dout(new_net_5483)
	);

	bfr new_net_5484_bfr_after (
		.din(new_net_5483),
		.dout(new_net_5484)
	);

	bfr new_net_5485_bfr_after (
		.din(new_net_5484),
		.dout(new_net_5485)
	);

	bfr new_net_5486_bfr_after (
		.din(new_net_5485),
		.dout(new_net_5486)
	);

	bfr new_net_5487_bfr_after (
		.din(new_net_5486),
		.dout(new_net_5487)
	);

	bfr new_net_5488_bfr_after (
		.din(new_net_5487),
		.dout(new_net_5488)
	);

	bfr new_net_5489_bfr_after (
		.din(new_net_5488),
		.dout(new_net_5489)
	);

	bfr new_net_5490_bfr_after (
		.din(new_net_5489),
		.dout(new_net_5490)
	);

	bfr new_net_5491_bfr_after (
		.din(new_net_5490),
		.dout(new_net_5491)
	);

	bfr new_net_5492_bfr_after (
		.din(new_net_5491),
		.dout(new_net_5492)
	);

	bfr new_net_5493_bfr_after (
		.din(new_net_5492),
		.dout(new_net_5493)
	);

	bfr new_net_5494_bfr_after (
		.din(new_net_5493),
		.dout(new_net_5494)
	);

	bfr new_net_5495_bfr_after (
		.din(new_net_5494),
		.dout(new_net_5495)
	);

	bfr new_net_5496_bfr_after (
		.din(new_net_5495),
		.dout(new_net_5496)
	);

	bfr new_net_5497_bfr_after (
		.din(new_net_5496),
		.dout(new_net_5497)
	);

	bfr new_net_5498_bfr_after (
		.din(new_net_5497),
		.dout(new_net_5498)
	);

	bfr new_net_5499_bfr_after (
		.din(new_net_5498),
		.dout(new_net_5499)
	);

	bfr new_net_5500_bfr_after (
		.din(new_net_5499),
		.dout(new_net_5500)
	);

	bfr new_net_5501_bfr_after (
		.din(new_net_5500),
		.dout(new_net_5501)
	);

	bfr new_net_5502_bfr_after (
		.din(new_net_5501),
		.dout(new_net_5502)
	);

	bfr new_net_5503_bfr_after (
		.din(new_net_5502),
		.dout(new_net_5503)
	);

	bfr new_net_5504_bfr_after (
		.din(new_net_5503),
		.dout(new_net_5504)
	);

	bfr new_net_2231_bfr_after (
		.din(new_net_5504),
		.dout(new_net_2231)
	);

	bfr new_net_2252_bfr_after (
		.din(_0225_),
		.dout(new_net_2252)
	);

	bfr new_net_5505_bfr_after (
		.din(_0448_),
		.dout(new_net_5505)
	);

	bfr new_net_5506_bfr_after (
		.din(new_net_5505),
		.dout(new_net_5506)
	);

	bfr new_net_5507_bfr_after (
		.din(new_net_5506),
		.dout(new_net_5507)
	);

	bfr new_net_5508_bfr_after (
		.din(new_net_5507),
		.dout(new_net_5508)
	);

	bfr new_net_5509_bfr_after (
		.din(new_net_5508),
		.dout(new_net_5509)
	);

	bfr new_net_5510_bfr_after (
		.din(new_net_5509),
		.dout(new_net_5510)
	);

	bfr new_net_5511_bfr_after (
		.din(new_net_5510),
		.dout(new_net_5511)
	);

	bfr new_net_5512_bfr_after (
		.din(new_net_5511),
		.dout(new_net_5512)
	);

	bfr new_net_5513_bfr_after (
		.din(new_net_5512),
		.dout(new_net_5513)
	);

	bfr new_net_5514_bfr_after (
		.din(new_net_5513),
		.dout(new_net_5514)
	);

	bfr new_net_5515_bfr_after (
		.din(new_net_5514),
		.dout(new_net_5515)
	);

	bfr new_net_5516_bfr_after (
		.din(new_net_5515),
		.dout(new_net_5516)
	);

	bfr new_net_5517_bfr_after (
		.din(new_net_5516),
		.dout(new_net_5517)
	);

	bfr new_net_5518_bfr_after (
		.din(new_net_5517),
		.dout(new_net_5518)
	);

	bfr new_net_5519_bfr_after (
		.din(new_net_5518),
		.dout(new_net_5519)
	);

	bfr new_net_5520_bfr_after (
		.din(new_net_5519),
		.dout(new_net_5520)
	);

	bfr new_net_5521_bfr_after (
		.din(new_net_5520),
		.dout(new_net_5521)
	);

	bfr new_net_5522_bfr_after (
		.din(new_net_5521),
		.dout(new_net_5522)
	);

	bfr new_net_5523_bfr_after (
		.din(new_net_5522),
		.dout(new_net_5523)
	);

	bfr new_net_5524_bfr_after (
		.din(new_net_5523),
		.dout(new_net_5524)
	);

	bfr new_net_5525_bfr_after (
		.din(new_net_5524),
		.dout(new_net_5525)
	);

	bfr new_net_5526_bfr_after (
		.din(new_net_5525),
		.dout(new_net_5526)
	);

	bfr new_net_5527_bfr_after (
		.din(new_net_5526),
		.dout(new_net_5527)
	);

	bfr new_net_5528_bfr_after (
		.din(new_net_5527),
		.dout(new_net_5528)
	);

	bfr new_net_5529_bfr_after (
		.din(new_net_5528),
		.dout(new_net_5529)
	);

	bfr new_net_5530_bfr_after (
		.din(new_net_5529),
		.dout(new_net_5530)
	);

	bfr new_net_5531_bfr_after (
		.din(new_net_5530),
		.dout(new_net_5531)
	);

	bfr new_net_5532_bfr_after (
		.din(new_net_5531),
		.dout(new_net_5532)
	);

	bfr new_net_5533_bfr_after (
		.din(new_net_5532),
		.dout(new_net_5533)
	);

	bfr new_net_5534_bfr_after (
		.din(new_net_5533),
		.dout(new_net_5534)
	);

	bfr new_net_2315_bfr_after (
		.din(new_net_5534),
		.dout(new_net_2315)
	);

	bfr new_net_2273_bfr_after (
		.din(_0281_),
		.dout(new_net_2273)
	);

	bfr new_net_5535_bfr_after (
		.din(_0544_),
		.dout(new_net_5535)
	);

	bfr new_net_5536_bfr_after (
		.din(new_net_5535),
		.dout(new_net_5536)
	);

	bfr new_net_5537_bfr_after (
		.din(new_net_5536),
		.dout(new_net_5537)
	);

	bfr new_net_5538_bfr_after (
		.din(new_net_5537),
		.dout(new_net_5538)
	);

	bfr new_net_5539_bfr_after (
		.din(new_net_5538),
		.dout(new_net_5539)
	);

	bfr new_net_5540_bfr_after (
		.din(new_net_5539),
		.dout(new_net_5540)
	);

	bfr new_net_5541_bfr_after (
		.din(new_net_5540),
		.dout(new_net_5541)
	);

	bfr new_net_5542_bfr_after (
		.din(new_net_5541),
		.dout(new_net_5542)
	);

	bfr new_net_5543_bfr_after (
		.din(new_net_5542),
		.dout(new_net_5543)
	);

	bfr new_net_5544_bfr_after (
		.din(new_net_5543),
		.dout(new_net_5544)
	);

	bfr new_net_5545_bfr_after (
		.din(new_net_5544),
		.dout(new_net_5545)
	);

	bfr new_net_5546_bfr_after (
		.din(new_net_5545),
		.dout(new_net_5546)
	);

	bfr new_net_5547_bfr_after (
		.din(new_net_5546),
		.dout(new_net_5547)
	);

	bfr new_net_5548_bfr_after (
		.din(new_net_5547),
		.dout(new_net_5548)
	);

	bfr new_net_5549_bfr_after (
		.din(new_net_5548),
		.dout(new_net_5549)
	);

	bfr new_net_5550_bfr_after (
		.din(new_net_5549),
		.dout(new_net_5550)
	);

	bfr new_net_5551_bfr_after (
		.din(new_net_5550),
		.dout(new_net_5551)
	);

	bfr new_net_5552_bfr_after (
		.din(new_net_5551),
		.dout(new_net_5552)
	);

	bfr new_net_5553_bfr_after (
		.din(new_net_5552),
		.dout(new_net_5553)
	);

	bfr new_net_5554_bfr_after (
		.din(new_net_5553),
		.dout(new_net_5554)
	);

	bfr new_net_5555_bfr_after (
		.din(new_net_5554),
		.dout(new_net_5555)
	);

	bfr new_net_5556_bfr_after (
		.din(new_net_5555),
		.dout(new_net_5556)
	);

	bfr new_net_5557_bfr_after (
		.din(new_net_5556),
		.dout(new_net_5557)
	);

	bfr new_net_5558_bfr_after (
		.din(new_net_5557),
		.dout(new_net_5558)
	);

	bfr new_net_5559_bfr_after (
		.din(new_net_5558),
		.dout(new_net_5559)
	);

	bfr new_net_5560_bfr_after (
		.din(new_net_5559),
		.dout(new_net_5560)
	);

	bfr new_net_5561_bfr_after (
		.din(new_net_5560),
		.dout(new_net_5561)
	);

	bfr new_net_5562_bfr_after (
		.din(new_net_5561),
		.dout(new_net_5562)
	);

	bfr new_net_5563_bfr_after (
		.din(new_net_5562),
		.dout(new_net_5563)
	);

	bfr new_net_5564_bfr_after (
		.din(new_net_5563),
		.dout(new_net_5564)
	);

	bfr new_net_2336_bfr_after (
		.din(new_net_5564),
		.dout(new_net_2336)
	);

	bfr new_net_5565_bfr_after (
		.din(_0608_),
		.dout(new_net_5565)
	);

	bfr new_net_5566_bfr_after (
		.din(new_net_5565),
		.dout(new_net_5566)
	);

	bfr new_net_5567_bfr_after (
		.din(new_net_5566),
		.dout(new_net_5567)
	);

	bfr new_net_5568_bfr_after (
		.din(new_net_5567),
		.dout(new_net_5568)
	);

	bfr new_net_5569_bfr_after (
		.din(new_net_5568),
		.dout(new_net_5569)
	);

	bfr new_net_5570_bfr_after (
		.din(new_net_5569),
		.dout(new_net_5570)
	);

	bfr new_net_5571_bfr_after (
		.din(new_net_5570),
		.dout(new_net_5571)
	);

	bfr new_net_5572_bfr_after (
		.din(new_net_5571),
		.dout(new_net_5572)
	);

	bfr new_net_5573_bfr_after (
		.din(new_net_5572),
		.dout(new_net_5573)
	);

	bfr new_net_5574_bfr_after (
		.din(new_net_5573),
		.dout(new_net_5574)
	);

	bfr new_net_2126_bfr_after (
		.din(new_net_5574),
		.dout(new_net_2126)
	);

	bfr new_net_5575_bfr_after (
		.din(G108),
		.dout(new_net_5575)
	);

	bfr new_net_2147_bfr_after (
		.din(new_net_5575),
		.dout(new_net_2147)
	);

	bfr new_net_5576_bfr_after (
		.din(_0857_),
		.dout(new_net_5576)
	);

	bfr new_net_5577_bfr_after (
		.din(new_net_5576),
		.dout(new_net_5577)
	);

	bfr new_net_5578_bfr_after (
		.din(new_net_5577),
		.dout(new_net_5578)
	);

	bfr new_net_5579_bfr_after (
		.din(new_net_5578),
		.dout(new_net_5579)
	);

	bfr new_net_2168_bfr_after (
		.din(new_net_5579),
		.dout(new_net_2168)
	);

	bfr new_net_5580_bfr_after (
		.din(G30),
		.dout(new_net_5580)
	);

	bfr new_net_2246_bfr_after (
		.din(new_net_5580),
		.dout(new_net_2246)
	);

	bfr new_net_5581_bfr_after (
		.din(_0407_),
		.dout(new_net_5581)
	);

	bfr new_net_5582_bfr_after (
		.din(new_net_5581),
		.dout(new_net_5582)
	);

	bfr new_net_2304_bfr_after (
		.din(new_net_5582),
		.dout(new_net_2304)
	);

	bfr new_net_5583_bfr_after (
		.din(_0429_),
		.dout(new_net_5583)
	);

	bfr new_net_5584_bfr_after (
		.din(new_net_5583),
		.dout(new_net_5584)
	);

	bfr new_net_5585_bfr_after (
		.din(new_net_5584),
		.dout(new_net_5585)
	);

	bfr new_net_5586_bfr_after (
		.din(new_net_5585),
		.dout(new_net_5586)
	);

	bfr new_net_2309_bfr_after (
		.din(new_net_5586),
		.dout(new_net_2309)
	);

	bfr new_net_5587_bfr_after (
		.din(new_net_2485),
		.dout(new_net_5587)
	);

	bfr new_net_5588_bfr_after (
		.din(new_net_5587),
		.dout(new_net_5588)
	);

	bfr new_net_5589_bfr_after (
		.din(new_net_5588),
		.dout(new_net_5589)
	);

	bfr new_net_5590_bfr_after (
		.din(new_net_5589),
		.dout(new_net_5590)
	);

	bfr new_net_5591_bfr_after (
		.din(new_net_5590),
		.dout(new_net_5591)
	);

	bfr new_net_5592_bfr_after (
		.din(new_net_5591),
		.dout(new_net_5592)
	);

	bfr new_net_5593_bfr_after (
		.din(new_net_5592),
		.dout(new_net_5593)
	);

	bfr new_net_5594_bfr_after (
		.din(new_net_5593),
		.dout(new_net_5594)
	);

	bfr new_net_5595_bfr_after (
		.din(new_net_5594),
		.dout(new_net_5595)
	);

	bfr new_net_5596_bfr_after (
		.din(new_net_5595),
		.dout(new_net_5596)
	);

	bfr new_net_5597_bfr_after (
		.din(new_net_5596),
		.dout(new_net_5597)
	);

	bfr new_net_5598_bfr_after (
		.din(new_net_5597),
		.dout(new_net_5598)
	);

	bfr new_net_5599_bfr_after (
		.din(new_net_5598),
		.dout(new_net_5599)
	);

	bfr new_net_5600_bfr_after (
		.din(new_net_5599),
		.dout(new_net_5600)
	);

	bfr new_net_5601_bfr_after (
		.din(new_net_5600),
		.dout(new_net_5601)
	);

	bfr new_net_5602_bfr_after (
		.din(new_net_5601),
		.dout(new_net_5602)
	);

	bfr new_net_5603_bfr_after (
		.din(new_net_5602),
		.dout(new_net_5603)
	);

	bfr new_net_5604_bfr_after (
		.din(new_net_5603),
		.dout(new_net_5604)
	);

	bfr new_net_5605_bfr_after (
		.din(new_net_5604),
		.dout(new_net_5605)
	);

	bfr new_net_5606_bfr_after (
		.din(new_net_5605),
		.dout(new_net_5606)
	);

	bfr new_net_5607_bfr_after (
		.din(new_net_5606),
		.dout(new_net_5607)
	);

	bfr new_net_5608_bfr_after (
		.din(new_net_5607),
		.dout(new_net_5608)
	);

	bfr new_net_5609_bfr_after (
		.din(new_net_5608),
		.dout(new_net_5609)
	);

	bfr new_net_5610_bfr_after (
		.din(new_net_5609),
		.dout(new_net_5610)
	);

	bfr new_net_5611_bfr_after (
		.din(new_net_5610),
		.dout(new_net_5611)
	);

	bfr G5283_bfr_after (
		.din(new_net_5611),
		.dout(G5283)
	);

	bfr new_net_5612_bfr_after (
		.din(G9),
		.dout(new_net_5612)
	);

	bfr new_net_2242_bfr_after (
		.din(new_net_5612),
		.dout(new_net_2242)
	);

	bfr new_net_2185_bfr_after (
		.din(_0939_),
		.dout(new_net_2185)
	);

	bfr new_net_2272_bfr_after (
		.din(_0280_),
		.dout(new_net_2272)
	);

	bfr new_net_5613_bfr_after (
		.din(_0536_),
		.dout(new_net_5613)
	);

	bfr new_net_5614_bfr_after (
		.din(new_net_5613),
		.dout(new_net_5614)
	);

	bfr new_net_5615_bfr_after (
		.din(new_net_5614),
		.dout(new_net_5615)
	);

	bfr new_net_5616_bfr_after (
		.din(new_net_5615),
		.dout(new_net_5616)
	);

	bfr new_net_5617_bfr_after (
		.din(new_net_5616),
		.dout(new_net_5617)
	);

	bfr new_net_5618_bfr_after (
		.din(new_net_5617),
		.dout(new_net_5618)
	);

	bfr new_net_5619_bfr_after (
		.din(new_net_5618),
		.dout(new_net_5619)
	);

	bfr new_net_5620_bfr_after (
		.din(new_net_5619),
		.dout(new_net_5620)
	);

	bfr new_net_5621_bfr_after (
		.din(new_net_5620),
		.dout(new_net_5621)
	);

	bfr new_net_5622_bfr_after (
		.din(new_net_5621),
		.dout(new_net_5622)
	);

	bfr new_net_5623_bfr_after (
		.din(new_net_5622),
		.dout(new_net_5623)
	);

	bfr new_net_5624_bfr_after (
		.din(new_net_5623),
		.dout(new_net_5624)
	);

	bfr new_net_5625_bfr_after (
		.din(new_net_5624),
		.dout(new_net_5625)
	);

	bfr new_net_5626_bfr_after (
		.din(new_net_5625),
		.dout(new_net_5626)
	);

	bfr new_net_5627_bfr_after (
		.din(new_net_5626),
		.dout(new_net_5627)
	);

	bfr new_net_5628_bfr_after (
		.din(new_net_5627),
		.dout(new_net_5628)
	);

	bfr new_net_5629_bfr_after (
		.din(new_net_5628),
		.dout(new_net_5629)
	);

	bfr new_net_5630_bfr_after (
		.din(new_net_5629),
		.dout(new_net_5630)
	);

	bfr new_net_5631_bfr_after (
		.din(new_net_5630),
		.dout(new_net_5631)
	);

	bfr new_net_5632_bfr_after (
		.din(new_net_5631),
		.dout(new_net_5632)
	);

	bfr new_net_5633_bfr_after (
		.din(new_net_5632),
		.dout(new_net_5633)
	);

	bfr new_net_5634_bfr_after (
		.din(new_net_5633),
		.dout(new_net_5634)
	);

	bfr new_net_5635_bfr_after (
		.din(new_net_5634),
		.dout(new_net_5635)
	);

	bfr new_net_5636_bfr_after (
		.din(new_net_5635),
		.dout(new_net_5636)
	);

	bfr new_net_5637_bfr_after (
		.din(new_net_5636),
		.dout(new_net_5637)
	);

	bfr new_net_5638_bfr_after (
		.din(new_net_5637),
		.dout(new_net_5638)
	);

	bfr new_net_5639_bfr_after (
		.din(new_net_5638),
		.dout(new_net_5639)
	);

	bfr new_net_2335_bfr_after (
		.din(new_net_5639),
		.dout(new_net_2335)
	);

	bfr new_net_5640_bfr_after (
		.din(_0765_),
		.dout(new_net_5640)
	);

	bfr new_net_5641_bfr_after (
		.din(new_net_5640),
		.dout(new_net_5641)
	);

	bfr new_net_2152_bfr_after (
		.din(new_net_5641),
		.dout(new_net_2152)
	);

	bfr new_net_5642_bfr_after (
		.din(_1223_),
		.dout(new_net_5642)
	);

	bfr new_net_5643_bfr_after (
		.din(new_net_5642),
		.dout(new_net_5643)
	);

	bfr new_net_5644_bfr_after (
		.din(new_net_5643),
		.dout(new_net_5644)
	);

	bfr new_net_5645_bfr_after (
		.din(new_net_5644),
		.dout(new_net_5645)
	);

	bfr new_net_5646_bfr_after (
		.din(new_net_5645),
		.dout(new_net_5646)
	);

	bfr new_net_5647_bfr_after (
		.din(new_net_5646),
		.dout(new_net_5647)
	);

	bfr new_net_5648_bfr_after (
		.din(new_net_5647),
		.dout(new_net_5648)
	);

	bfr new_net_5649_bfr_after (
		.din(new_net_5648),
		.dout(new_net_5649)
	);

	bfr new_net_5650_bfr_after (
		.din(new_net_5649),
		.dout(new_net_5650)
	);

	bfr new_net_5651_bfr_after (
		.din(new_net_5650),
		.dout(new_net_5651)
	);

	bfr new_net_5652_bfr_after (
		.din(new_net_5651),
		.dout(new_net_5652)
	);

	bfr new_net_2215_bfr_after (
		.din(new_net_5652),
		.dout(new_net_2215)
	);

	bfr new_net_5653_bfr_after (
		.din(_1111_),
		.dout(new_net_5653)
	);

	bfr new_net_5654_bfr_after (
		.din(new_net_5653),
		.dout(new_net_5654)
	);

	bfr new_net_2211_bfr_after (
		.din(new_net_5654),
		.dout(new_net_2211)
	);

	bfr new_net_5655_bfr_after (
		.din(_0593_),
		.dout(new_net_5655)
	);

	bfr new_net_5656_bfr_after (
		.din(new_net_5655),
		.dout(new_net_5656)
	);

	bfr new_net_5657_bfr_after (
		.din(new_net_5656),
		.dout(new_net_5657)
	);

	bfr new_net_5658_bfr_after (
		.din(new_net_5657),
		.dout(new_net_5658)
	);

	bfr new_net_5659_bfr_after (
		.din(new_net_5658),
		.dout(new_net_5659)
	);

	bfr new_net_2121_bfr_after (
		.din(new_net_5659),
		.dout(new_net_2121)
	);

	bfr new_net_5660_bfr_after (
		.din(_0730_),
		.dout(new_net_5660)
	);

	bfr new_net_5661_bfr_after (
		.din(new_net_5660),
		.dout(new_net_5661)
	);

	bfr new_net_5662_bfr_after (
		.din(new_net_5661),
		.dout(new_net_5662)
	);

	bfr new_net_5663_bfr_after (
		.din(new_net_5662),
		.dout(new_net_5663)
	);

	bfr new_net_5664_bfr_after (
		.din(new_net_5663),
		.dout(new_net_5664)
	);

	bfr new_net_5665_bfr_after (
		.din(new_net_5664),
		.dout(new_net_5665)
	);

	bfr new_net_5666_bfr_after (
		.din(new_net_5665),
		.dout(new_net_5666)
	);

	bfr new_net_5667_bfr_after (
		.din(new_net_5666),
		.dout(new_net_5667)
	);

	bfr new_net_5668_bfr_after (
		.din(new_net_5667),
		.dout(new_net_5668)
	);

	bfr new_net_2142_bfr_after (
		.din(new_net_5668),
		.dout(new_net_2142)
	);

	bfr new_net_5669_bfr_after (
		.din(_0813_),
		.dout(new_net_5669)
	);

	bfr new_net_5670_bfr_after (
		.din(new_net_5669),
		.dout(new_net_5670)
	);

	bfr new_net_5671_bfr_after (
		.din(new_net_5670),
		.dout(new_net_5671)
	);

	bfr new_net_5672_bfr_after (
		.din(new_net_5671),
		.dout(new_net_5672)
	);

	bfr new_net_5673_bfr_after (
		.din(new_net_5672),
		.dout(new_net_5673)
	);

	bfr new_net_5674_bfr_after (
		.din(new_net_5673),
		.dout(new_net_5674)
	);

	bfr new_net_5675_bfr_after (
		.din(new_net_5674),
		.dout(new_net_5675)
	);

	bfr new_net_5676_bfr_after (
		.din(new_net_5675),
		.dout(new_net_5676)
	);

	bfr new_net_5677_bfr_after (
		.din(new_net_5676),
		.dout(new_net_5677)
	);

	bfr new_net_5678_bfr_after (
		.din(new_net_5677),
		.dout(new_net_5678)
	);

	bfr new_net_5679_bfr_after (
		.din(new_net_5678),
		.dout(new_net_5679)
	);

	bfr new_net_5680_bfr_after (
		.din(new_net_5679),
		.dout(new_net_5680)
	);

	bfr new_net_5681_bfr_after (
		.din(new_net_5680),
		.dout(new_net_5681)
	);

	bfr new_net_5682_bfr_after (
		.din(new_net_5681),
		.dout(new_net_5682)
	);

	bfr new_net_5683_bfr_after (
		.din(new_net_5682),
		.dout(new_net_5683)
	);

	bfr new_net_5684_bfr_after (
		.din(new_net_5683),
		.dout(new_net_5684)
	);

	bfr new_net_5685_bfr_after (
		.din(new_net_5684),
		.dout(new_net_5685)
	);

	bfr new_net_2163_bfr_after (
		.din(new_net_5685),
		.dout(new_net_2163)
	);

	bfr new_net_5686_bfr_after (
		.din(G91),
		.dout(new_net_5686)
	);

	bfr new_net_2184_bfr_after (
		.din(new_net_5686),
		.dout(new_net_2184)
	);

	bfr new_net_5687_bfr_after (
		.din(_0342_),
		.dout(new_net_5687)
	);

	bfr new_net_5688_bfr_after (
		.din(new_net_5687),
		.dout(new_net_5688)
	);

	bfr new_net_5689_bfr_after (
		.din(new_net_5688),
		.dout(new_net_5689)
	);

	bfr new_net_5690_bfr_after (
		.din(new_net_5689),
		.dout(new_net_5690)
	);

	bfr new_net_5691_bfr_after (
		.din(new_net_5690),
		.dout(new_net_5691)
	);

	bfr new_net_5692_bfr_after (
		.din(new_net_5691),
		.dout(new_net_5692)
	);

	bfr new_net_5693_bfr_after (
		.din(new_net_5692),
		.dout(new_net_5693)
	);

	bfr new_net_5694_bfr_after (
		.din(new_net_5693),
		.dout(new_net_5694)
	);

	bfr new_net_5695_bfr_after (
		.din(new_net_5694),
		.dout(new_net_5695)
	);

	bfr new_net_5696_bfr_after (
		.din(new_net_5695),
		.dout(new_net_5696)
	);

	bfr new_net_5697_bfr_after (
		.din(new_net_5696),
		.dout(new_net_5697)
	);

	bfr new_net_5698_bfr_after (
		.din(new_net_5697),
		.dout(new_net_5698)
	);

	bfr new_net_5699_bfr_after (
		.din(new_net_5698),
		.dout(new_net_5699)
	);

	bfr new_net_5700_bfr_after (
		.din(new_net_5699),
		.dout(new_net_5700)
	);

	bfr new_net_5701_bfr_after (
		.din(new_net_5700),
		.dout(new_net_5701)
	);

	bfr new_net_5702_bfr_after (
		.din(new_net_5701),
		.dout(new_net_5702)
	);

	bfr new_net_5703_bfr_after (
		.din(new_net_5702),
		.dout(new_net_5703)
	);

	bfr new_net_5704_bfr_after (
		.din(new_net_5703),
		.dout(new_net_5704)
	);

	bfr new_net_5705_bfr_after (
		.din(new_net_5704),
		.dout(new_net_5705)
	);

	bfr new_net_5706_bfr_after (
		.din(new_net_5705),
		.dout(new_net_5706)
	);

	bfr new_net_5707_bfr_after (
		.din(new_net_5706),
		.dout(new_net_5707)
	);

	bfr new_net_5708_bfr_after (
		.din(new_net_5707),
		.dout(new_net_5708)
	);

	bfr new_net_2289_bfr_after (
		.din(new_net_5708),
		.dout(new_net_2289)
	);

	bfr new_net_2205_bfr_after (
		.din(_1058_),
		.dout(new_net_2205)
	);

	bfr new_net_2226_bfr_after (
		.din(_0072_),
		.dout(new_net_2226)
	);

	bfr new_net_5709_bfr_after (
		.din(G10),
		.dout(new_net_5709)
	);

	bfr new_net_2247_bfr_after (
		.din(new_net_5709),
		.dout(new_net_2247)
	);

	bfr new_net_5710_bfr_after (
		.din(_0428_),
		.dout(new_net_5710)
	);

	bfr new_net_5711_bfr_after (
		.din(new_net_5710),
		.dout(new_net_5711)
	);

	bfr new_net_5712_bfr_after (
		.din(new_net_5711),
		.dout(new_net_5712)
	);

	bfr new_net_5713_bfr_after (
		.din(new_net_5712),
		.dout(new_net_5713)
	);

	bfr new_net_5714_bfr_after (
		.din(new_net_5713),
		.dout(new_net_5714)
	);

	bfr new_net_5715_bfr_after (
		.din(new_net_5714),
		.dout(new_net_5715)
	);

	bfr new_net_5716_bfr_after (
		.din(new_net_5715),
		.dout(new_net_5716)
	);

	bfr new_net_2310_bfr_after (
		.din(new_net_5716),
		.dout(new_net_2310)
	);

	bfr new_net_5717_bfr_after (
		.din(_0274_),
		.dout(new_net_5717)
	);

	bfr new_net_2268_bfr_after (
		.din(new_net_5717),
		.dout(new_net_2268)
	);

	bfr new_net_5718_bfr_after (
		.din(_0254_),
		.dout(new_net_5718)
	);

	bfr new_net_5719_bfr_after (
		.din(new_net_5718),
		.dout(new_net_5719)
	);

	bfr new_net_2263_bfr_after (
		.din(new_net_5719),
		.dout(new_net_2263)
	);

	bfr new_net_5720_bfr_after (
		.din(_0658_),
		.dout(new_net_5720)
	);

	bfr new_net_5721_bfr_after (
		.din(new_net_5720),
		.dout(new_net_5721)
	);

	bfr new_net_5722_bfr_after (
		.din(new_net_5721),
		.dout(new_net_5722)
	);

	bfr new_net_5723_bfr_after (
		.din(new_net_5722),
		.dout(new_net_5723)
	);

	bfr new_net_5724_bfr_after (
		.din(new_net_5723),
		.dout(new_net_5724)
	);

	bfr new_net_5725_bfr_after (
		.din(new_net_5724),
		.dout(new_net_5725)
	);

	bfr new_net_5726_bfr_after (
		.din(new_net_5725),
		.dout(new_net_5726)
	);

	bfr new_net_5727_bfr_after (
		.din(new_net_5726),
		.dout(new_net_5727)
	);

	bfr new_net_5728_bfr_after (
		.din(new_net_5727),
		.dout(new_net_5728)
	);

	bfr new_net_5729_bfr_after (
		.din(new_net_5728),
		.dout(new_net_5729)
	);

	bfr new_net_5730_bfr_after (
		.din(new_net_5729),
		.dout(new_net_5730)
	);

	bfr new_net_5731_bfr_after (
		.din(new_net_5730),
		.dout(new_net_5731)
	);

	bfr new_net_5732_bfr_after (
		.din(new_net_5731),
		.dout(new_net_5732)
	);

	bfr new_net_5733_bfr_after (
		.din(new_net_5732),
		.dout(new_net_5733)
	);

	bfr new_net_5734_bfr_after (
		.din(new_net_5733),
		.dout(new_net_5734)
	);

	bfr new_net_5735_bfr_after (
		.din(new_net_5734),
		.dout(new_net_5735)
	);

	bfr new_net_5736_bfr_after (
		.din(new_net_5735),
		.dout(new_net_5736)
	);

	bfr new_net_2137_bfr_after (
		.din(new_net_5736),
		.dout(new_net_2137)
	);

	bfr new_net_5737_bfr_after (
		.din(_0811_),
		.dout(new_net_5737)
	);

	bfr new_net_5738_bfr_after (
		.din(new_net_5737),
		.dout(new_net_5738)
	);

	bfr new_net_5739_bfr_after (
		.din(new_net_5738),
		.dout(new_net_5739)
	);

	bfr new_net_5740_bfr_after (
		.din(new_net_5739),
		.dout(new_net_5740)
	);

	bfr new_net_5741_bfr_after (
		.din(new_net_5740),
		.dout(new_net_5741)
	);

	bfr new_net_5742_bfr_after (
		.din(new_net_5741),
		.dout(new_net_5742)
	);

	bfr new_net_5743_bfr_after (
		.din(new_net_5742),
		.dout(new_net_5743)
	);

	bfr new_net_5744_bfr_after (
		.din(new_net_5743),
		.dout(new_net_5744)
	);

	bfr new_net_5745_bfr_after (
		.din(new_net_5744),
		.dout(new_net_5745)
	);

	bfr new_net_5746_bfr_after (
		.din(new_net_5745),
		.dout(new_net_5746)
	);

	bfr new_net_5747_bfr_after (
		.din(new_net_5746),
		.dout(new_net_5747)
	);

	bfr new_net_5748_bfr_after (
		.din(new_net_5747),
		.dout(new_net_5748)
	);

	bfr new_net_2158_bfr_after (
		.din(new_net_5748),
		.dout(new_net_2158)
	);

	bfr new_net_5749_bfr_after (
		.din(G43),
		.dout(new_net_5749)
	);

	bfr new_net_5750_bfr_after (
		.din(new_net_5749),
		.dout(new_net_5750)
	);

	bfr new_net_5751_bfr_after (
		.din(new_net_5750),
		.dout(new_net_5751)
	);

	bfr new_net_5752_bfr_after (
		.din(new_net_5751),
		.dout(new_net_5752)
	);

	bfr new_net_2179_bfr_after (
		.din(new_net_5752),
		.dout(new_net_2179)
	);

	bfr new_net_5753_bfr_after (
		.din(G35),
		.dout(new_net_5753)
	);

	bfr new_net_2116_bfr_after (
		.din(new_net_5753),
		.dout(new_net_2116)
	);

	bfr new_net_5754_bfr_after (
		.din(_1044_),
		.dout(new_net_5754)
	);

	bfr new_net_5755_bfr_after (
		.din(new_net_5754),
		.dout(new_net_5755)
	);

	bfr new_net_5756_bfr_after (
		.din(new_net_5755),
		.dout(new_net_5756)
	);

	bfr new_net_5757_bfr_after (
		.din(new_net_5756),
		.dout(new_net_5757)
	);

	bfr new_net_5758_bfr_after (
		.din(new_net_5757),
		.dout(new_net_5758)
	);

	bfr new_net_5759_bfr_after (
		.din(new_net_5758),
		.dout(new_net_5759)
	);

	bfr new_net_5760_bfr_after (
		.din(new_net_5759),
		.dout(new_net_5760)
	);

	bfr new_net_5761_bfr_after (
		.din(new_net_5760),
		.dout(new_net_5761)
	);

	bfr new_net_5762_bfr_after (
		.din(new_net_5761),
		.dout(new_net_5762)
	);

	bfr new_net_5763_bfr_after (
		.din(new_net_5762),
		.dout(new_net_5763)
	);

	bfr new_net_5764_bfr_after (
		.din(new_net_5763),
		.dout(new_net_5764)
	);

	bfr new_net_5765_bfr_after (
		.din(new_net_5764),
		.dout(new_net_5765)
	);

	bfr new_net_5766_bfr_after (
		.din(new_net_5765),
		.dout(new_net_5766)
	);

	bfr new_net_5767_bfr_after (
		.din(new_net_5766),
		.dout(new_net_5767)
	);

	bfr new_net_5768_bfr_after (
		.din(new_net_5767),
		.dout(new_net_5768)
	);

	bfr new_net_5769_bfr_after (
		.din(new_net_5768),
		.dout(new_net_5769)
	);

	bfr new_net_5770_bfr_after (
		.din(new_net_5769),
		.dout(new_net_5770)
	);

	bfr new_net_5771_bfr_after (
		.din(new_net_5770),
		.dout(new_net_5771)
	);

	bfr new_net_2200_bfr_after (
		.din(new_net_5771),
		.dout(new_net_2200)
	);

	bfr new_net_5772_bfr_after (
		.din(_0321_),
		.dout(new_net_5772)
	);

	bfr new_net_5773_bfr_after (
		.din(new_net_5772),
		.dout(new_net_5773)
	);

	bfr new_net_5774_bfr_after (
		.din(new_net_5773),
		.dout(new_net_5774)
	);

	bfr new_net_5775_bfr_after (
		.din(new_net_5774),
		.dout(new_net_5775)
	);

	bfr new_net_5776_bfr_after (
		.din(new_net_5775),
		.dout(new_net_5776)
	);

	bfr new_net_5777_bfr_after (
		.din(new_net_5776),
		.dout(new_net_5777)
	);

	bfr new_net_5778_bfr_after (
		.din(new_net_5777),
		.dout(new_net_5778)
	);

	bfr new_net_5779_bfr_after (
		.din(new_net_5778),
		.dout(new_net_5779)
	);

	bfr new_net_5780_bfr_after (
		.din(new_net_5779),
		.dout(new_net_5780)
	);

	bfr new_net_5781_bfr_after (
		.din(new_net_5780),
		.dout(new_net_5781)
	);

	bfr new_net_5782_bfr_after (
		.din(new_net_5781),
		.dout(new_net_5782)
	);

	bfr new_net_5783_bfr_after (
		.din(new_net_5782),
		.dout(new_net_5783)
	);

	bfr new_net_5784_bfr_after (
		.din(new_net_5783),
		.dout(new_net_5784)
	);

	bfr new_net_5785_bfr_after (
		.din(new_net_5784),
		.dout(new_net_5785)
	);

	bfr new_net_5786_bfr_after (
		.din(new_net_5785),
		.dout(new_net_5786)
	);

	bfr new_net_5787_bfr_after (
		.din(new_net_5786),
		.dout(new_net_5787)
	);

	bfr new_net_5788_bfr_after (
		.din(new_net_5787),
		.dout(new_net_5788)
	);

	bfr new_net_5789_bfr_after (
		.din(new_net_5788),
		.dout(new_net_5789)
	);

	bfr new_net_5790_bfr_after (
		.din(new_net_5789),
		.dout(new_net_5790)
	);

	bfr new_net_5791_bfr_after (
		.din(new_net_5790),
		.dout(new_net_5791)
	);

	bfr new_net_5792_bfr_after (
		.din(new_net_5791),
		.dout(new_net_5792)
	);

	bfr new_net_5793_bfr_after (
		.din(new_net_5792),
		.dout(new_net_5793)
	);

	bfr new_net_2284_bfr_after (
		.din(new_net_5793),
		.dout(new_net_2284)
	);

	bfr new_net_5794_bfr_after (
		.din(_0573_),
		.dout(new_net_5794)
	);

	bfr new_net_5795_bfr_after (
		.din(new_net_5794),
		.dout(new_net_5795)
	);

	bfr new_net_2347_bfr_after (
		.din(new_net_5795),
		.dout(new_net_2347)
	);

	bfr new_net_5796_bfr_after (
		.din(_0002_),
		.dout(new_net_5796)
	);

	bfr new_net_5797_bfr_after (
		.din(new_net_5796),
		.dout(new_net_5797)
	);

	bfr new_net_5798_bfr_after (
		.din(new_net_5797),
		.dout(new_net_5798)
	);

	bfr new_net_5799_bfr_after (
		.din(new_net_5798),
		.dout(new_net_5799)
	);

	bfr new_net_5800_bfr_after (
		.din(new_net_5799),
		.dout(new_net_5800)
	);

	bfr new_net_5801_bfr_after (
		.din(new_net_5800),
		.dout(new_net_5801)
	);

	bfr new_net_5802_bfr_after (
		.din(new_net_5801),
		.dout(new_net_5802)
	);

	bfr new_net_5803_bfr_after (
		.din(new_net_5802),
		.dout(new_net_5803)
	);

	bfr new_net_2221_bfr_after (
		.din(new_net_5803),
		.dout(new_net_2221)
	);

	bfr new_net_5804_bfr_after (
		.din(_0411_),
		.dout(new_net_5804)
	);

	bfr new_net_5805_bfr_after (
		.din(new_net_5804),
		.dout(new_net_5805)
	);

	bfr new_net_5806_bfr_after (
		.din(new_net_5805),
		.dout(new_net_5806)
	);

	bfr new_net_5807_bfr_after (
		.din(new_net_5806),
		.dout(new_net_5807)
	);

	bfr new_net_5808_bfr_after (
		.din(new_net_5807),
		.dout(new_net_5808)
	);

	bfr new_net_5809_bfr_after (
		.din(new_net_5808),
		.dout(new_net_5809)
	);

	bfr new_net_5810_bfr_after (
		.din(new_net_5809),
		.dout(new_net_5810)
	);

	bfr new_net_5811_bfr_after (
		.din(new_net_5810),
		.dout(new_net_5811)
	);

	bfr new_net_5812_bfr_after (
		.din(new_net_5811),
		.dout(new_net_5812)
	);

	bfr new_net_5813_bfr_after (
		.din(new_net_5812),
		.dout(new_net_5813)
	);

	bfr new_net_5814_bfr_after (
		.din(new_net_5813),
		.dout(new_net_5814)
	);

	bfr new_net_5815_bfr_after (
		.din(new_net_5814),
		.dout(new_net_5815)
	);

	bfr new_net_5816_bfr_after (
		.din(new_net_5815),
		.dout(new_net_5816)
	);

	bfr new_net_5817_bfr_after (
		.din(new_net_5816),
		.dout(new_net_5817)
	);

	bfr new_net_5818_bfr_after (
		.din(new_net_5817),
		.dout(new_net_5818)
	);

	bfr new_net_5819_bfr_after (
		.din(new_net_5818),
		.dout(new_net_5819)
	);

	bfr new_net_5820_bfr_after (
		.din(new_net_5819),
		.dout(new_net_5820)
	);

	bfr new_net_5821_bfr_after (
		.din(new_net_5820),
		.dout(new_net_5821)
	);

	bfr new_net_5822_bfr_after (
		.din(new_net_5821),
		.dout(new_net_5822)
	);

	bfr new_net_5823_bfr_after (
		.din(new_net_5822),
		.dout(new_net_5823)
	);

	bfr new_net_5824_bfr_after (
		.din(new_net_5823),
		.dout(new_net_5824)
	);

	bfr new_net_5825_bfr_after (
		.din(new_net_5824),
		.dout(new_net_5825)
	);

	bfr new_net_2305_bfr_after (
		.din(new_net_5825),
		.dout(new_net_2305)
	);

	bfr new_net_5826_bfr_after (
		.din(G120),
		.dout(new_net_5826)
	);

	bfr new_net_5827_bfr_after (
		.din(new_net_5826),
		.dout(new_net_5827)
	);

	bfr new_net_2172_bfr_after (
		.din(new_net_5827),
		.dout(new_net_2172)
	);

	bfr new_net_5828_bfr_after (
		.din(new_net_2497),
		.dout(new_net_5828)
	);

	bfr new_net_5829_bfr_after (
		.din(new_net_5828),
		.dout(new_net_5829)
	);

	bfr new_net_5830_bfr_after (
		.din(new_net_5829),
		.dout(new_net_5830)
	);

	bfr new_net_5831_bfr_after (
		.din(new_net_5830),
		.dout(new_net_5831)
	);

	bfr new_net_5832_bfr_after (
		.din(new_net_5831),
		.dout(new_net_5832)
	);

	bfr new_net_5833_bfr_after (
		.din(new_net_5832),
		.dout(new_net_5833)
	);

	bfr new_net_5834_bfr_after (
		.din(new_net_5833),
		.dout(new_net_5834)
	);

	bfr new_net_5835_bfr_after (
		.din(new_net_5834),
		.dout(new_net_5835)
	);

	bfr new_net_5836_bfr_after (
		.din(new_net_5835),
		.dout(new_net_5836)
	);

	bfr new_net_5837_bfr_after (
		.din(new_net_5836),
		.dout(new_net_5837)
	);

	bfr new_net_5838_bfr_after (
		.din(new_net_5837),
		.dout(new_net_5838)
	);

	bfr new_net_5839_bfr_after (
		.din(new_net_5838),
		.dout(new_net_5839)
	);

	bfr new_net_5840_bfr_after (
		.din(new_net_5839),
		.dout(new_net_5840)
	);

	bfr new_net_5841_bfr_after (
		.din(new_net_5840),
		.dout(new_net_5841)
	);

	bfr new_net_5842_bfr_after (
		.din(new_net_5841),
		.dout(new_net_5842)
	);

	bfr new_net_5843_bfr_after (
		.din(new_net_5842),
		.dout(new_net_5843)
	);

	bfr new_net_5844_bfr_after (
		.din(new_net_5843),
		.dout(new_net_5844)
	);

	bfr new_net_5845_bfr_after (
		.din(new_net_5844),
		.dout(new_net_5845)
	);

	bfr new_net_5846_bfr_after (
		.din(new_net_5845),
		.dout(new_net_5846)
	);

	bfr new_net_5847_bfr_after (
		.din(new_net_5846),
		.dout(new_net_5847)
	);

	bfr new_net_5848_bfr_after (
		.din(new_net_5847),
		.dout(new_net_5848)
	);

	bfr new_net_5849_bfr_after (
		.din(new_net_5848),
		.dout(new_net_5849)
	);

	bfr new_net_5850_bfr_after (
		.din(new_net_5849),
		.dout(new_net_5850)
	);

	bfr new_net_5851_bfr_after (
		.din(new_net_5850),
		.dout(new_net_5851)
	);

	bfr new_net_5852_bfr_after (
		.din(new_net_5851),
		.dout(new_net_5852)
	);

	bfr new_net_5853_bfr_after (
		.din(new_net_5852),
		.dout(new_net_5853)
	);

	bfr new_net_5854_bfr_after (
		.din(new_net_5853),
		.dout(new_net_5854)
	);

	bfr new_net_5855_bfr_after (
		.din(new_net_5854),
		.dout(new_net_5855)
	);

	bfr new_net_5856_bfr_after (
		.din(new_net_5855),
		.dout(new_net_5856)
	);

	bfr new_net_5857_bfr_after (
		.din(new_net_5856),
		.dout(new_net_5857)
	);

	bfr new_net_5858_bfr_after (
		.din(new_net_5857),
		.dout(new_net_5858)
	);

	bfr new_net_5859_bfr_after (
		.din(new_net_5858),
		.dout(new_net_5859)
	);

	bfr new_net_5860_bfr_after (
		.din(new_net_5859),
		.dout(new_net_5860)
	);

	bfr G5247_bfr_after (
		.din(new_net_5860),
		.dout(G5247)
	);

	bfr new_net_5861_bfr_after (
		.din(new_net_2423),
		.dout(new_net_5861)
	);

	bfr new_net_5862_bfr_after (
		.din(new_net_5861),
		.dout(new_net_5862)
	);

	bfr new_net_5863_bfr_after (
		.din(new_net_5862),
		.dout(new_net_5863)
	);

	bfr new_net_5864_bfr_after (
		.din(new_net_5863),
		.dout(new_net_5864)
	);

	bfr new_net_5865_bfr_after (
		.din(new_net_5864),
		.dout(new_net_5865)
	);

	bfr new_net_5866_bfr_after (
		.din(new_net_5865),
		.dout(new_net_5866)
	);

	bfr new_net_5867_bfr_after (
		.din(new_net_5866),
		.dout(new_net_5867)
	);

	bfr new_net_5868_bfr_after (
		.din(new_net_5867),
		.dout(new_net_5868)
	);

	bfr new_net_5869_bfr_after (
		.din(new_net_5868),
		.dout(new_net_5869)
	);

	bfr new_net_5870_bfr_after (
		.din(new_net_5869),
		.dout(new_net_5870)
	);

	bfr new_net_5871_bfr_after (
		.din(new_net_5870),
		.dout(new_net_5871)
	);

	bfr new_net_5872_bfr_after (
		.din(new_net_5871),
		.dout(new_net_5872)
	);

	bfr new_net_5873_bfr_after (
		.din(new_net_5872),
		.dout(new_net_5873)
	);

	bfr new_net_5874_bfr_after (
		.din(new_net_5873),
		.dout(new_net_5874)
	);

	bfr new_net_5875_bfr_after (
		.din(new_net_5874),
		.dout(new_net_5875)
	);

	bfr new_net_5876_bfr_after (
		.din(new_net_5875),
		.dout(new_net_5876)
	);

	bfr new_net_5877_bfr_after (
		.din(new_net_5876),
		.dout(new_net_5877)
	);

	bfr new_net_5878_bfr_after (
		.din(new_net_5877),
		.dout(new_net_5878)
	);

	bfr new_net_5879_bfr_after (
		.din(new_net_5878),
		.dout(new_net_5879)
	);

	bfr new_net_5880_bfr_after (
		.din(new_net_5879),
		.dout(new_net_5880)
	);

	bfr G5289_bfr_after (
		.din(new_net_5880),
		.dout(G5289)
	);

	bfr new_net_5881_bfr_after (
		.din(_0232_),
		.dout(new_net_5881)
	);

	bfr new_net_2258_bfr_after (
		.din(new_net_5881),
		.dout(new_net_2258)
	);

	bfr new_net_2153_bfr_after (
		.din(_0783_),
		.dout(new_net_2153)
	);

	bfr new_net_5882_bfr_after (
		.din(_0887_),
		.dout(new_net_5882)
	);

	bfr new_net_5883_bfr_after (
		.din(new_net_5882),
		.dout(new_net_5883)
	);

	bfr new_net_5884_bfr_after (
		.din(new_net_5883),
		.dout(new_net_5884)
	);

	bfr new_net_5885_bfr_after (
		.din(new_net_5884),
		.dout(new_net_5885)
	);

	bfr new_net_5886_bfr_after (
		.din(new_net_5885),
		.dout(new_net_5886)
	);

	bfr new_net_5887_bfr_after (
		.din(new_net_5886),
		.dout(new_net_5887)
	);

	bfr new_net_5888_bfr_after (
		.din(new_net_5887),
		.dout(new_net_5888)
	);

	bfr new_net_5889_bfr_after (
		.din(new_net_5888),
		.dout(new_net_5889)
	);

	bfr new_net_5890_bfr_after (
		.din(new_net_5889),
		.dout(new_net_5890)
	);

	bfr new_net_5891_bfr_after (
		.din(new_net_5890),
		.dout(new_net_5891)
	);

	bfr new_net_5892_bfr_after (
		.din(new_net_5891),
		.dout(new_net_5892)
	);

	bfr new_net_5893_bfr_after (
		.din(new_net_5892),
		.dout(new_net_5893)
	);

	bfr new_net_5894_bfr_after (
		.din(new_net_5893),
		.dout(new_net_5894)
	);

	bfr new_net_5895_bfr_after (
		.din(new_net_5894),
		.dout(new_net_5895)
	);

	bfr new_net_5896_bfr_after (
		.din(new_net_5895),
		.dout(new_net_5896)
	);

	bfr new_net_5897_bfr_after (
		.din(new_net_5896),
		.dout(new_net_5897)
	);

	bfr new_net_5898_bfr_after (
		.din(new_net_5897),
		.dout(new_net_5898)
	);

	bfr new_net_5899_bfr_after (
		.din(new_net_5898),
		.dout(new_net_5899)
	);

	bfr new_net_5900_bfr_after (
		.din(new_net_5899),
		.dout(new_net_5900)
	);

	bfr new_net_5901_bfr_after (
		.din(new_net_5900),
		.dout(new_net_5901)
	);

	bfr new_net_5902_bfr_after (
		.din(new_net_5901),
		.dout(new_net_5902)
	);

	bfr new_net_5903_bfr_after (
		.din(new_net_5902),
		.dout(new_net_5903)
	);

	bfr new_net_2174_bfr_after (
		.din(new_net_5903),
		.dout(new_net_2174)
	);

	bfr new_net_5904_bfr_after (
		.din(G65),
		.dout(new_net_5904)
	);

	bfr new_net_5905_bfr_after (
		.din(new_net_5904),
		.dout(new_net_5905)
	);

	bfr new_net_5906_bfr_after (
		.din(new_net_5905),
		.dout(new_net_5906)
	);

	bfr new_net_2111_bfr_after (
		.din(new_net_5906),
		.dout(new_net_2111)
	);

	bfr new_net_5907_bfr_after (
		.din(_0634_),
		.dout(new_net_5907)
	);

	bfr new_net_5908_bfr_after (
		.din(new_net_5907),
		.dout(new_net_5908)
	);

	bfr new_net_5909_bfr_after (
		.din(new_net_5908),
		.dout(new_net_5909)
	);

	bfr new_net_5910_bfr_after (
		.din(new_net_5909),
		.dout(new_net_5910)
	);

	bfr new_net_5911_bfr_after (
		.din(new_net_5910),
		.dout(new_net_5911)
	);

	bfr new_net_5912_bfr_after (
		.din(new_net_5911),
		.dout(new_net_5912)
	);

	bfr new_net_5913_bfr_after (
		.din(new_net_5912),
		.dout(new_net_5913)
	);

	bfr new_net_5914_bfr_after (
		.din(new_net_5913),
		.dout(new_net_5914)
	);

	bfr new_net_5915_bfr_after (
		.din(new_net_5914),
		.dout(new_net_5915)
	);

	bfr new_net_2132_bfr_after (
		.din(new_net_5915),
		.dout(new_net_2132)
	);

	bfr new_net_5916_bfr_after (
		.din(_0989_),
		.dout(new_net_5916)
	);

	bfr new_net_5917_bfr_after (
		.din(new_net_5916),
		.dout(new_net_5917)
	);

	bfr new_net_5918_bfr_after (
		.din(new_net_5917),
		.dout(new_net_5918)
	);

	bfr new_net_5919_bfr_after (
		.din(new_net_5918),
		.dout(new_net_5919)
	);

	bfr new_net_5920_bfr_after (
		.din(new_net_5919),
		.dout(new_net_5920)
	);

	bfr new_net_5921_bfr_after (
		.din(new_net_5920),
		.dout(new_net_5921)
	);

	bfr new_net_5922_bfr_after (
		.din(new_net_5921),
		.dout(new_net_5922)
	);

	bfr new_net_5923_bfr_after (
		.din(new_net_5922),
		.dout(new_net_5923)
	);

	bfr new_net_5924_bfr_after (
		.din(new_net_5923),
		.dout(new_net_5924)
	);

	bfr new_net_5925_bfr_after (
		.din(new_net_5924),
		.dout(new_net_5925)
	);

	bfr new_net_5926_bfr_after (
		.din(new_net_5925),
		.dout(new_net_5926)
	);

	bfr new_net_5927_bfr_after (
		.din(new_net_5926),
		.dout(new_net_5927)
	);

	bfr new_net_5928_bfr_after (
		.din(new_net_5927),
		.dout(new_net_5928)
	);

	bfr new_net_5929_bfr_after (
		.din(new_net_5928),
		.dout(new_net_5929)
	);

	bfr new_net_5930_bfr_after (
		.din(new_net_5929),
		.dout(new_net_5930)
	);

	bfr new_net_5931_bfr_after (
		.din(new_net_5930),
		.dout(new_net_5931)
	);

	bfr new_net_5932_bfr_after (
		.din(new_net_5931),
		.dout(new_net_5932)
	);

	bfr new_net_5933_bfr_after (
		.din(new_net_5932),
		.dout(new_net_5933)
	);

	bfr new_net_5934_bfr_after (
		.din(new_net_5933),
		.dout(new_net_5934)
	);

	bfr new_net_5935_bfr_after (
		.din(new_net_5934),
		.dout(new_net_5935)
	);

	bfr new_net_5936_bfr_after (
		.din(new_net_5935),
		.dout(new_net_5936)
	);

	bfr new_net_5937_bfr_after (
		.din(new_net_5936),
		.dout(new_net_5937)
	);

	bfr new_net_5938_bfr_after (
		.din(new_net_5937),
		.dout(new_net_5938)
	);

	bfr new_net_5939_bfr_after (
		.din(new_net_5938),
		.dout(new_net_5939)
	);

	bfr new_net_5940_bfr_after (
		.din(new_net_5939),
		.dout(new_net_5940)
	);

	bfr new_net_2195_bfr_after (
		.din(new_net_5940),
		.dout(new_net_2195)
	);

	bfr new_net_5941_bfr_after (
		.din(_0299_),
		.dout(new_net_5941)
	);

	bfr new_net_5942_bfr_after (
		.din(new_net_5941),
		.dout(new_net_5942)
	);

	bfr new_net_5943_bfr_after (
		.din(new_net_5942),
		.dout(new_net_5943)
	);

	bfr new_net_5944_bfr_after (
		.din(new_net_5943),
		.dout(new_net_5944)
	);

	bfr new_net_5945_bfr_after (
		.din(new_net_5944),
		.dout(new_net_5945)
	);

	bfr new_net_5946_bfr_after (
		.din(new_net_5945),
		.dout(new_net_5946)
	);

	bfr new_net_5947_bfr_after (
		.din(new_net_5946),
		.dout(new_net_5947)
	);

	bfr new_net_5948_bfr_after (
		.din(new_net_5947),
		.dout(new_net_5948)
	);

	bfr new_net_5949_bfr_after (
		.din(new_net_5948),
		.dout(new_net_5949)
	);

	bfr new_net_5950_bfr_after (
		.din(new_net_5949),
		.dout(new_net_5950)
	);

	bfr new_net_5951_bfr_after (
		.din(new_net_5950),
		.dout(new_net_5951)
	);

	bfr new_net_5952_bfr_after (
		.din(new_net_5951),
		.dout(new_net_5952)
	);

	bfr new_net_5953_bfr_after (
		.din(new_net_5952),
		.dout(new_net_5953)
	);

	bfr new_net_5954_bfr_after (
		.din(new_net_5953),
		.dout(new_net_5954)
	);

	bfr new_net_2279_bfr_after (
		.din(new_net_5954),
		.dout(new_net_2279)
	);

	bfr new_net_5955_bfr_after (
		.din(_0562_),
		.dout(new_net_5955)
	);

	bfr new_net_5956_bfr_after (
		.din(new_net_5955),
		.dout(new_net_5956)
	);

	bfr new_net_5957_bfr_after (
		.din(new_net_5956),
		.dout(new_net_5957)
	);

	bfr new_net_5958_bfr_after (
		.din(new_net_5957),
		.dout(new_net_5958)
	);

	bfr new_net_5959_bfr_after (
		.din(new_net_5958),
		.dout(new_net_5959)
	);

	bfr new_net_5960_bfr_after (
		.din(new_net_5959),
		.dout(new_net_5960)
	);

	bfr new_net_5961_bfr_after (
		.din(new_net_5960),
		.dout(new_net_5961)
	);

	bfr new_net_5962_bfr_after (
		.din(new_net_5961),
		.dout(new_net_5962)
	);

	bfr new_net_5963_bfr_after (
		.din(new_net_5962),
		.dout(new_net_5963)
	);

	bfr new_net_5964_bfr_after (
		.din(new_net_5963),
		.dout(new_net_5964)
	);

	bfr new_net_5965_bfr_after (
		.din(new_net_5964),
		.dout(new_net_5965)
	);

	bfr new_net_5966_bfr_after (
		.din(new_net_5965),
		.dout(new_net_5966)
	);

	bfr new_net_5967_bfr_after (
		.din(new_net_5966),
		.dout(new_net_5967)
	);

	bfr new_net_5968_bfr_after (
		.din(new_net_5967),
		.dout(new_net_5968)
	);

	bfr new_net_5969_bfr_after (
		.din(new_net_5968),
		.dout(new_net_5969)
	);

	bfr new_net_5970_bfr_after (
		.din(new_net_5969),
		.dout(new_net_5970)
	);

	bfr new_net_5971_bfr_after (
		.din(new_net_5970),
		.dout(new_net_5971)
	);

	bfr new_net_5972_bfr_after (
		.din(new_net_5971),
		.dout(new_net_5972)
	);

	bfr new_net_5973_bfr_after (
		.din(new_net_5972),
		.dout(new_net_5973)
	);

	bfr new_net_5974_bfr_after (
		.din(new_net_5973),
		.dout(new_net_5974)
	);

	bfr new_net_5975_bfr_after (
		.din(new_net_5974),
		.dout(new_net_5975)
	);

	bfr new_net_5976_bfr_after (
		.din(new_net_5975),
		.dout(new_net_5976)
	);

	bfr new_net_5977_bfr_after (
		.din(new_net_5976),
		.dout(new_net_5977)
	);

	bfr new_net_5978_bfr_after (
		.din(new_net_5977),
		.dout(new_net_5978)
	);

	bfr new_net_2342_bfr_after (
		.din(new_net_5978),
		.dout(new_net_2342)
	);

	bfr new_net_5979_bfr_after (
		.din(_0469_),
		.dout(new_net_5979)
	);

	bfr new_net_5980_bfr_after (
		.din(new_net_5979),
		.dout(new_net_5980)
	);

	bfr new_net_5981_bfr_after (
		.din(new_net_5980),
		.dout(new_net_5981)
	);

	bfr new_net_5982_bfr_after (
		.din(new_net_5981),
		.dout(new_net_5982)
	);

	bfr new_net_5983_bfr_after (
		.din(new_net_5982),
		.dout(new_net_5983)
	);

	bfr new_net_5984_bfr_after (
		.din(new_net_5983),
		.dout(new_net_5984)
	);

	bfr new_net_5985_bfr_after (
		.din(new_net_5984),
		.dout(new_net_5985)
	);

	bfr new_net_5986_bfr_after (
		.din(new_net_5985),
		.dout(new_net_5986)
	);

	bfr new_net_5987_bfr_after (
		.din(new_net_5986),
		.dout(new_net_5987)
	);

	bfr new_net_5988_bfr_after (
		.din(new_net_5987),
		.dout(new_net_5988)
	);

	bfr new_net_5989_bfr_after (
		.din(new_net_5988),
		.dout(new_net_5989)
	);

	bfr new_net_5990_bfr_after (
		.din(new_net_5989),
		.dout(new_net_5990)
	);

	bfr new_net_5991_bfr_after (
		.din(new_net_5990),
		.dout(new_net_5991)
	);

	bfr new_net_5992_bfr_after (
		.din(new_net_5991),
		.dout(new_net_5992)
	);

	bfr new_net_5993_bfr_after (
		.din(new_net_5992),
		.dout(new_net_5993)
	);

	bfr new_net_5994_bfr_after (
		.din(new_net_5993),
		.dout(new_net_5994)
	);

	bfr new_net_5995_bfr_after (
		.din(new_net_5994),
		.dout(new_net_5995)
	);

	bfr new_net_5996_bfr_after (
		.din(new_net_5995),
		.dout(new_net_5996)
	);

	bfr new_net_5997_bfr_after (
		.din(new_net_5996),
		.dout(new_net_5997)
	);

	bfr new_net_5998_bfr_after (
		.din(new_net_5997),
		.dout(new_net_5998)
	);

	bfr new_net_5999_bfr_after (
		.din(new_net_5998),
		.dout(new_net_5999)
	);

	bfr new_net_6000_bfr_after (
		.din(new_net_5999),
		.dout(new_net_6000)
	);

	bfr new_net_6001_bfr_after (
		.din(new_net_6000),
		.dout(new_net_6001)
	);

	bfr new_net_6002_bfr_after (
		.din(new_net_6001),
		.dout(new_net_6002)
	);

	bfr new_net_6003_bfr_after (
		.din(new_net_6002),
		.dout(new_net_6003)
	);

	bfr new_net_6004_bfr_after (
		.din(new_net_6003),
		.dout(new_net_6004)
	);

	bfr new_net_6005_bfr_after (
		.din(new_net_6004),
		.dout(new_net_6005)
	);

	bfr new_net_6006_bfr_after (
		.din(new_net_6005),
		.dout(new_net_6006)
	);

	bfr new_net_6007_bfr_after (
		.din(new_net_6006),
		.dout(new_net_6007)
	);

	bfr new_net_6008_bfr_after (
		.din(new_net_6007),
		.dout(new_net_6008)
	);

	bfr new_net_6009_bfr_after (
		.din(new_net_6008),
		.dout(new_net_6009)
	);

	bfr new_net_2321_bfr_after (
		.din(new_net_6009),
		.dout(new_net_2321)
	);

	bfr new_net_2216_bfr_after (
		.din(G38),
		.dout(new_net_2216)
	);

	bfr new_net_6010_bfr_after (
		.din(G47),
		.dout(new_net_6010)
	);

	bfr new_net_6011_bfr_after (
		.din(new_net_6010),
		.dout(new_net_6011)
	);

	bfr new_net_6012_bfr_after (
		.din(new_net_6011),
		.dout(new_net_6012)
	);

	bfr new_net_6013_bfr_after (
		.din(new_net_6012),
		.dout(new_net_6013)
	);

	bfr new_net_2176_bfr_after (
		.din(new_net_6013),
		.dout(new_net_2176)
	);

	bfr new_net_6014_bfr_after (
		.din(G33),
		.dout(new_net_6014)
	);

	bfr new_net_2113_bfr_after (
		.din(new_net_6014),
		.dout(new_net_2113)
	);

	bfr new_net_6015_bfr_after (
		.din(_0089_),
		.dout(new_net_6015)
	);

	bfr new_net_6016_bfr_after (
		.din(new_net_6015),
		.dout(new_net_6016)
	);

	bfr new_net_2232_bfr_after (
		.din(new_net_6016),
		.dout(new_net_2232)
	);

	bfr new_net_6017_bfr_after (
		.din(_0224_),
		.dout(new_net_6017)
	);

	bfr new_net_2253_bfr_after (
		.din(new_net_6017),
		.dout(new_net_2253)
	);

	bfr new_net_6018_bfr_after (
		.din(_0451_),
		.dout(new_net_6018)
	);

	bfr new_net_6019_bfr_after (
		.din(new_net_6018),
		.dout(new_net_6019)
	);

	bfr new_net_6020_bfr_after (
		.din(new_net_6019),
		.dout(new_net_6020)
	);

	bfr new_net_6021_bfr_after (
		.din(new_net_6020),
		.dout(new_net_6021)
	);

	bfr new_net_6022_bfr_after (
		.din(new_net_6021),
		.dout(new_net_6022)
	);

	bfr new_net_6023_bfr_after (
		.din(new_net_6022),
		.dout(new_net_6023)
	);

	bfr new_net_6024_bfr_after (
		.din(new_net_6023),
		.dout(new_net_6024)
	);

	bfr new_net_6025_bfr_after (
		.din(new_net_6024),
		.dout(new_net_6025)
	);

	bfr new_net_6026_bfr_after (
		.din(new_net_6025),
		.dout(new_net_6026)
	);

	bfr new_net_6027_bfr_after (
		.din(new_net_6026),
		.dout(new_net_6027)
	);

	bfr new_net_6028_bfr_after (
		.din(new_net_6027),
		.dout(new_net_6028)
	);

	bfr new_net_6029_bfr_after (
		.din(new_net_6028),
		.dout(new_net_6029)
	);

	bfr new_net_6030_bfr_after (
		.din(new_net_6029),
		.dout(new_net_6030)
	);

	bfr new_net_6031_bfr_after (
		.din(new_net_6030),
		.dout(new_net_6031)
	);

	bfr new_net_6032_bfr_after (
		.din(new_net_6031),
		.dout(new_net_6032)
	);

	bfr new_net_6033_bfr_after (
		.din(new_net_6032),
		.dout(new_net_6033)
	);

	bfr new_net_2316_bfr_after (
		.din(new_net_6033),
		.dout(new_net_2316)
	);

	bfr new_net_6034_bfr_after (
		.din(_0282_),
		.dout(new_net_6034)
	);

	bfr new_net_6035_bfr_after (
		.din(new_net_6034),
		.dout(new_net_6035)
	);

	bfr new_net_2274_bfr_after (
		.din(new_net_6035),
		.dout(new_net_2274)
	);

	bfr new_net_6036_bfr_after (
		.din(_0546_),
		.dout(new_net_6036)
	);

	bfr new_net_2337_bfr_after (
		.din(new_net_6036),
		.dout(new_net_2337)
	);

	bfr new_net_6037_bfr_after (
		.din(new_net_2445),
		.dout(new_net_6037)
	);

	bfr new_net_6038_bfr_after (
		.din(new_net_6037),
		.dout(new_net_6038)
	);

	bfr new_net_6039_bfr_after (
		.din(new_net_6038),
		.dout(new_net_6039)
	);

	bfr new_net_6040_bfr_after (
		.din(new_net_6039),
		.dout(new_net_6040)
	);

	bfr new_net_6041_bfr_after (
		.din(new_net_6040),
		.dout(new_net_6041)
	);

	bfr new_net_6042_bfr_after (
		.din(new_net_6041),
		.dout(new_net_6042)
	);

	bfr new_net_6043_bfr_after (
		.din(new_net_6042),
		.dout(new_net_6043)
	);

	bfr new_net_6044_bfr_after (
		.din(new_net_6043),
		.dout(new_net_6044)
	);

	bfr new_net_6045_bfr_after (
		.din(new_net_6044),
		.dout(new_net_6045)
	);

	bfr G5279_bfr_after (
		.din(new_net_6045),
		.dout(G5279)
	);

	bfr new_net_6046_bfr_after (
		.din(new_net_2457),
		.dout(new_net_6046)
	);

	bfr new_net_6047_bfr_after (
		.din(new_net_6046),
		.dout(new_net_6047)
	);

	bfr G5297_bfr_after (
		.din(new_net_6047),
		.dout(G5297)
	);

	bfr new_net_6048_bfr_after (
		.din(G106),
		.dout(new_net_6048)
	);

	bfr new_net_2148_bfr_after (
		.din(new_net_6048),
		.dout(new_net_2148)
	);

	bfr new_net_6049_bfr_after (
		.din(_0850_),
		.dout(new_net_6049)
	);

	bfr new_net_6050_bfr_after (
		.din(new_net_6049),
		.dout(new_net_6050)
	);

	bfr new_net_6051_bfr_after (
		.din(new_net_6050),
		.dout(new_net_6051)
	);

	bfr new_net_6052_bfr_after (
		.din(new_net_6051),
		.dout(new_net_6052)
	);

	bfr new_net_6053_bfr_after (
		.din(new_net_6052),
		.dout(new_net_6053)
	);

	bfr new_net_6054_bfr_after (
		.din(new_net_6053),
		.dout(new_net_6054)
	);

	bfr new_net_6055_bfr_after (
		.din(new_net_6054),
		.dout(new_net_6055)
	);

	bfr new_net_2169_bfr_after (
		.din(new_net_6055),
		.dout(new_net_2169)
	);

	bfr new_net_6056_bfr_after (
		.din(G48),
		.dout(new_net_6056)
	);

	bfr new_net_6057_bfr_after (
		.din(new_net_6056),
		.dout(new_net_6057)
	);

	bfr new_net_6058_bfr_after (
		.din(new_net_6057),
		.dout(new_net_6058)
	);

	bfr new_net_6059_bfr_after (
		.din(new_net_6058),
		.dout(new_net_6059)
	);

	bfr new_net_2127_bfr_after (
		.din(new_net_6059),
		.dout(new_net_2127)
	);

	bfr new_net_6060_bfr_after (
		.din(new_net_2463),
		.dout(new_net_6060)
	);

	bfr new_net_6061_bfr_after (
		.din(new_net_6060),
		.dout(new_net_6061)
	);

	bfr new_net_6062_bfr_after (
		.din(new_net_6061),
		.dout(new_net_6062)
	);

	bfr new_net_6063_bfr_after (
		.din(new_net_6062),
		.dout(new_net_6063)
	);

	bfr new_net_6064_bfr_after (
		.din(new_net_6063),
		.dout(new_net_6064)
	);

	bfr new_net_6065_bfr_after (
		.din(new_net_6064),
		.dout(new_net_6065)
	);

	bfr new_net_6066_bfr_after (
		.din(new_net_6065),
		.dout(new_net_6066)
	);

	bfr new_net_6067_bfr_after (
		.din(new_net_6066),
		.dout(new_net_6067)
	);

	bfr new_net_6068_bfr_after (
		.din(new_net_6067),
		.dout(new_net_6068)
	);

	bfr new_net_6069_bfr_after (
		.din(new_net_6068),
		.dout(new_net_6069)
	);

	bfr new_net_6070_bfr_after (
		.din(new_net_6069),
		.dout(new_net_6070)
	);

	bfr new_net_6071_bfr_after (
		.din(new_net_6070),
		.dout(new_net_6071)
	);

	bfr new_net_6072_bfr_after (
		.din(new_net_6071),
		.dout(new_net_6072)
	);

	bfr new_net_6073_bfr_after (
		.din(new_net_6072),
		.dout(new_net_6073)
	);

	bfr new_net_6074_bfr_after (
		.din(new_net_6073),
		.dout(new_net_6074)
	);

	bfr new_net_6075_bfr_after (
		.din(new_net_6074),
		.dout(new_net_6075)
	);

	bfr new_net_6076_bfr_after (
		.din(new_net_6075),
		.dout(new_net_6076)
	);

	bfr new_net_6077_bfr_after (
		.din(new_net_6076),
		.dout(new_net_6077)
	);

	bfr new_net_6078_bfr_after (
		.din(new_net_6077),
		.dout(new_net_6078)
	);

	bfr new_net_6079_bfr_after (
		.din(new_net_6078),
		.dout(new_net_6079)
	);

	bfr new_net_6080_bfr_after (
		.din(new_net_6079),
		.dout(new_net_6080)
	);

	bfr new_net_6081_bfr_after (
		.din(new_net_6080),
		.dout(new_net_6081)
	);

	bfr new_net_6082_bfr_after (
		.din(new_net_6081),
		.dout(new_net_6082)
	);

	bfr new_net_6083_bfr_after (
		.din(new_net_6082),
		.dout(new_net_6083)
	);

	bfr new_net_6084_bfr_after (
		.din(new_net_6083),
		.dout(new_net_6084)
	);

	bfr new_net_6085_bfr_after (
		.din(new_net_6084),
		.dout(new_net_6085)
	);

	bfr new_net_6086_bfr_after (
		.din(new_net_6085),
		.dout(new_net_6086)
	);

	bfr new_net_6087_bfr_after (
		.din(new_net_6086),
		.dout(new_net_6087)
	);

	bfr new_net_6088_bfr_after (
		.din(new_net_6087),
		.dout(new_net_6088)
	);

	bfr new_net_6089_bfr_after (
		.din(new_net_6088),
		.dout(new_net_6089)
	);

	bfr new_net_6090_bfr_after (
		.din(new_net_6089),
		.dout(new_net_6090)
	);

	bfr new_net_6091_bfr_after (
		.din(new_net_6090),
		.dout(new_net_6091)
	);

	bfr new_net_6092_bfr_after (
		.din(new_net_6091),
		.dout(new_net_6092)
	);

	bfr new_net_6093_bfr_after (
		.din(new_net_6092),
		.dout(new_net_6093)
	);

	bfr new_net_6094_bfr_after (
		.din(new_net_6093),
		.dout(new_net_6094)
	);

	bfr new_net_6095_bfr_after (
		.din(new_net_6094),
		.dout(new_net_6095)
	);

	bfr new_net_6096_bfr_after (
		.din(new_net_6095),
		.dout(new_net_6096)
	);

	bfr new_net_6097_bfr_after (
		.din(new_net_6096),
		.dout(new_net_6097)
	);

	bfr new_net_6098_bfr_after (
		.din(new_net_6097),
		.dout(new_net_6098)
	);

	bfr G5198_bfr_after (
		.din(new_net_6098),
		.dout(G5198)
	);

	bfr new_net_6099_bfr_after (
		.din(new_net_2421),
		.dout(new_net_6099)
	);

	bfr new_net_6100_bfr_after (
		.din(new_net_6099),
		.dout(new_net_6100)
	);

	bfr new_net_6101_bfr_after (
		.din(new_net_6100),
		.dout(new_net_6101)
	);

	bfr new_net_6102_bfr_after (
		.din(new_net_6101),
		.dout(new_net_6102)
	);

	bfr new_net_6103_bfr_after (
		.din(new_net_6102),
		.dout(new_net_6103)
	);

	bfr new_net_6104_bfr_after (
		.din(new_net_6103),
		.dout(new_net_6104)
	);

	bfr new_net_6105_bfr_after (
		.din(new_net_6104),
		.dout(new_net_6105)
	);

	bfr new_net_6106_bfr_after (
		.din(new_net_6105),
		.dout(new_net_6106)
	);

	bfr new_net_6107_bfr_after (
		.din(new_net_6106),
		.dout(new_net_6107)
	);

	bfr new_net_6108_bfr_after (
		.din(new_net_6107),
		.dout(new_net_6108)
	);

	bfr new_net_6109_bfr_after (
		.din(new_net_6108),
		.dout(new_net_6109)
	);

	bfr new_net_6110_bfr_after (
		.din(new_net_6109),
		.dout(new_net_6110)
	);

	bfr new_net_6111_bfr_after (
		.din(new_net_6110),
		.dout(new_net_6111)
	);

	bfr new_net_6112_bfr_after (
		.din(new_net_6111),
		.dout(new_net_6112)
	);

	bfr new_net_6113_bfr_after (
		.din(new_net_6112),
		.dout(new_net_6113)
	);

	bfr new_net_6114_bfr_after (
		.din(new_net_6113),
		.dout(new_net_6114)
	);

	bfr new_net_6115_bfr_after (
		.din(new_net_6114),
		.dout(new_net_6115)
	);

	bfr new_net_6116_bfr_after (
		.din(new_net_6115),
		.dout(new_net_6116)
	);

	bfr new_net_6117_bfr_after (
		.din(new_net_6116),
		.dout(new_net_6117)
	);

	bfr new_net_6118_bfr_after (
		.din(new_net_6117),
		.dout(new_net_6118)
	);

	bfr new_net_6119_bfr_after (
		.din(new_net_6118),
		.dout(new_net_6119)
	);

	bfr G5241_bfr_after (
		.din(new_net_6119),
		.dout(G5241)
	);

	bfr new_net_6120_bfr_after (
		.din(new_net_2439),
		.dout(new_net_6120)
	);

	bfr new_net_6121_bfr_after (
		.din(new_net_6120),
		.dout(new_net_6121)
	);

	bfr new_net_6122_bfr_after (
		.din(new_net_6121),
		.dout(new_net_6122)
	);

	bfr G5294_bfr_after (
		.din(new_net_6122),
		.dout(G5294)
	);

	bfr new_net_6123_bfr_after (
		.din(new_net_2451),
		.dout(new_net_6123)
	);

	bfr new_net_6124_bfr_after (
		.din(new_net_6123),
		.dout(new_net_6124)
	);

	bfr new_net_6125_bfr_after (
		.din(new_net_6124),
		.dout(new_net_6125)
	);

	bfr new_net_6126_bfr_after (
		.din(new_net_6125),
		.dout(new_net_6126)
	);

	bfr new_net_6127_bfr_after (
		.din(new_net_6126),
		.dout(new_net_6127)
	);

	bfr new_net_6128_bfr_after (
		.din(new_net_6127),
		.dout(new_net_6128)
	);

	bfr new_net_6129_bfr_after (
		.din(new_net_6128),
		.dout(new_net_6129)
	);

	bfr new_net_6130_bfr_after (
		.din(new_net_6129),
		.dout(new_net_6130)
	);

	bfr new_net_6131_bfr_after (
		.din(new_net_6130),
		.dout(new_net_6131)
	);

	bfr new_net_6132_bfr_after (
		.din(new_net_6131),
		.dout(new_net_6132)
	);

	bfr new_net_6133_bfr_after (
		.din(new_net_6132),
		.dout(new_net_6133)
	);

	bfr new_net_6134_bfr_after (
		.din(new_net_6133),
		.dout(new_net_6134)
	);

	bfr new_net_6135_bfr_after (
		.din(new_net_6134),
		.dout(new_net_6135)
	);

	bfr new_net_6136_bfr_after (
		.din(new_net_6135),
		.dout(new_net_6136)
	);

	bfr new_net_6137_bfr_after (
		.din(new_net_6136),
		.dout(new_net_6137)
	);

	bfr new_net_6138_bfr_after (
		.din(new_net_6137),
		.dout(new_net_6138)
	);

	bfr new_net_6139_bfr_after (
		.din(new_net_6138),
		.dout(new_net_6139)
	);

	bfr new_net_6140_bfr_after (
		.din(new_net_6139),
		.dout(new_net_6140)
	);

	bfr new_net_6141_bfr_after (
		.din(new_net_6140),
		.dout(new_net_6141)
	);

	bfr G5256_bfr_after (
		.din(new_net_6141),
		.dout(G5256)
	);

	bfr new_net_6142_bfr_after (
		.din(new_net_2475),
		.dout(new_net_6142)
	);

	bfr new_net_6143_bfr_after (
		.din(new_net_6142),
		.dout(new_net_6143)
	);

	bfr new_net_6144_bfr_after (
		.din(new_net_6143),
		.dout(new_net_6144)
	);

	bfr new_net_6145_bfr_after (
		.din(new_net_6144),
		.dout(new_net_6145)
	);

	bfr new_net_6146_bfr_after (
		.din(new_net_6145),
		.dout(new_net_6146)
	);

	bfr new_net_6147_bfr_after (
		.din(new_net_6146),
		.dout(new_net_6147)
	);

	bfr new_net_6148_bfr_after (
		.din(new_net_6147),
		.dout(new_net_6148)
	);

	bfr new_net_6149_bfr_after (
		.din(new_net_6148),
		.dout(new_net_6149)
	);

	bfr new_net_6150_bfr_after (
		.din(new_net_6149),
		.dout(new_net_6150)
	);

	bfr new_net_6151_bfr_after (
		.din(new_net_6150),
		.dout(new_net_6151)
	);

	bfr new_net_6152_bfr_after (
		.din(new_net_6151),
		.dout(new_net_6152)
	);

	bfr new_net_6153_bfr_after (
		.din(new_net_6152),
		.dout(new_net_6153)
	);

	bfr new_net_6154_bfr_after (
		.din(new_net_6153),
		.dout(new_net_6154)
	);

	bfr new_net_6155_bfr_after (
		.din(new_net_6154),
		.dout(new_net_6155)
	);

	bfr G5280_bfr_after (
		.din(new_net_6155),
		.dout(G5280)
	);

	bfr new_net_6156_bfr_after (
		.din(new_net_2487),
		.dout(new_net_6156)
	);

	bfr new_net_6157_bfr_after (
		.din(new_net_6156),
		.dout(new_net_6157)
	);

	bfr new_net_6158_bfr_after (
		.din(new_net_6157),
		.dout(new_net_6158)
	);

	bfr new_net_6159_bfr_after (
		.din(new_net_6158),
		.dout(new_net_6159)
	);

	bfr new_net_6160_bfr_after (
		.din(new_net_6159),
		.dout(new_net_6160)
	);

	bfr new_net_6161_bfr_after (
		.din(new_net_6160),
		.dout(new_net_6161)
	);

	bfr new_net_6162_bfr_after (
		.din(new_net_6161),
		.dout(new_net_6162)
	);

	bfr new_net_6163_bfr_after (
		.din(new_net_6162),
		.dout(new_net_6163)
	);

	bfr new_net_6164_bfr_after (
		.din(new_net_6163),
		.dout(new_net_6164)
	);

	bfr new_net_6165_bfr_after (
		.din(new_net_6164),
		.dout(new_net_6165)
	);

	bfr new_net_6166_bfr_after (
		.din(new_net_6165),
		.dout(new_net_6166)
	);

	bfr new_net_6167_bfr_after (
		.din(new_net_6166),
		.dout(new_net_6167)
	);

	bfr new_net_6168_bfr_after (
		.din(new_net_6167),
		.dout(new_net_6168)
	);

	bfr new_net_6169_bfr_after (
		.din(new_net_6168),
		.dout(new_net_6169)
	);

	bfr new_net_6170_bfr_after (
		.din(new_net_6169),
		.dout(new_net_6170)
	);

	bfr new_net_6171_bfr_after (
		.din(new_net_6170),
		.dout(new_net_6171)
	);

	bfr new_net_6172_bfr_after (
		.din(new_net_6171),
		.dout(new_net_6172)
	);

	bfr new_net_6173_bfr_after (
		.din(new_net_6172),
		.dout(new_net_6173)
	);

	bfr new_net_6174_bfr_after (
		.din(new_net_6173),
		.dout(new_net_6174)
	);

	bfr new_net_6175_bfr_after (
		.din(new_net_6174),
		.dout(new_net_6175)
	);

	bfr new_net_6176_bfr_after (
		.din(new_net_6175),
		.dout(new_net_6176)
	);

	bfr new_net_6177_bfr_after (
		.din(new_net_6176),
		.dout(new_net_6177)
	);

	bfr new_net_6178_bfr_after (
		.din(new_net_6177),
		.dout(new_net_6178)
	);

	bfr new_net_6179_bfr_after (
		.din(new_net_6178),
		.dout(new_net_6179)
	);

	bfr new_net_6180_bfr_after (
		.din(new_net_6179),
		.dout(new_net_6180)
	);

	bfr new_net_6181_bfr_after (
		.din(new_net_6180),
		.dout(new_net_6181)
	);

	bfr new_net_6182_bfr_after (
		.din(new_net_6181),
		.dout(new_net_6182)
	);

	bfr new_net_6183_bfr_after (
		.din(new_net_6182),
		.dout(new_net_6183)
	);

	bfr new_net_6184_bfr_after (
		.din(new_net_6183),
		.dout(new_net_6184)
	);

	bfr new_net_6185_bfr_after (
		.din(new_net_6184),
		.dout(new_net_6185)
	);

	bfr new_net_6186_bfr_after (
		.din(new_net_6185),
		.dout(new_net_6186)
	);

	bfr new_net_6187_bfr_after (
		.din(new_net_6186),
		.dout(new_net_6187)
	);

	bfr new_net_6188_bfr_after (
		.din(new_net_6187),
		.dout(new_net_6188)
	);

	bfr new_net_6189_bfr_after (
		.din(new_net_6188),
		.dout(new_net_6189)
	);

	bfr new_net_6190_bfr_after (
		.din(new_net_6189),
		.dout(new_net_6190)
	);

	bfr new_net_6191_bfr_after (
		.din(new_net_6190),
		.dout(new_net_6191)
	);

	bfr new_net_6192_bfr_after (
		.din(new_net_6191),
		.dout(new_net_6192)
	);

	bfr new_net_6193_bfr_after (
		.din(new_net_6192),
		.dout(new_net_6193)
	);

	bfr G5194_bfr_after (
		.din(new_net_6193),
		.dout(G5194)
	);

	bfr new_net_6194_bfr_after (
		.din(new_net_2499),
		.dout(new_net_6194)
	);

	bfr new_net_6195_bfr_after (
		.din(new_net_6194),
		.dout(new_net_6195)
	);

	bfr new_net_6196_bfr_after (
		.din(new_net_6195),
		.dout(new_net_6196)
	);

	bfr new_net_6197_bfr_after (
		.din(new_net_6196),
		.dout(new_net_6197)
	);

	bfr new_net_6198_bfr_after (
		.din(new_net_6197),
		.dout(new_net_6198)
	);

	bfr new_net_6199_bfr_after (
		.din(new_net_6198),
		.dout(new_net_6199)
	);

	bfr new_net_6200_bfr_after (
		.din(new_net_6199),
		.dout(new_net_6200)
	);

	bfr new_net_6201_bfr_after (
		.din(new_net_6200),
		.dout(new_net_6201)
	);

	bfr new_net_6202_bfr_after (
		.din(new_net_6201),
		.dout(new_net_6202)
	);

	bfr new_net_6203_bfr_after (
		.din(new_net_6202),
		.dout(new_net_6203)
	);

	bfr new_net_6204_bfr_after (
		.din(new_net_6203),
		.dout(new_net_6204)
	);

	bfr new_net_6205_bfr_after (
		.din(new_net_6204),
		.dout(new_net_6205)
	);

	bfr new_net_6206_bfr_after (
		.din(new_net_6205),
		.dout(new_net_6206)
	);

	bfr new_net_6207_bfr_after (
		.din(new_net_6206),
		.dout(new_net_6207)
	);

	bfr new_net_6208_bfr_after (
		.din(new_net_6207),
		.dout(new_net_6208)
	);

	bfr new_net_6209_bfr_after (
		.din(new_net_6208),
		.dout(new_net_6209)
	);

	bfr new_net_6210_bfr_after (
		.din(new_net_6209),
		.dout(new_net_6210)
	);

	bfr new_net_6211_bfr_after (
		.din(new_net_6210),
		.dout(new_net_6211)
	);

	bfr new_net_6212_bfr_after (
		.din(new_net_6211),
		.dout(new_net_6212)
	);

	bfr new_net_6213_bfr_after (
		.din(new_net_6212),
		.dout(new_net_6213)
	);

	bfr new_net_6214_bfr_after (
		.din(new_net_6213),
		.dout(new_net_6214)
	);

	bfr new_net_6215_bfr_after (
		.din(new_net_6214),
		.dout(new_net_6215)
	);

	bfr new_net_6216_bfr_after (
		.din(new_net_6215),
		.dout(new_net_6216)
	);

	bfr new_net_6217_bfr_after (
		.din(new_net_6216),
		.dout(new_net_6217)
	);

	bfr new_net_6218_bfr_after (
		.din(new_net_6217),
		.dout(new_net_6218)
	);

	bfr new_net_6219_bfr_after (
		.din(new_net_6218),
		.dout(new_net_6219)
	);

	bfr new_net_6220_bfr_after (
		.din(new_net_6219),
		.dout(new_net_6220)
	);

	bfr new_net_6221_bfr_after (
		.din(new_net_6220),
		.dout(new_net_6221)
	);

	bfr new_net_6222_bfr_after (
		.din(new_net_6221),
		.dout(new_net_6222)
	);

	bfr G5237_bfr_after (
		.din(new_net_6222),
		.dout(G5237)
	);

	bfr new_net_6223_bfr_after (
		.din(new_net_2511),
		.dout(new_net_6223)
	);

	bfr new_net_6224_bfr_after (
		.din(new_net_6223),
		.dout(new_net_6224)
	);

	bfr new_net_6225_bfr_after (
		.din(new_net_6224),
		.dout(new_net_6225)
	);

	bfr new_net_6226_bfr_after (
		.din(new_net_6225),
		.dout(new_net_6226)
	);

	bfr new_net_6227_bfr_after (
		.din(new_net_6226),
		.dout(new_net_6227)
	);

	bfr new_net_6228_bfr_after (
		.din(new_net_6227),
		.dout(new_net_6228)
	);

	bfr G5301_bfr_after (
		.din(new_net_6228),
		.dout(G5301)
	);

	bfr new_net_6229_bfr_after (
		.din(new_net_2363),
		.dout(new_net_6229)
	);

	bfr G5308_bfr_after (
		.din(new_net_6229),
		.dout(G5308)
	);

	bfr new_net_6230_bfr_after (
		.din(_0387_),
		.dout(new_net_6230)
	);

	bfr new_net_6231_bfr_after (
		.din(new_net_6230),
		.dout(new_net_6231)
	);

	bfr new_net_6232_bfr_after (
		.din(new_net_6231),
		.dout(new_net_6232)
	);

	bfr new_net_6233_bfr_after (
		.din(new_net_6232),
		.dout(new_net_6233)
	);

	bfr new_net_6234_bfr_after (
		.din(new_net_6233),
		.dout(new_net_6234)
	);

	bfr new_net_6235_bfr_after (
		.din(new_net_6234),
		.dout(new_net_6235)
	);

	bfr new_net_6236_bfr_after (
		.din(new_net_6235),
		.dout(new_net_6236)
	);

	bfr new_net_6237_bfr_after (
		.din(new_net_6236),
		.dout(new_net_6237)
	);

	bfr new_net_6238_bfr_after (
		.din(new_net_6237),
		.dout(new_net_6238)
	);

	bfr new_net_6239_bfr_after (
		.din(new_net_6238),
		.dout(new_net_6239)
	);

	bfr new_net_6240_bfr_after (
		.din(new_net_6239),
		.dout(new_net_6240)
	);

	bfr new_net_6241_bfr_after (
		.din(new_net_6240),
		.dout(new_net_6241)
	);

	bfr new_net_6242_bfr_after (
		.din(new_net_6241),
		.dout(new_net_6242)
	);

	bfr new_net_6243_bfr_after (
		.din(new_net_6242),
		.dout(new_net_6243)
	);

	bfr new_net_6244_bfr_after (
		.din(new_net_6243),
		.dout(new_net_6244)
	);

	bfr new_net_6245_bfr_after (
		.din(new_net_6244),
		.dout(new_net_6245)
	);

	bfr new_net_6246_bfr_after (
		.din(new_net_6245),
		.dout(new_net_6246)
	);

	bfr new_net_6247_bfr_after (
		.din(new_net_6246),
		.dout(new_net_6247)
	);

	bfr new_net_6248_bfr_after (
		.din(new_net_6247),
		.dout(new_net_6248)
	);

	bfr new_net_6249_bfr_after (
		.din(new_net_6248),
		.dout(new_net_6249)
	);

	bfr new_net_6250_bfr_after (
		.din(new_net_6249),
		.dout(new_net_6250)
	);

	bfr new_net_6251_bfr_after (
		.din(new_net_6250),
		.dout(new_net_6251)
	);

	bfr new_net_2300_bfr_after (
		.din(new_net_6251),
		.dout(new_net_2300)
	);

	bfr new_net_6252_bfr_after (
		.din(_0367_),
		.dout(new_net_6252)
	);

	bfr new_net_2295_bfr_after (
		.din(new_net_6252),
		.dout(new_net_2295)
	);

	bfr new_net_6253_bfr_after (
		.din(new_net_2413),
		.dout(new_net_6253)
	);

	bfr new_net_6254_bfr_after (
		.din(new_net_6253),
		.dout(new_net_6254)
	);

	bfr new_net_6255_bfr_after (
		.din(new_net_6254),
		.dout(new_net_6255)
	);

	bfr new_net_6256_bfr_after (
		.din(new_net_6255),
		.dout(new_net_6256)
	);

	bfr new_net_6257_bfr_after (
		.din(new_net_6256),
		.dout(new_net_6257)
	);

	bfr new_net_6258_bfr_after (
		.din(new_net_6257),
		.dout(new_net_6258)
	);

	bfr new_net_6259_bfr_after (
		.din(new_net_6258),
		.dout(new_net_6259)
	);

	bfr new_net_6260_bfr_after (
		.din(new_net_6259),
		.dout(new_net_6260)
	);

	bfr new_net_6261_bfr_after (
		.din(new_net_6260),
		.dout(new_net_6261)
	);

	bfr new_net_6262_bfr_after (
		.din(new_net_6261),
		.dout(new_net_6262)
	);

	bfr G5277_bfr_after (
		.din(new_net_6262),
		.dout(G5277)
	);

	bfr new_net_6263_bfr_after (
		.din(_0176_),
		.dout(new_net_6263)
	);

	bfr new_net_2238_bfr_after (
		.din(new_net_6263),
		.dout(new_net_2238)
	);

	bfr new_net_6264_bfr_after (
		.din(_1062_),
		.dout(new_net_6264)
	);

	bfr new_net_2206_bfr_after (
		.din(new_net_6264),
		.dout(new_net_2206)
	);

	bfr new_net_2227_bfr_after (
		.din(_0075_),
		.dout(new_net_2227)
	);

	bfr new_net_2248_bfr_after (
		.din(_0221_),
		.dout(new_net_2248)
	);

	bfr new_net_6265_bfr_after (
		.din(_0433_),
		.dout(new_net_6265)
	);

	bfr new_net_6266_bfr_after (
		.din(new_net_6265),
		.dout(new_net_6266)
	);

	bfr new_net_6267_bfr_after (
		.din(new_net_6266),
		.dout(new_net_6267)
	);

	bfr new_net_6268_bfr_after (
		.din(new_net_6267),
		.dout(new_net_6268)
	);

	bfr new_net_2311_bfr_after (
		.din(new_net_6268),
		.dout(new_net_2311)
	);

	bfr new_net_6269_bfr_after (
		.din(new_net_2431),
		.dout(new_net_6269)
	);

	bfr new_net_6270_bfr_after (
		.din(new_net_6269),
		.dout(new_net_6270)
	);

	bfr new_net_6271_bfr_after (
		.din(new_net_6270),
		.dout(new_net_6271)
	);

	bfr new_net_6272_bfr_after (
		.din(new_net_6271),
		.dout(new_net_6272)
	);

	bfr new_net_6273_bfr_after (
		.din(new_net_6272),
		.dout(new_net_6273)
	);

	bfr new_net_6274_bfr_after (
		.din(new_net_6273),
		.dout(new_net_6274)
	);

	bfr new_net_6275_bfr_after (
		.din(new_net_6274),
		.dout(new_net_6275)
	);

	bfr new_net_6276_bfr_after (
		.din(new_net_6275),
		.dout(new_net_6276)
	);

	bfr new_net_6277_bfr_after (
		.din(new_net_6276),
		.dout(new_net_6277)
	);

	bfr new_net_6278_bfr_after (
		.din(new_net_6277),
		.dout(new_net_6278)
	);

	bfr G5281_bfr_after (
		.din(new_net_6278),
		.dout(G5281)
	);

	bfr new_net_6279_bfr_after (
		.din(_0275_),
		.dout(new_net_6279)
	);

	bfr new_net_2269_bfr_after (
		.din(new_net_6279),
		.dout(new_net_2269)
	);

	bfr new_net_6280_bfr_after (
		.din(_0520_),
		.dout(new_net_6280)
	);

	bfr new_net_6281_bfr_after (
		.din(new_net_6280),
		.dout(new_net_6281)
	);

	bfr new_net_6282_bfr_after (
		.din(new_net_6281),
		.dout(new_net_6282)
	);

	bfr new_net_6283_bfr_after (
		.din(new_net_6282),
		.dout(new_net_6283)
	);

	bfr new_net_6284_bfr_after (
		.din(new_net_6283),
		.dout(new_net_6284)
	);

	bfr new_net_6285_bfr_after (
		.din(new_net_6284),
		.dout(new_net_6285)
	);

	bfr new_net_6286_bfr_after (
		.din(new_net_6285),
		.dout(new_net_6286)
	);

	bfr new_net_6287_bfr_after (
		.din(new_net_6286),
		.dout(new_net_6287)
	);

	bfr new_net_6288_bfr_after (
		.din(new_net_6287),
		.dout(new_net_6288)
	);

	bfr new_net_6289_bfr_after (
		.din(new_net_6288),
		.dout(new_net_6289)
	);

	bfr new_net_6290_bfr_after (
		.din(new_net_6289),
		.dout(new_net_6290)
	);

	bfr new_net_6291_bfr_after (
		.din(new_net_6290),
		.dout(new_net_6291)
	);

	bfr new_net_6292_bfr_after (
		.din(new_net_6291),
		.dout(new_net_6292)
	);

	bfr new_net_6293_bfr_after (
		.din(new_net_6292),
		.dout(new_net_6293)
	);

	bfr new_net_6294_bfr_after (
		.din(new_net_6293),
		.dout(new_net_6294)
	);

	bfr new_net_6295_bfr_after (
		.din(new_net_6294),
		.dout(new_net_6295)
	);

	bfr new_net_6296_bfr_after (
		.din(new_net_6295),
		.dout(new_net_6296)
	);

	bfr new_net_6297_bfr_after (
		.din(new_net_6296),
		.dout(new_net_6297)
	);

	bfr new_net_6298_bfr_after (
		.din(new_net_6297),
		.dout(new_net_6298)
	);

	bfr new_net_6299_bfr_after (
		.din(new_net_6298),
		.dout(new_net_6299)
	);

	bfr new_net_6300_bfr_after (
		.din(new_net_6299),
		.dout(new_net_6300)
	);

	bfr new_net_6301_bfr_after (
		.din(new_net_6300),
		.dout(new_net_6301)
	);

	bfr new_net_6302_bfr_after (
		.din(new_net_6301),
		.dout(new_net_6302)
	);

	bfr new_net_6303_bfr_after (
		.din(new_net_6302),
		.dout(new_net_6303)
	);

	bfr new_net_6304_bfr_after (
		.din(new_net_6303),
		.dout(new_net_6304)
	);

	bfr new_net_6305_bfr_after (
		.din(new_net_6304),
		.dout(new_net_6305)
	);

	bfr new_net_6306_bfr_after (
		.din(new_net_6305),
		.dout(new_net_6306)
	);

	bfr new_net_6307_bfr_after (
		.din(new_net_6306),
		.dout(new_net_6307)
	);

	bfr new_net_6308_bfr_after (
		.din(new_net_6307),
		.dout(new_net_6308)
	);

	bfr new_net_6309_bfr_after (
		.din(new_net_6308),
		.dout(new_net_6309)
	);

	bfr new_net_6310_bfr_after (
		.din(new_net_6309),
		.dout(new_net_6310)
	);

	bfr new_net_2332_bfr_after (
		.din(new_net_6310),
		.dout(new_net_2332)
	);

	bfr new_net_6311_bfr_after (
		.din(G58),
		.dout(new_net_6311)
	);

	bfr new_net_6312_bfr_after (
		.din(new_net_6311),
		.dout(new_net_6312)
	);

	bfr new_net_6313_bfr_after (
		.din(new_net_6312),
		.dout(new_net_6313)
	);

	bfr new_net_6314_bfr_after (
		.din(new_net_6313),
		.dout(new_net_6314)
	);

	bfr new_net_2122_bfr_after (
		.din(new_net_6314),
		.dout(new_net_2122)
	);

	bfr new_net_6315_bfr_after (
		.din(_0714_),
		.dout(new_net_6315)
	);

	bfr new_net_6316_bfr_after (
		.din(new_net_6315),
		.dout(new_net_6316)
	);

	bfr new_net_6317_bfr_after (
		.din(new_net_6316),
		.dout(new_net_6317)
	);

	bfr new_net_6318_bfr_after (
		.din(new_net_6317),
		.dout(new_net_6318)
	);

	bfr new_net_6319_bfr_after (
		.din(new_net_6318),
		.dout(new_net_6319)
	);

	bfr new_net_6320_bfr_after (
		.din(new_net_6319),
		.dout(new_net_6320)
	);

	bfr new_net_6321_bfr_after (
		.din(new_net_6320),
		.dout(new_net_6321)
	);

	bfr new_net_6322_bfr_after (
		.din(new_net_6321),
		.dout(new_net_6322)
	);

	bfr new_net_6323_bfr_after (
		.din(new_net_6322),
		.dout(new_net_6323)
	);

	bfr new_net_6324_bfr_after (
		.din(new_net_6323),
		.dout(new_net_6324)
	);

	bfr new_net_6325_bfr_after (
		.din(new_net_6324),
		.dout(new_net_6325)
	);

	bfr new_net_6326_bfr_after (
		.din(new_net_6325),
		.dout(new_net_6326)
	);

	bfr new_net_6327_bfr_after (
		.din(new_net_6326),
		.dout(new_net_6327)
	);

	bfr new_net_2143_bfr_after (
		.din(new_net_6327),
		.dout(new_net_2143)
	);

	bfr new_net_6328_bfr_after (
		.din(G55),
		.dout(new_net_6328)
	);

	bfr new_net_6329_bfr_after (
		.din(new_net_6328),
		.dout(new_net_6329)
	);

	bfr new_net_6330_bfr_after (
		.din(new_net_6329),
		.dout(new_net_6330)
	);

	bfr new_net_6331_bfr_after (
		.din(new_net_6330),
		.dout(new_net_6331)
	);

	bfr new_net_2164_bfr_after (
		.din(new_net_6331),
		.dout(new_net_2164)
	);

	bfr new_net_6332_bfr_after (
		.din(new_net_2419),
		.dout(new_net_6332)
	);

	bfr new_net_6333_bfr_after (
		.din(new_net_6332),
		.dout(new_net_6333)
	);

	bfr new_net_6334_bfr_after (
		.din(new_net_6333),
		.dout(new_net_6334)
	);

	bfr new_net_6335_bfr_after (
		.din(new_net_6334),
		.dout(new_net_6335)
	);

	bfr new_net_6336_bfr_after (
		.din(new_net_6335),
		.dout(new_net_6336)
	);

	bfr new_net_6337_bfr_after (
		.din(new_net_6336),
		.dout(new_net_6337)
	);

	bfr new_net_6338_bfr_after (
		.din(new_net_6337),
		.dout(new_net_6338)
	);

	bfr new_net_6339_bfr_after (
		.din(new_net_6338),
		.dout(new_net_6339)
	);

	bfr new_net_6340_bfr_after (
		.din(new_net_6339),
		.dout(new_net_6340)
	);

	bfr new_net_6341_bfr_after (
		.din(new_net_6340),
		.dout(new_net_6341)
	);

	bfr new_net_6342_bfr_after (
		.din(new_net_6341),
		.dout(new_net_6342)
	);

	bfr new_net_6343_bfr_after (
		.din(new_net_6342),
		.dout(new_net_6343)
	);

	bfr new_net_6344_bfr_after (
		.din(new_net_6343),
		.dout(new_net_6344)
	);

	bfr new_net_6345_bfr_after (
		.din(new_net_6344),
		.dout(new_net_6345)
	);

	bfr new_net_6346_bfr_after (
		.din(new_net_6345),
		.dout(new_net_6346)
	);

	bfr new_net_6347_bfr_after (
		.din(new_net_6346),
		.dout(new_net_6347)
	);

	bfr new_net_6348_bfr_after (
		.din(new_net_6347),
		.dout(new_net_6348)
	);

	bfr new_net_6349_bfr_after (
		.din(new_net_6348),
		.dout(new_net_6349)
	);

	bfr new_net_6350_bfr_after (
		.din(new_net_6349),
		.dout(new_net_6350)
	);

	bfr new_net_6351_bfr_after (
		.din(new_net_6350),
		.dout(new_net_6351)
	);

	bfr new_net_6352_bfr_after (
		.din(new_net_6351),
		.dout(new_net_6352)
	);

	bfr new_net_6353_bfr_after (
		.din(new_net_6352),
		.dout(new_net_6353)
	);

	bfr new_net_6354_bfr_after (
		.din(new_net_6353),
		.dout(new_net_6354)
	);

	bfr new_net_6355_bfr_after (
		.din(new_net_6354),
		.dout(new_net_6355)
	);

	bfr new_net_6356_bfr_after (
		.din(new_net_6355),
		.dout(new_net_6356)
	);

	bfr new_net_6357_bfr_after (
		.din(new_net_6356),
		.dout(new_net_6357)
	);

	bfr new_net_6358_bfr_after (
		.din(new_net_6357),
		.dout(new_net_6358)
	);

	bfr new_net_6359_bfr_after (
		.din(new_net_6358),
		.dout(new_net_6359)
	);

	bfr new_net_6360_bfr_after (
		.din(new_net_6359),
		.dout(new_net_6360)
	);

	bfr new_net_6361_bfr_after (
		.din(new_net_6360),
		.dout(new_net_6361)
	);

	bfr new_net_6362_bfr_after (
		.din(new_net_6361),
		.dout(new_net_6362)
	);

	bfr new_net_6363_bfr_after (
		.din(new_net_6362),
		.dout(new_net_6363)
	);

	bfr new_net_6364_bfr_after (
		.din(new_net_6363),
		.dout(new_net_6364)
	);

	bfr new_net_6365_bfr_after (
		.din(new_net_6364),
		.dout(new_net_6365)
	);

	bfr new_net_6366_bfr_after (
		.din(new_net_6365),
		.dout(new_net_6366)
	);

	bfr new_net_6367_bfr_after (
		.din(new_net_6366),
		.dout(new_net_6367)
	);

	bfr new_net_6368_bfr_after (
		.din(new_net_6367),
		.dout(new_net_6368)
	);

	bfr new_net_6369_bfr_after (
		.din(new_net_6368),
		.dout(new_net_6369)
	);

	bfr new_net_6370_bfr_after (
		.din(new_net_6369),
		.dout(new_net_6370)
	);

	bfr G5208_bfr_after (
		.din(new_net_6370),
		.dout(G5208)
	);

	bfr new_net_6371_bfr_after (
		.din(new_net_2509),
		.dout(new_net_6371)
	);

	bfr new_net_6372_bfr_after (
		.din(new_net_6371),
		.dout(new_net_6372)
	);

	bfr new_net_6373_bfr_after (
		.din(new_net_6372),
		.dout(new_net_6373)
	);

	bfr new_net_6374_bfr_after (
		.din(new_net_6373),
		.dout(new_net_6374)
	);

	bfr new_net_6375_bfr_after (
		.din(new_net_6374),
		.dout(new_net_6375)
	);

	bfr new_net_6376_bfr_after (
		.din(new_net_6375),
		.dout(new_net_6376)
	);

	bfr new_net_6377_bfr_after (
		.din(new_net_6376),
		.dout(new_net_6377)
	);

	bfr new_net_6378_bfr_after (
		.din(new_net_6377),
		.dout(new_net_6378)
	);

	bfr new_net_6379_bfr_after (
		.din(new_net_6378),
		.dout(new_net_6379)
	);

	bfr new_net_6380_bfr_after (
		.din(new_net_6379),
		.dout(new_net_6380)
	);

	bfr new_net_6381_bfr_after (
		.din(new_net_6380),
		.dout(new_net_6381)
	);

	bfr new_net_6382_bfr_after (
		.din(new_net_6381),
		.dout(new_net_6382)
	);

	bfr new_net_6383_bfr_after (
		.din(new_net_6382),
		.dout(new_net_6383)
	);

	bfr new_net_6384_bfr_after (
		.din(new_net_6383),
		.dout(new_net_6384)
	);

	bfr new_net_6385_bfr_after (
		.din(new_net_6384),
		.dout(new_net_6385)
	);

	bfr new_net_6386_bfr_after (
		.din(new_net_6385),
		.dout(new_net_6386)
	);

	bfr new_net_6387_bfr_after (
		.din(new_net_6386),
		.dout(new_net_6387)
	);

	bfr new_net_6388_bfr_after (
		.din(new_net_6387),
		.dout(new_net_6388)
	);

	bfr new_net_6389_bfr_after (
		.din(new_net_6388),
		.dout(new_net_6389)
	);

	bfr G5252_bfr_after (
		.din(new_net_6389),
		.dout(G5252)
	);

	bfr new_net_6390_bfr_after (
		.din(_0514_),
		.dout(new_net_6390)
	);

	bfr new_net_2331_bfr_after (
		.din(new_net_6390),
		.dout(new_net_2331)
	);

	bfr new_net_6391_bfr_after (
		.din(_0497_),
		.dout(new_net_6391)
	);

	bfr new_net_6392_bfr_after (
		.din(new_net_6391),
		.dout(new_net_6392)
	);

	bfr new_net_6393_bfr_after (
		.din(new_net_6392),
		.dout(new_net_6393)
	);

	bfr new_net_6394_bfr_after (
		.din(new_net_6393),
		.dout(new_net_6394)
	);

	bfr new_net_6395_bfr_after (
		.din(new_net_6394),
		.dout(new_net_6395)
	);

	bfr new_net_6396_bfr_after (
		.din(new_net_6395),
		.dout(new_net_6396)
	);

	bfr new_net_6397_bfr_after (
		.din(new_net_6396),
		.dout(new_net_6397)
	);

	bfr new_net_6398_bfr_after (
		.din(new_net_6397),
		.dout(new_net_6398)
	);

	bfr new_net_6399_bfr_after (
		.din(new_net_6398),
		.dout(new_net_6399)
	);

	bfr new_net_6400_bfr_after (
		.din(new_net_6399),
		.dout(new_net_6400)
	);

	bfr new_net_6401_bfr_after (
		.din(new_net_6400),
		.dout(new_net_6401)
	);

	bfr new_net_6402_bfr_after (
		.din(new_net_6401),
		.dout(new_net_6402)
	);

	bfr new_net_6403_bfr_after (
		.din(new_net_6402),
		.dout(new_net_6403)
	);

	bfr new_net_6404_bfr_after (
		.din(new_net_6403),
		.dout(new_net_6404)
	);

	bfr new_net_6405_bfr_after (
		.din(new_net_6404),
		.dout(new_net_6405)
	);

	bfr new_net_6406_bfr_after (
		.din(new_net_6405),
		.dout(new_net_6406)
	);

	bfr new_net_6407_bfr_after (
		.din(new_net_6406),
		.dout(new_net_6407)
	);

	bfr new_net_6408_bfr_after (
		.din(new_net_6407),
		.dout(new_net_6408)
	);

	bfr new_net_6409_bfr_after (
		.din(new_net_6408),
		.dout(new_net_6409)
	);

	bfr new_net_6410_bfr_after (
		.din(new_net_6409),
		.dout(new_net_6410)
	);

	bfr new_net_6411_bfr_after (
		.din(new_net_6410),
		.dout(new_net_6411)
	);

	bfr new_net_6412_bfr_after (
		.din(new_net_6411),
		.dout(new_net_6412)
	);

	bfr new_net_6413_bfr_after (
		.din(new_net_6412),
		.dout(new_net_6413)
	);

	bfr new_net_6414_bfr_after (
		.din(new_net_6413),
		.dout(new_net_6414)
	);

	bfr new_net_6415_bfr_after (
		.din(new_net_6414),
		.dout(new_net_6415)
	);

	bfr new_net_6416_bfr_after (
		.din(new_net_6415),
		.dout(new_net_6416)
	);

	bfr new_net_6417_bfr_after (
		.din(new_net_6416),
		.dout(new_net_6417)
	);

	bfr new_net_2326_bfr_after (
		.din(new_net_6417),
		.dout(new_net_2326)
	);

	bfr new_net_6418_bfr_after (
		.din(new_net_2407),
		.dout(new_net_6418)
	);

	bfr new_net_6419_bfr_after (
		.din(new_net_6418),
		.dout(new_net_6419)
	);

	bfr new_net_6420_bfr_after (
		.din(new_net_6419),
		.dout(new_net_6420)
	);

	bfr new_net_6421_bfr_after (
		.din(new_net_6420),
		.dout(new_net_6421)
	);

	bfr new_net_6422_bfr_after (
		.din(new_net_6421),
		.dout(new_net_6422)
	);

	bfr new_net_6423_bfr_after (
		.din(new_net_6422),
		.dout(new_net_6423)
	);

	bfr new_net_6424_bfr_after (
		.din(new_net_6423),
		.dout(new_net_6424)
	);

	bfr new_net_6425_bfr_after (
		.din(new_net_6424),
		.dout(new_net_6425)
	);

	bfr new_net_6426_bfr_after (
		.din(new_net_6425),
		.dout(new_net_6426)
	);

	bfr new_net_6427_bfr_after (
		.din(new_net_6426),
		.dout(new_net_6427)
	);

	bfr new_net_6428_bfr_after (
		.din(new_net_6427),
		.dout(new_net_6428)
	);

	bfr new_net_6429_bfr_after (
		.din(new_net_6428),
		.dout(new_net_6429)
	);

	bfr new_net_6430_bfr_after (
		.din(new_net_6429),
		.dout(new_net_6430)
	);

	bfr new_net_6431_bfr_after (
		.din(new_net_6430),
		.dout(new_net_6431)
	);

	bfr G5276_bfr_after (
		.din(new_net_6431),
		.dout(G5276)
	);

	bfr new_net_2207_bfr_after (
		.din(_1075_),
		.dout(new_net_2207)
	);

	bfr new_net_2202_bfr_after (
		.din(_1049_),
		.dout(new_net_2202)
	);

	bfr new_net_6432_bfr_after (
		.din(_0324_),
		.dout(new_net_6432)
	);

	bfr new_net_2285_bfr_after (
		.din(new_net_6432),
		.dout(new_net_2285)
	);

	bfr new_net_6433_bfr_after (
		.din(_0577_),
		.dout(new_net_6433)
	);

	bfr new_net_6434_bfr_after (
		.din(new_net_6433),
		.dout(new_net_6434)
	);

	bfr new_net_6435_bfr_after (
		.din(new_net_6434),
		.dout(new_net_6435)
	);

	bfr new_net_6436_bfr_after (
		.din(new_net_6435),
		.dout(new_net_6436)
	);

	bfr new_net_6437_bfr_after (
		.din(new_net_6436),
		.dout(new_net_6437)
	);

	bfr new_net_6438_bfr_after (
		.din(new_net_6437),
		.dout(new_net_6438)
	);

	bfr new_net_6439_bfr_after (
		.din(new_net_6438),
		.dout(new_net_6439)
	);

	bfr new_net_6440_bfr_after (
		.din(new_net_6439),
		.dout(new_net_6440)
	);

	bfr new_net_6441_bfr_after (
		.din(new_net_6440),
		.dout(new_net_6441)
	);

	bfr new_net_6442_bfr_after (
		.din(new_net_6441),
		.dout(new_net_6442)
	);

	bfr new_net_6443_bfr_after (
		.din(new_net_6442),
		.dout(new_net_6443)
	);

	bfr new_net_6444_bfr_after (
		.din(new_net_6443),
		.dout(new_net_6444)
	);

	bfr new_net_6445_bfr_after (
		.din(new_net_6444),
		.dout(new_net_6445)
	);

	bfr new_net_6446_bfr_after (
		.din(new_net_6445),
		.dout(new_net_6446)
	);

	bfr new_net_6447_bfr_after (
		.din(new_net_6446),
		.dout(new_net_6447)
	);

	bfr new_net_6448_bfr_after (
		.din(new_net_6447),
		.dout(new_net_6448)
	);

	bfr new_net_6449_bfr_after (
		.din(new_net_6448),
		.dout(new_net_6449)
	);

	bfr new_net_6450_bfr_after (
		.din(new_net_6449),
		.dout(new_net_6450)
	);

	bfr new_net_6451_bfr_after (
		.din(new_net_6450),
		.dout(new_net_6451)
	);

	bfr new_net_6452_bfr_after (
		.din(new_net_6451),
		.dout(new_net_6452)
	);

	bfr new_net_6453_bfr_after (
		.din(new_net_6452),
		.dout(new_net_6453)
	);

	bfr new_net_6454_bfr_after (
		.din(new_net_6453),
		.dout(new_net_6454)
	);

	bfr new_net_6455_bfr_after (
		.din(new_net_6454),
		.dout(new_net_6455)
	);

	bfr new_net_6456_bfr_after (
		.din(new_net_6455),
		.dout(new_net_6456)
	);

	bfr new_net_6457_bfr_after (
		.din(new_net_6456),
		.dout(new_net_6457)
	);

	bfr new_net_6458_bfr_after (
		.din(new_net_6457),
		.dout(new_net_6458)
	);

	bfr new_net_6459_bfr_after (
		.din(new_net_6458),
		.dout(new_net_6459)
	);

	bfr new_net_6460_bfr_after (
		.din(new_net_6459),
		.dout(new_net_6460)
	);

	bfr new_net_6461_bfr_after (
		.din(new_net_6460),
		.dout(new_net_6461)
	);

	bfr new_net_6462_bfr_after (
		.din(new_net_6461),
		.dout(new_net_6462)
	);

	bfr new_net_6463_bfr_after (
		.din(new_net_6462),
		.dout(new_net_6463)
	);

	bfr new_net_6464_bfr_after (
		.din(new_net_6463),
		.dout(new_net_6464)
	);

	bfr new_net_2348_bfr_after (
		.din(new_net_6464),
		.dout(new_net_2348)
	);

	bfr new_net_6465_bfr_after (
		.din(new_net_2371),
		.dout(new_net_6465)
	);

	bfr new_net_6466_bfr_after (
		.din(new_net_6465),
		.dout(new_net_6466)
	);

	bfr new_net_6467_bfr_after (
		.din(new_net_6466),
		.dout(new_net_6467)
	);

	bfr new_net_6468_bfr_after (
		.din(new_net_6467),
		.dout(new_net_6468)
	);

	bfr new_net_6469_bfr_after (
		.din(new_net_6468),
		.dout(new_net_6469)
	);

	bfr new_net_6470_bfr_after (
		.din(new_net_6469),
		.dout(new_net_6470)
	);

	bfr new_net_6471_bfr_after (
		.din(new_net_6470),
		.dout(new_net_6471)
	);

	bfr new_net_6472_bfr_after (
		.din(new_net_6471),
		.dout(new_net_6472)
	);

	bfr new_net_6473_bfr_after (
		.din(new_net_6472),
		.dout(new_net_6473)
	);

	bfr new_net_6474_bfr_after (
		.din(new_net_6473),
		.dout(new_net_6474)
	);

	bfr new_net_6475_bfr_after (
		.din(new_net_6474),
		.dout(new_net_6475)
	);

	bfr new_net_6476_bfr_after (
		.din(new_net_6475),
		.dout(new_net_6476)
	);

	bfr new_net_6477_bfr_after (
		.din(new_net_6476),
		.dout(new_net_6477)
	);

	bfr new_net_6478_bfr_after (
		.din(new_net_6477),
		.dout(new_net_6478)
	);

	bfr new_net_6479_bfr_after (
		.din(new_net_6478),
		.dout(new_net_6479)
	);

	bfr new_net_6480_bfr_after (
		.din(new_net_6479),
		.dout(new_net_6480)
	);

	bfr new_net_6481_bfr_after (
		.din(new_net_6480),
		.dout(new_net_6481)
	);

	bfr new_net_6482_bfr_after (
		.din(new_net_6481),
		.dout(new_net_6482)
	);

	bfr new_net_6483_bfr_after (
		.din(new_net_6482),
		.dout(new_net_6483)
	);

	bfr new_net_6484_bfr_after (
		.din(new_net_6483),
		.dout(new_net_6484)
	);

	bfr new_net_6485_bfr_after (
		.din(new_net_6484),
		.dout(new_net_6485)
	);

	bfr G5238_bfr_after (
		.din(new_net_6485),
		.dout(G5238)
	);

	bfr new_net_2222_bfr_after (
		.din(_0008_),
		.dout(new_net_2222)
	);

	bfr new_net_2306_bfr_after (
		.din(_0415_),
		.dout(new_net_2306)
	);

	bfr new_net_6486_bfr_after (
		.din(new_net_2395),
		.dout(new_net_6486)
	);

	bfr G5304_bfr_after (
		.din(new_net_6486),
		.dout(G5304)
	);

	bfr new_net_6487_bfr_after (
		.din(G8),
		.dout(new_net_6487)
	);

	bfr new_net_2243_bfr_after (
		.din(new_net_6487),
		.dout(new_net_2243)
	);

	bfr new_net_6488_bfr_after (
		.din(_0498_),
		.dout(new_net_6488)
	);

	bfr new_net_2327_bfr_after (
		.din(new_net_6488),
		.dout(new_net_2327)
	);

	bfr new_net_6489_bfr_after (
		.din(new_net_2383),
		.dout(new_net_6489)
	);

	bfr new_net_6490_bfr_after (
		.din(new_net_6489),
		.dout(new_net_6490)
	);

	bfr new_net_6491_bfr_after (
		.din(new_net_6490),
		.dout(new_net_6491)
	);

	bfr new_net_6492_bfr_after (
		.din(new_net_6491),
		.dout(new_net_6492)
	);

	bfr new_net_6493_bfr_after (
		.din(new_net_6492),
		.dout(new_net_6493)
	);

	bfr new_net_6494_bfr_after (
		.din(new_net_6493),
		.dout(new_net_6494)
	);

	bfr new_net_6495_bfr_after (
		.din(new_net_6494),
		.dout(new_net_6495)
	);

	bfr new_net_6496_bfr_after (
		.din(new_net_6495),
		.dout(new_net_6496)
	);

	bfr new_net_6497_bfr_after (
		.din(new_net_6496),
		.dout(new_net_6497)
	);

	bfr new_net_6498_bfr_after (
		.din(new_net_6497),
		.dout(new_net_6498)
	);

	bfr new_net_6499_bfr_after (
		.din(new_net_6498),
		.dout(new_net_6499)
	);

	bfr G5269_bfr_after (
		.din(new_net_6499),
		.dout(G5269)
	);

	bfr new_net_6500_bfr_after (
		.din(_0260_),
		.dout(new_net_6500)
	);

	bfr new_net_6501_bfr_after (
		.din(new_net_6500),
		.dout(new_net_6501)
	);

	bfr new_net_6502_bfr_after (
		.din(new_net_6501),
		.dout(new_net_6502)
	);

	bfr new_net_6503_bfr_after (
		.din(new_net_6502),
		.dout(new_net_6503)
	);

	bfr new_net_6504_bfr_after (
		.din(new_net_6503),
		.dout(new_net_6504)
	);

	bfr new_net_6505_bfr_after (
		.din(new_net_6504),
		.dout(new_net_6505)
	);

	bfr new_net_6506_bfr_after (
		.din(new_net_6505),
		.dout(new_net_6506)
	);

	bfr new_net_6507_bfr_after (
		.din(new_net_6506),
		.dout(new_net_6507)
	);

	bfr new_net_6508_bfr_after (
		.din(new_net_6507),
		.dout(new_net_6508)
	);

	bfr new_net_6509_bfr_after (
		.din(new_net_6508),
		.dout(new_net_6509)
	);

	bfr new_net_6510_bfr_after (
		.din(new_net_6509),
		.dout(new_net_6510)
	);

	bfr new_net_6511_bfr_after (
		.din(new_net_6510),
		.dout(new_net_6511)
	);

	bfr new_net_6512_bfr_after (
		.din(new_net_6511),
		.dout(new_net_6512)
	);

	bfr new_net_6513_bfr_after (
		.din(new_net_6512),
		.dout(new_net_6513)
	);

	bfr new_net_2264_bfr_after (
		.din(new_net_6513),
		.dout(new_net_2264)
	);

	bfr new_net_2299_bfr_after (
		.din(_0383_),
		.dout(new_net_2299)
	);

	bfr new_net_6514_bfr_after (
		.din(_0363_),
		.dout(new_net_6514)
	);

	bfr new_net_6515_bfr_after (
		.din(new_net_6514),
		.dout(new_net_6515)
	);

	bfr new_net_6516_bfr_after (
		.din(new_net_6515),
		.dout(new_net_6516)
	);

	bfr new_net_6517_bfr_after (
		.din(new_net_6516),
		.dout(new_net_6517)
	);

	bfr new_net_6518_bfr_after (
		.din(new_net_6517),
		.dout(new_net_6518)
	);

	bfr new_net_6519_bfr_after (
		.din(new_net_6518),
		.dout(new_net_6519)
	);

	bfr new_net_6520_bfr_after (
		.din(new_net_6519),
		.dout(new_net_6520)
	);

	bfr new_net_6521_bfr_after (
		.din(new_net_6520),
		.dout(new_net_6521)
	);

	bfr new_net_6522_bfr_after (
		.din(new_net_6521),
		.dout(new_net_6522)
	);

	bfr new_net_6523_bfr_after (
		.din(new_net_6522),
		.dout(new_net_6523)
	);

	bfr new_net_6524_bfr_after (
		.din(new_net_6523),
		.dout(new_net_6524)
	);

	bfr new_net_6525_bfr_after (
		.din(new_net_6524),
		.dout(new_net_6525)
	);

	bfr new_net_6526_bfr_after (
		.din(new_net_6525),
		.dout(new_net_6526)
	);

	bfr new_net_6527_bfr_after (
		.din(new_net_6526),
		.dout(new_net_6527)
	);

	bfr new_net_6528_bfr_after (
		.din(new_net_6527),
		.dout(new_net_6528)
	);

	bfr new_net_6529_bfr_after (
		.din(new_net_6528),
		.dout(new_net_6529)
	);

	bfr new_net_6530_bfr_after (
		.din(new_net_6529),
		.dout(new_net_6530)
	);

	bfr new_net_6531_bfr_after (
		.din(new_net_6530),
		.dout(new_net_6531)
	);

	bfr new_net_6532_bfr_after (
		.din(new_net_6531),
		.dout(new_net_6532)
	);

	bfr new_net_6533_bfr_after (
		.din(new_net_6532),
		.dout(new_net_6533)
	);

	bfr new_net_6534_bfr_after (
		.din(new_net_6533),
		.dout(new_net_6534)
	);

	bfr new_net_6535_bfr_after (
		.din(new_net_6534),
		.dout(new_net_6535)
	);

	bfr new_net_6536_bfr_after (
		.din(new_net_6535),
		.dout(new_net_6536)
	);

	bfr new_net_2294_bfr_after (
		.din(new_net_6536),
		.dout(new_net_2294)
	);

	bfr new_net_6537_bfr_after (
		.din(G133),
		.dout(new_net_6537)
	);

	bfr new_net_6538_bfr_after (
		.din(new_net_6537),
		.dout(new_net_6538)
	);

	bfr new_net_2237_bfr_after (
		.din(new_net_6538),
		.dout(new_net_2237)
	);

	bfr new_net_6539_bfr_after (
		.din(new_net_2469),
		.dout(new_net_6539)
	);

	bfr new_net_6540_bfr_after (
		.din(new_net_6539),
		.dout(new_net_6540)
	);

	bfr new_net_6541_bfr_after (
		.din(new_net_6540),
		.dout(new_net_6541)
	);

	bfr new_net_6542_bfr_after (
		.din(new_net_6541),
		.dout(new_net_6542)
	);

	bfr new_net_6543_bfr_after (
		.din(new_net_6542),
		.dout(new_net_6543)
	);

	bfr new_net_6544_bfr_after (
		.din(new_net_6543),
		.dout(new_net_6544)
	);

	bfr new_net_6545_bfr_after (
		.din(new_net_6544),
		.dout(new_net_6545)
	);

	bfr new_net_6546_bfr_after (
		.din(new_net_6545),
		.dout(new_net_6546)
	);

	bfr new_net_6547_bfr_after (
		.din(new_net_6546),
		.dout(new_net_6547)
	);

	bfr new_net_6548_bfr_after (
		.din(new_net_6547),
		.dout(new_net_6548)
	);

	bfr G5264_bfr_after (
		.din(new_net_6548),
		.dout(G5264)
	);

	bfr new_net_6549_bfr_after (
		.din(new_net_2353),
		.dout(new_net_6549)
	);

	bfr new_net_6550_bfr_after (
		.din(new_net_6549),
		.dout(new_net_6550)
	);

	bfr new_net_6551_bfr_after (
		.din(new_net_6550),
		.dout(new_net_6551)
	);

	bfr new_net_6552_bfr_after (
		.din(new_net_6551),
		.dout(new_net_6552)
	);

	bfr new_net_6553_bfr_after (
		.din(new_net_6552),
		.dout(new_net_6553)
	);

	bfr new_net_6554_bfr_after (
		.din(new_net_6553),
		.dout(new_net_6554)
	);

	bfr new_net_6555_bfr_after (
		.din(new_net_6554),
		.dout(new_net_6555)
	);

	bfr new_net_6556_bfr_after (
		.din(new_net_6555),
		.dout(new_net_6556)
	);

	bfr new_net_6557_bfr_after (
		.din(new_net_6556),
		.dout(new_net_6557)
	);

	bfr G5310_bfr_after (
		.din(new_net_6557),
		.dout(G5310)
	);

	bfr new_net_6558_bfr_after (
		.din(new_net_2365),
		.dout(new_net_6558)
	);

	bfr new_net_6559_bfr_after (
		.din(new_net_6558),
		.dout(new_net_6559)
	);

	bfr new_net_6560_bfr_after (
		.din(new_net_6559),
		.dout(new_net_6560)
	);

	bfr new_net_6561_bfr_after (
		.din(new_net_6560),
		.dout(new_net_6561)
	);

	bfr new_net_6562_bfr_after (
		.din(new_net_6561),
		.dout(new_net_6562)
	);

	bfr new_net_6563_bfr_after (
		.din(new_net_6562),
		.dout(new_net_6563)
	);

	bfr new_net_6564_bfr_after (
		.din(new_net_6563),
		.dout(new_net_6564)
	);

	bfr new_net_6565_bfr_after (
		.din(new_net_6564),
		.dout(new_net_6565)
	);

	bfr new_net_6566_bfr_after (
		.din(new_net_6565),
		.dout(new_net_6566)
	);

	bfr new_net_6567_bfr_after (
		.din(new_net_6566),
		.dout(new_net_6567)
	);

	bfr new_net_6568_bfr_after (
		.din(new_net_6567),
		.dout(new_net_6568)
	);

	bfr new_net_6569_bfr_after (
		.din(new_net_6568),
		.dout(new_net_6569)
	);

	bfr new_net_6570_bfr_after (
		.din(new_net_6569),
		.dout(new_net_6570)
	);

	bfr new_net_6571_bfr_after (
		.din(new_net_6570),
		.dout(new_net_6571)
	);

	bfr new_net_6572_bfr_after (
		.din(new_net_6571),
		.dout(new_net_6572)
	);

	bfr G5274_bfr_after (
		.din(new_net_6572),
		.dout(G5274)
	);

	bfr new_net_6573_bfr_after (
		.din(new_net_2377),
		.dout(new_net_6573)
	);

	bfr new_net_6574_bfr_after (
		.din(new_net_6573),
		.dout(new_net_6574)
	);

	bfr new_net_6575_bfr_after (
		.din(new_net_6574),
		.dout(new_net_6575)
	);

	bfr new_net_6576_bfr_after (
		.din(new_net_6575),
		.dout(new_net_6576)
	);

	bfr new_net_6577_bfr_after (
		.din(new_net_6576),
		.dout(new_net_6577)
	);

	bfr new_net_6578_bfr_after (
		.din(new_net_6577),
		.dout(new_net_6578)
	);

	bfr new_net_6579_bfr_after (
		.din(new_net_6578),
		.dout(new_net_6579)
	);

	bfr new_net_6580_bfr_after (
		.din(new_net_6579),
		.dout(new_net_6580)
	);

	bfr new_net_6581_bfr_after (
		.din(new_net_6580),
		.dout(new_net_6581)
	);

	bfr new_net_6582_bfr_after (
		.din(new_net_6581),
		.dout(new_net_6582)
	);

	bfr new_net_6583_bfr_after (
		.din(new_net_6582),
		.dout(new_net_6583)
	);

	bfr new_net_6584_bfr_after (
		.din(new_net_6583),
		.dout(new_net_6584)
	);

	bfr new_net_6585_bfr_after (
		.din(new_net_6584),
		.dout(new_net_6585)
	);

	bfr new_net_6586_bfr_after (
		.din(new_net_6585),
		.dout(new_net_6586)
	);

	bfr new_net_6587_bfr_after (
		.din(new_net_6586),
		.dout(new_net_6587)
	);

	bfr new_net_6588_bfr_after (
		.din(new_net_6587),
		.dout(new_net_6588)
	);

	bfr new_net_6589_bfr_after (
		.din(new_net_6588),
		.dout(new_net_6589)
	);

	bfr new_net_6590_bfr_after (
		.din(new_net_6589),
		.dout(new_net_6590)
	);

	bfr new_net_6591_bfr_after (
		.din(new_net_6590),
		.dout(new_net_6591)
	);

	bfr new_net_6592_bfr_after (
		.din(new_net_6591),
		.dout(new_net_6592)
	);

	bfr new_net_6593_bfr_after (
		.din(new_net_6592),
		.dout(new_net_6593)
	);

	bfr new_net_6594_bfr_after (
		.din(new_net_6593),
		.dout(new_net_6594)
	);

	bfr new_net_6595_bfr_after (
		.din(new_net_6594),
		.dout(new_net_6595)
	);

	bfr new_net_6596_bfr_after (
		.din(new_net_6595),
		.dout(new_net_6596)
	);

	bfr new_net_6597_bfr_after (
		.din(new_net_6596),
		.dout(new_net_6597)
	);

	bfr new_net_6598_bfr_after (
		.din(new_net_6597),
		.dout(new_net_6598)
	);

	bfr new_net_6599_bfr_after (
		.din(new_net_6598),
		.dout(new_net_6599)
	);

	bfr G5284_bfr_after (
		.din(new_net_6599),
		.dout(G5284)
	);

	bfr new_net_6600_bfr_after (
		.din(new_net_2389),
		.dout(new_net_6600)
	);

	bfr new_net_6601_bfr_after (
		.din(new_net_6600),
		.dout(new_net_6601)
	);

	bfr new_net_6602_bfr_after (
		.din(new_net_6601),
		.dout(new_net_6602)
	);

	bfr new_net_6603_bfr_after (
		.din(new_net_6602),
		.dout(new_net_6603)
	);

	bfr new_net_6604_bfr_after (
		.din(new_net_6603),
		.dout(new_net_6604)
	);

	bfr new_net_6605_bfr_after (
		.din(new_net_6604),
		.dout(new_net_6605)
	);

	bfr new_net_6606_bfr_after (
		.din(new_net_6605),
		.dout(new_net_6606)
	);

	bfr new_net_6607_bfr_after (
		.din(new_net_6606),
		.dout(new_net_6607)
	);

	bfr new_net_6608_bfr_after (
		.din(new_net_6607),
		.dout(new_net_6608)
	);

	bfr new_net_6609_bfr_after (
		.din(new_net_6608),
		.dout(new_net_6609)
	);

	bfr new_net_6610_bfr_after (
		.din(new_net_6609),
		.dout(new_net_6610)
	);

	bfr new_net_6611_bfr_after (
		.din(new_net_6610),
		.dout(new_net_6611)
	);

	bfr new_net_6612_bfr_after (
		.din(new_net_6611),
		.dout(new_net_6612)
	);

	bfr new_net_6613_bfr_after (
		.din(new_net_6612),
		.dout(new_net_6613)
	);

	bfr new_net_6614_bfr_after (
		.din(new_net_6613),
		.dout(new_net_6614)
	);

	bfr new_net_6615_bfr_after (
		.din(new_net_6614),
		.dout(new_net_6615)
	);

	bfr new_net_6616_bfr_after (
		.din(new_net_6615),
		.dout(new_net_6616)
	);

	bfr new_net_6617_bfr_after (
		.din(new_net_6616),
		.dout(new_net_6617)
	);

	bfr new_net_6618_bfr_after (
		.din(new_net_6617),
		.dout(new_net_6618)
	);

	bfr new_net_6619_bfr_after (
		.din(new_net_6618),
		.dout(new_net_6619)
	);

	bfr new_net_6620_bfr_after (
		.din(new_net_6619),
		.dout(new_net_6620)
	);

	bfr new_net_6621_bfr_after (
		.din(new_net_6620),
		.dout(new_net_6621)
	);

	bfr new_net_6622_bfr_after (
		.din(new_net_6621),
		.dout(new_net_6622)
	);

	bfr new_net_6623_bfr_after (
		.din(new_net_6622),
		.dout(new_net_6623)
	);

	bfr new_net_6624_bfr_after (
		.din(new_net_6623),
		.dout(new_net_6624)
	);

	bfr new_net_6625_bfr_after (
		.din(new_net_6624),
		.dout(new_net_6625)
	);

	bfr new_net_6626_bfr_after (
		.din(new_net_6625),
		.dout(new_net_6626)
	);

	bfr new_net_6627_bfr_after (
		.din(new_net_6626),
		.dout(new_net_6627)
	);

	bfr new_net_6628_bfr_after (
		.din(new_net_6627),
		.dout(new_net_6628)
	);

	bfr new_net_6629_bfr_after (
		.din(new_net_6628),
		.dout(new_net_6629)
	);

	bfr new_net_6630_bfr_after (
		.din(new_net_6629),
		.dout(new_net_6630)
	);

	bfr new_net_6631_bfr_after (
		.din(new_net_6630),
		.dout(new_net_6631)
	);

	bfr new_net_6632_bfr_after (
		.din(new_net_6631),
		.dout(new_net_6632)
	);

	bfr new_net_6633_bfr_after (
		.din(new_net_6632),
		.dout(new_net_6633)
	);

	bfr new_net_6634_bfr_after (
		.din(new_net_6633),
		.dout(new_net_6634)
	);

	bfr new_net_6635_bfr_after (
		.din(new_net_6634),
		.dout(new_net_6635)
	);

	bfr new_net_6636_bfr_after (
		.din(new_net_6635),
		.dout(new_net_6636)
	);

	bfr new_net_6637_bfr_after (
		.din(new_net_6636),
		.dout(new_net_6637)
	);

	bfr new_net_6638_bfr_after (
		.din(new_net_6637),
		.dout(new_net_6638)
	);

	bfr G5212_bfr_after (
		.din(new_net_6638),
		.dout(G5212)
	);

	bfr new_net_6639_bfr_after (
		.din(new_net_2401),
		.dout(new_net_6639)
	);

	bfr new_net_6640_bfr_after (
		.din(new_net_6639),
		.dout(new_net_6640)
	);

	bfr new_net_6641_bfr_after (
		.din(new_net_6640),
		.dout(new_net_6641)
	);

	bfr G5295_bfr_after (
		.din(new_net_6641),
		.dout(G5295)
	);

	bfr new_net_6642_bfr_after (
		.din(new_net_2489),
		.dout(new_net_6642)
	);

	bfr G5312_bfr_after (
		.din(new_net_6642),
		.dout(G5312)
	);

	bfr new_net_6643_bfr_after (
		.din(G59),
		.dout(new_net_6643)
	);

	bfr new_net_6644_bfr_after (
		.din(new_net_6643),
		.dout(new_net_6644)
	);

	bfr new_net_6645_bfr_after (
		.din(new_net_6644),
		.dout(new_net_6645)
	);

	bfr new_net_6646_bfr_after (
		.din(new_net_6645),
		.dout(new_net_6646)
	);

	bfr new_net_2138_bfr_after (
		.din(new_net_6646),
		.dout(new_net_2138)
	);

	bfr new_net_6647_bfr_after (
		.din(_1029_),
		.dout(new_net_6647)
	);

	bfr new_net_6648_bfr_after (
		.din(new_net_6647),
		.dout(new_net_6648)
	);

	bfr new_net_6649_bfr_after (
		.din(new_net_6648),
		.dout(new_net_6649)
	);

	bfr new_net_6650_bfr_after (
		.din(new_net_6649),
		.dout(new_net_6650)
	);

	bfr new_net_6651_bfr_after (
		.din(new_net_6650),
		.dout(new_net_6651)
	);

	bfr new_net_6652_bfr_after (
		.din(new_net_6651),
		.dout(new_net_6652)
	);

	bfr new_net_6653_bfr_after (
		.din(new_net_6652),
		.dout(new_net_6653)
	);

	bfr new_net_6654_bfr_after (
		.din(new_net_6653),
		.dout(new_net_6654)
	);

	bfr new_net_6655_bfr_after (
		.din(new_net_6654),
		.dout(new_net_6655)
	);

	bfr new_net_6656_bfr_after (
		.din(new_net_6655),
		.dout(new_net_6656)
	);

	bfr new_net_6657_bfr_after (
		.din(new_net_6656),
		.dout(new_net_6657)
	);

	bfr new_net_6658_bfr_after (
		.din(new_net_6657),
		.dout(new_net_6658)
	);

	bfr new_net_6659_bfr_after (
		.din(new_net_6658),
		.dout(new_net_6659)
	);

	bfr new_net_6660_bfr_after (
		.din(new_net_6659),
		.dout(new_net_6660)
	);

	bfr new_net_6661_bfr_after (
		.din(new_net_6660),
		.dout(new_net_6661)
	);

	bfr new_net_6662_bfr_after (
		.din(new_net_6661),
		.dout(new_net_6662)
	);

	bfr new_net_6663_bfr_after (
		.din(new_net_6662),
		.dout(new_net_6663)
	);

	bfr new_net_6664_bfr_after (
		.din(new_net_6663),
		.dout(new_net_6664)
	);

	bfr new_net_6665_bfr_after (
		.din(new_net_6664),
		.dout(new_net_6665)
	);

	bfr new_net_6666_bfr_after (
		.din(new_net_6665),
		.dout(new_net_6666)
	);

	bfr new_net_6667_bfr_after (
		.din(new_net_6666),
		.dout(new_net_6667)
	);

	bfr new_net_6668_bfr_after (
		.din(new_net_6667),
		.dout(new_net_6668)
	);

	bfr new_net_2201_bfr_after (
		.din(new_net_6668),
		.dout(new_net_2201)
	);

	bfr new_net_2259_bfr_after (
		.din(_0235_),
		.dout(new_net_2259)
	);

	bfr new_net_6669_bfr_after (
		.din(G19),
		.dout(new_net_6669)
	);

	bfr new_net_6670_bfr_after (
		.din(new_net_6669),
		.dout(new_net_6670)
	);

	bfr new_net_6671_bfr_after (
		.din(new_net_6670),
		.dout(new_net_6671)
	);

	bfr new_net_6672_bfr_after (
		.din(new_net_6671),
		.dout(new_net_6672)
	);

	bfr new_net_2133_bfr_after (
		.din(new_net_6672),
		.dout(new_net_2133)
	);

	bfr new_net_6673_bfr_after (
		.din(_0789_),
		.dout(new_net_6673)
	);

	bfr new_net_6674_bfr_after (
		.din(new_net_6673),
		.dout(new_net_6674)
	);

	bfr new_net_6675_bfr_after (
		.din(new_net_6674),
		.dout(new_net_6675)
	);

	bfr new_net_6676_bfr_after (
		.din(new_net_6675),
		.dout(new_net_6676)
	);

	bfr new_net_6677_bfr_after (
		.din(new_net_6676),
		.dout(new_net_6677)
	);

	bfr new_net_6678_bfr_after (
		.din(new_net_6677),
		.dout(new_net_6678)
	);

	bfr new_net_6679_bfr_after (
		.din(new_net_6678),
		.dout(new_net_6679)
	);

	bfr new_net_6680_bfr_after (
		.din(new_net_6679),
		.dout(new_net_6680)
	);

	bfr new_net_6681_bfr_after (
		.din(new_net_6680),
		.dout(new_net_6681)
	);

	bfr new_net_6682_bfr_after (
		.din(new_net_6681),
		.dout(new_net_6682)
	);

	bfr new_net_6683_bfr_after (
		.din(new_net_6682),
		.dout(new_net_6683)
	);

	bfr new_net_6684_bfr_after (
		.din(new_net_6683),
		.dout(new_net_6684)
	);

	bfr new_net_6685_bfr_after (
		.din(new_net_6684),
		.dout(new_net_6685)
	);

	bfr new_net_2154_bfr_after (
		.din(new_net_6685),
		.dout(new_net_2154)
	);

	bfr new_net_6686_bfr_after (
		.din(_0859_),
		.dout(new_net_6686)
	);

	bfr new_net_6687_bfr_after (
		.din(new_net_6686),
		.dout(new_net_6687)
	);

	bfr new_net_6688_bfr_after (
		.din(new_net_6687),
		.dout(new_net_6688)
	);

	bfr new_net_6689_bfr_after (
		.din(new_net_6688),
		.dout(new_net_6689)
	);

	bfr new_net_6690_bfr_after (
		.din(new_net_6689),
		.dout(new_net_6690)
	);

	bfr new_net_6691_bfr_after (
		.din(new_net_6690),
		.dout(new_net_6691)
	);

	bfr new_net_6692_bfr_after (
		.din(new_net_6691),
		.dout(new_net_6692)
	);

	bfr new_net_6693_bfr_after (
		.din(new_net_6692),
		.dout(new_net_6693)
	);

	bfr new_net_6694_bfr_after (
		.din(new_net_6693),
		.dout(new_net_6694)
	);

	bfr new_net_6695_bfr_after (
		.din(new_net_6694),
		.dout(new_net_6695)
	);

	bfr new_net_6696_bfr_after (
		.din(new_net_6695),
		.dout(new_net_6696)
	);

	bfr new_net_6697_bfr_after (
		.din(new_net_6696),
		.dout(new_net_6697)
	);

	bfr new_net_6698_bfr_after (
		.din(new_net_6697),
		.dout(new_net_6698)
	);

	bfr new_net_6699_bfr_after (
		.din(new_net_6698),
		.dout(new_net_6699)
	);

	bfr new_net_6700_bfr_after (
		.din(new_net_6699),
		.dout(new_net_6700)
	);

	bfr new_net_6701_bfr_after (
		.din(new_net_6700),
		.dout(new_net_6701)
	);

	bfr new_net_6702_bfr_after (
		.din(new_net_6701),
		.dout(new_net_6702)
	);

	bfr new_net_6703_bfr_after (
		.din(new_net_6702),
		.dout(new_net_6703)
	);

	bfr new_net_6704_bfr_after (
		.din(new_net_6703),
		.dout(new_net_6704)
	);

	bfr new_net_6705_bfr_after (
		.din(new_net_6704),
		.dout(new_net_6705)
	);

	bfr new_net_6706_bfr_after (
		.din(new_net_6705),
		.dout(new_net_6706)
	);

	bfr new_net_6707_bfr_after (
		.din(new_net_6706),
		.dout(new_net_6707)
	);

	bfr new_net_6708_bfr_after (
		.din(new_net_6707),
		.dout(new_net_6708)
	);

	bfr new_net_6709_bfr_after (
		.din(new_net_6708),
		.dout(new_net_6709)
	);

	bfr new_net_2175_bfr_after (
		.din(new_net_6709),
		.dout(new_net_2175)
	);

	bfr new_net_6710_bfr_after (
		.din(G34),
		.dout(new_net_6710)
	);

	bfr new_net_2112_bfr_after (
		.din(new_net_6710),
		.dout(new_net_2112)
	);

	bfr new_net_6711_bfr_after (
		.din(G20),
		.dout(new_net_6711)
	);

	bfr new_net_6712_bfr_after (
		.din(new_net_6711),
		.dout(new_net_6712)
	);

	bfr new_net_6713_bfr_after (
		.din(new_net_6712),
		.dout(new_net_6713)
	);

	bfr new_net_6714_bfr_after (
		.din(new_net_6713),
		.dout(new_net_6714)
	);

	bfr new_net_2196_bfr_after (
		.din(new_net_6714),
		.dout(new_net_2196)
	);

	bfr new_net_6715_bfr_after (
		.din(_0307_),
		.dout(new_net_6715)
	);

	bfr new_net_6716_bfr_after (
		.din(new_net_6715),
		.dout(new_net_6716)
	);

	bfr new_net_6717_bfr_after (
		.din(new_net_6716),
		.dout(new_net_6717)
	);

	bfr new_net_6718_bfr_after (
		.din(new_net_6717),
		.dout(new_net_6718)
	);

	bfr new_net_6719_bfr_after (
		.din(new_net_6718),
		.dout(new_net_6719)
	);

	bfr new_net_6720_bfr_after (
		.din(new_net_6719),
		.dout(new_net_6720)
	);

	bfr new_net_6721_bfr_after (
		.din(new_net_6720),
		.dout(new_net_6721)
	);

	bfr new_net_6722_bfr_after (
		.din(new_net_6721),
		.dout(new_net_6722)
	);

	bfr new_net_6723_bfr_after (
		.din(new_net_6722),
		.dout(new_net_6723)
	);

	bfr new_net_6724_bfr_after (
		.din(new_net_6723),
		.dout(new_net_6724)
	);

	bfr new_net_6725_bfr_after (
		.din(new_net_6724),
		.dout(new_net_6725)
	);

	bfr new_net_6726_bfr_after (
		.din(new_net_6725),
		.dout(new_net_6726)
	);

	bfr new_net_6727_bfr_after (
		.din(new_net_6726),
		.dout(new_net_6727)
	);

	bfr new_net_6728_bfr_after (
		.din(new_net_6727),
		.dout(new_net_6728)
	);

	bfr new_net_6729_bfr_after (
		.din(new_net_6728),
		.dout(new_net_6729)
	);

	bfr new_net_6730_bfr_after (
		.din(new_net_6729),
		.dout(new_net_6730)
	);

	bfr new_net_6731_bfr_after (
		.din(new_net_6730),
		.dout(new_net_6731)
	);

	bfr new_net_6732_bfr_after (
		.din(new_net_6731),
		.dout(new_net_6732)
	);

	bfr new_net_6733_bfr_after (
		.din(new_net_6732),
		.dout(new_net_6733)
	);

	bfr new_net_6734_bfr_after (
		.din(new_net_6733),
		.dout(new_net_6734)
	);

	bfr new_net_6735_bfr_after (
		.din(new_net_6734),
		.dout(new_net_6735)
	);

	bfr new_net_6736_bfr_after (
		.din(new_net_6735),
		.dout(new_net_6736)
	);

	bfr new_net_6737_bfr_after (
		.din(new_net_6736),
		.dout(new_net_6737)
	);

	bfr new_net_2280_bfr_after (
		.din(new_net_6737),
		.dout(new_net_2280)
	);

	bfr new_net_6738_bfr_after (
		.din(G49),
		.dout(new_net_6738)
	);

	bfr new_net_6739_bfr_after (
		.din(new_net_6738),
		.dout(new_net_6739)
	);

	bfr new_net_6740_bfr_after (
		.din(new_net_6739),
		.dout(new_net_6740)
	);

	bfr new_net_6741_bfr_after (
		.din(new_net_6740),
		.dout(new_net_6741)
	);

	bfr new_net_2343_bfr_after (
		.din(new_net_6741),
		.dout(new_net_2343)
	);

	bfr new_net_6742_bfr_after (
		.din(_1225_),
		.dout(new_net_6742)
	);

	bfr new_net_6743_bfr_after (
		.din(new_net_6742),
		.dout(new_net_6743)
	);

	bfr new_net_6744_bfr_after (
		.din(new_net_6743),
		.dout(new_net_6744)
	);

	bfr new_net_6745_bfr_after (
		.din(new_net_6744),
		.dout(new_net_6745)
	);

	bfr new_net_6746_bfr_after (
		.din(new_net_6745),
		.dout(new_net_6746)
	);

	bfr new_net_6747_bfr_after (
		.din(new_net_6746),
		.dout(new_net_6747)
	);

	bfr new_net_6748_bfr_after (
		.din(new_net_6747),
		.dout(new_net_6748)
	);

	bfr new_net_6749_bfr_after (
		.din(new_net_6748),
		.dout(new_net_6749)
	);

	bfr new_net_6750_bfr_after (
		.din(new_net_6749),
		.dout(new_net_6750)
	);

	bfr new_net_6751_bfr_after (
		.din(new_net_6750),
		.dout(new_net_6751)
	);

	bfr new_net_6752_bfr_after (
		.din(new_net_6751),
		.dout(new_net_6752)
	);

	bfr new_net_6753_bfr_after (
		.din(new_net_6752),
		.dout(new_net_6753)
	);

	bfr new_net_6754_bfr_after (
		.din(new_net_6753),
		.dout(new_net_6754)
	);

	bfr new_net_6755_bfr_after (
		.din(new_net_6754),
		.dout(new_net_6755)
	);

	bfr new_net_6756_bfr_after (
		.din(new_net_6755),
		.dout(new_net_6756)
	);

	bfr new_net_6757_bfr_after (
		.din(new_net_6756),
		.dout(new_net_6757)
	);

	bfr new_net_6758_bfr_after (
		.din(new_net_6757),
		.dout(new_net_6758)
	);

	bfr new_net_6759_bfr_after (
		.din(new_net_6758),
		.dout(new_net_6759)
	);

	bfr new_net_6760_bfr_after (
		.din(new_net_6759),
		.dout(new_net_6760)
	);

	bfr new_net_6761_bfr_after (
		.din(new_net_6760),
		.dout(new_net_6761)
	);

	bfr new_net_6762_bfr_after (
		.din(new_net_6761),
		.dout(new_net_6762)
	);

	bfr new_net_6763_bfr_after (
		.din(new_net_6762),
		.dout(new_net_6763)
	);

	bfr new_net_6764_bfr_after (
		.din(new_net_6763),
		.dout(new_net_6764)
	);

	bfr new_net_6765_bfr_after (
		.din(new_net_6764),
		.dout(new_net_6765)
	);

	bfr new_net_6766_bfr_after (
		.din(new_net_6765),
		.dout(new_net_6766)
	);

	bfr new_net_6767_bfr_after (
		.din(new_net_6766),
		.dout(new_net_6767)
	);

	bfr new_net_6768_bfr_after (
		.din(new_net_6767),
		.dout(new_net_6768)
	);

	bfr new_net_6769_bfr_after (
		.din(new_net_6768),
		.dout(new_net_6769)
	);

	bfr new_net_6770_bfr_after (
		.din(new_net_6769),
		.dout(new_net_6770)
	);

	bfr new_net_6771_bfr_after (
		.din(new_net_6770),
		.dout(new_net_6771)
	);

	bfr new_net_6772_bfr_after (
		.din(new_net_6771),
		.dout(new_net_6772)
	);

	bfr new_net_6773_bfr_after (
		.din(new_net_6772),
		.dout(new_net_6773)
	);

	bfr new_net_2217_bfr_after (
		.din(new_net_6773),
		.dout(new_net_2217)
	);

	bfr new_net_6774_bfr_after (
		.din(_0395_),
		.dout(new_net_6774)
	);

	bfr new_net_6775_bfr_after (
		.din(new_net_6774),
		.dout(new_net_6775)
	);

	bfr new_net_6776_bfr_after (
		.din(new_net_6775),
		.dout(new_net_6776)
	);

	bfr new_net_6777_bfr_after (
		.din(new_net_6776),
		.dout(new_net_6777)
	);

	bfr new_net_6778_bfr_after (
		.din(new_net_6777),
		.dout(new_net_6778)
	);

	bfr new_net_6779_bfr_after (
		.din(new_net_6778),
		.dout(new_net_6779)
	);

	bfr new_net_6780_bfr_after (
		.din(new_net_6779),
		.dout(new_net_6780)
	);

	bfr new_net_6781_bfr_after (
		.din(new_net_6780),
		.dout(new_net_6781)
	);

	bfr new_net_6782_bfr_after (
		.din(new_net_6781),
		.dout(new_net_6782)
	);

	bfr new_net_6783_bfr_after (
		.din(new_net_6782),
		.dout(new_net_6783)
	);

	bfr new_net_6784_bfr_after (
		.din(new_net_6783),
		.dout(new_net_6784)
	);

	bfr new_net_6785_bfr_after (
		.din(new_net_6784),
		.dout(new_net_6785)
	);

	bfr new_net_6786_bfr_after (
		.din(new_net_6785),
		.dout(new_net_6786)
	);

	bfr new_net_6787_bfr_after (
		.din(new_net_6786),
		.dout(new_net_6787)
	);

	bfr new_net_6788_bfr_after (
		.din(new_net_6787),
		.dout(new_net_6788)
	);

	bfr new_net_6789_bfr_after (
		.din(new_net_6788),
		.dout(new_net_6789)
	);

	bfr new_net_6790_bfr_after (
		.din(new_net_6789),
		.dout(new_net_6790)
	);

	bfr new_net_6791_bfr_after (
		.din(new_net_6790),
		.dout(new_net_6791)
	);

	bfr new_net_6792_bfr_after (
		.din(new_net_6791),
		.dout(new_net_6792)
	);

	bfr new_net_6793_bfr_after (
		.din(new_net_6792),
		.dout(new_net_6793)
	);

	bfr new_net_6794_bfr_after (
		.din(new_net_6793),
		.dout(new_net_6794)
	);

	bfr new_net_6795_bfr_after (
		.din(new_net_6794),
		.dout(new_net_6795)
	);

	bfr new_net_6796_bfr_after (
		.din(new_net_6795),
		.dout(new_net_6796)
	);

	bfr new_net_2301_bfr_after (
		.din(new_net_6796),
		.dout(new_net_2301)
	);

	bfr new_net_6797_bfr_after (
		.din(_0095_),
		.dout(new_net_6797)
	);

	bfr new_net_6798_bfr_after (
		.din(new_net_6797),
		.dout(new_net_6798)
	);

	bfr new_net_6799_bfr_after (
		.din(new_net_6798),
		.dout(new_net_6799)
	);

	bfr new_net_6800_bfr_after (
		.din(new_net_6799),
		.dout(new_net_6800)
	);

	bfr new_net_6801_bfr_after (
		.din(new_net_6800),
		.dout(new_net_6801)
	);

	bfr new_net_6802_bfr_after (
		.din(new_net_6801),
		.dout(new_net_6802)
	);

	bfr new_net_6803_bfr_after (
		.din(new_net_6802),
		.dout(new_net_6803)
	);

	bfr new_net_6804_bfr_after (
		.din(new_net_6803),
		.dout(new_net_6804)
	);

	bfr new_net_6805_bfr_after (
		.din(new_net_6804),
		.dout(new_net_6805)
	);

	bfr new_net_6806_bfr_after (
		.din(new_net_6805),
		.dout(new_net_6806)
	);

	bfr new_net_6807_bfr_after (
		.din(new_net_6806),
		.dout(new_net_6807)
	);

	bfr new_net_6808_bfr_after (
		.din(new_net_6807),
		.dout(new_net_6808)
	);

	bfr new_net_6809_bfr_after (
		.din(new_net_6808),
		.dout(new_net_6809)
	);

	bfr new_net_6810_bfr_after (
		.din(new_net_6809),
		.dout(new_net_6810)
	);

	bfr new_net_6811_bfr_after (
		.din(new_net_6810),
		.dout(new_net_6811)
	);

	bfr new_net_6812_bfr_after (
		.din(new_net_6811),
		.dout(new_net_6812)
	);

	bfr new_net_6813_bfr_after (
		.din(new_net_6812),
		.dout(new_net_6813)
	);

	bfr new_net_6814_bfr_after (
		.din(new_net_6813),
		.dout(new_net_6814)
	);

	bfr new_net_6815_bfr_after (
		.din(new_net_6814),
		.dout(new_net_6815)
	);

	bfr new_net_6816_bfr_after (
		.din(new_net_6815),
		.dout(new_net_6816)
	);

	bfr new_net_6817_bfr_after (
		.din(new_net_6816),
		.dout(new_net_6817)
	);

	bfr new_net_6818_bfr_after (
		.din(new_net_6817),
		.dout(new_net_6818)
	);

	bfr new_net_6819_bfr_after (
		.din(new_net_6818),
		.dout(new_net_6819)
	);

	bfr new_net_6820_bfr_after (
		.din(new_net_6819),
		.dout(new_net_6820)
	);

	bfr new_net_6821_bfr_after (
		.din(new_net_6820),
		.dout(new_net_6821)
	);

	bfr new_net_6822_bfr_after (
		.din(new_net_6821),
		.dout(new_net_6822)
	);

	bfr new_net_6823_bfr_after (
		.din(new_net_6822),
		.dout(new_net_6823)
	);

	bfr new_net_6824_bfr_after (
		.din(new_net_6823),
		.dout(new_net_6824)
	);

	bfr new_net_6825_bfr_after (
		.din(new_net_6824),
		.dout(new_net_6825)
	);

	bfr new_net_6826_bfr_after (
		.din(new_net_6825),
		.dout(new_net_6826)
	);

	bfr new_net_6827_bfr_after (
		.din(new_net_6826),
		.dout(new_net_6827)
	);

	bfr new_net_6828_bfr_after (
		.din(new_net_6827),
		.dout(new_net_6828)
	);

	bfr new_net_2233_bfr_after (
		.din(new_net_6828),
		.dout(new_net_2233)
	);

	bfr new_net_6829_bfr_after (
		.din(G29),
		.dout(new_net_6829)
	);

	bfr new_net_2254_bfr_after (
		.din(new_net_6829),
		.dout(new_net_2254)
	);

	bfr new_net_6830_bfr_after (
		.din(_0455_),
		.dout(new_net_6830)
	);

	bfr new_net_6831_bfr_after (
		.din(new_net_6830),
		.dout(new_net_6831)
	);

	bfr new_net_6832_bfr_after (
		.din(new_net_6831),
		.dout(new_net_6832)
	);

	bfr new_net_6833_bfr_after (
		.din(new_net_6832),
		.dout(new_net_6833)
	);

	bfr new_net_6834_bfr_after (
		.din(new_net_6833),
		.dout(new_net_6834)
	);

	bfr new_net_6835_bfr_after (
		.din(new_net_6834),
		.dout(new_net_6835)
	);

	bfr new_net_6836_bfr_after (
		.din(new_net_6835),
		.dout(new_net_6836)
	);

	bfr new_net_6837_bfr_after (
		.din(new_net_6836),
		.dout(new_net_6837)
	);

	bfr new_net_6838_bfr_after (
		.din(new_net_6837),
		.dout(new_net_6838)
	);

	bfr new_net_6839_bfr_after (
		.din(new_net_6838),
		.dout(new_net_6839)
	);

	bfr new_net_6840_bfr_after (
		.din(new_net_6839),
		.dout(new_net_6840)
	);

	bfr new_net_6841_bfr_after (
		.din(new_net_6840),
		.dout(new_net_6841)
	);

	bfr new_net_6842_bfr_after (
		.din(new_net_6841),
		.dout(new_net_6842)
	);

	bfr new_net_6843_bfr_after (
		.din(new_net_6842),
		.dout(new_net_6843)
	);

	bfr new_net_6844_bfr_after (
		.din(new_net_6843),
		.dout(new_net_6844)
	);

	bfr new_net_6845_bfr_after (
		.din(new_net_6844),
		.dout(new_net_6845)
	);

	bfr new_net_6846_bfr_after (
		.din(new_net_6845),
		.dout(new_net_6846)
	);

	bfr new_net_6847_bfr_after (
		.din(new_net_6846),
		.dout(new_net_6847)
	);

	bfr new_net_6848_bfr_after (
		.din(new_net_6847),
		.dout(new_net_6848)
	);

	bfr new_net_6849_bfr_after (
		.din(new_net_6848),
		.dout(new_net_6849)
	);

	bfr new_net_6850_bfr_after (
		.din(new_net_6849),
		.dout(new_net_6850)
	);

	bfr new_net_6851_bfr_after (
		.din(new_net_6850),
		.dout(new_net_6851)
	);

	bfr new_net_6852_bfr_after (
		.din(new_net_6851),
		.dout(new_net_6852)
	);

	bfr new_net_6853_bfr_after (
		.din(new_net_6852),
		.dout(new_net_6853)
	);

	bfr new_net_6854_bfr_after (
		.din(new_net_6853),
		.dout(new_net_6854)
	);

	bfr new_net_6855_bfr_after (
		.din(new_net_6854),
		.dout(new_net_6855)
	);

	bfr new_net_6856_bfr_after (
		.din(new_net_6855),
		.dout(new_net_6856)
	);

	bfr new_net_6857_bfr_after (
		.din(new_net_6856),
		.dout(new_net_6857)
	);

	bfr new_net_6858_bfr_after (
		.din(new_net_6857),
		.dout(new_net_6858)
	);

	bfr new_net_6859_bfr_after (
		.din(new_net_6858),
		.dout(new_net_6859)
	);

	bfr new_net_2317_bfr_after (
		.din(new_net_6859),
		.dout(new_net_2317)
	);

	bfr new_net_6860_bfr_after (
		.din(_0283_),
		.dout(new_net_6860)
	);

	bfr new_net_2275_bfr_after (
		.din(new_net_6860),
		.dout(new_net_2275)
	);

	bfr new_net_6861_bfr_after (
		.din(_0552_),
		.dout(new_net_6861)
	);

	bfr new_net_6862_bfr_after (
		.din(new_net_6861),
		.dout(new_net_6862)
	);

	bfr new_net_6863_bfr_after (
		.din(new_net_6862),
		.dout(new_net_6863)
	);

	bfr new_net_6864_bfr_after (
		.din(new_net_6863),
		.dout(new_net_6864)
	);

	bfr new_net_6865_bfr_after (
		.din(new_net_6864),
		.dout(new_net_6865)
	);

	bfr new_net_6866_bfr_after (
		.din(new_net_6865),
		.dout(new_net_6866)
	);

	bfr new_net_6867_bfr_after (
		.din(new_net_6866),
		.dout(new_net_6867)
	);

	bfr new_net_6868_bfr_after (
		.din(new_net_6867),
		.dout(new_net_6868)
	);

	bfr new_net_6869_bfr_after (
		.din(new_net_6868),
		.dout(new_net_6869)
	);

	bfr new_net_6870_bfr_after (
		.din(new_net_6869),
		.dout(new_net_6870)
	);

	bfr new_net_6871_bfr_after (
		.din(new_net_6870),
		.dout(new_net_6871)
	);

	bfr new_net_6872_bfr_after (
		.din(new_net_6871),
		.dout(new_net_6872)
	);

	bfr new_net_6873_bfr_after (
		.din(new_net_6872),
		.dout(new_net_6873)
	);

	bfr new_net_6874_bfr_after (
		.din(new_net_6873),
		.dout(new_net_6874)
	);

	bfr new_net_6875_bfr_after (
		.din(new_net_6874),
		.dout(new_net_6875)
	);

	bfr new_net_6876_bfr_after (
		.din(new_net_6875),
		.dout(new_net_6876)
	);

	bfr new_net_6877_bfr_after (
		.din(new_net_6876),
		.dout(new_net_6877)
	);

	bfr new_net_6878_bfr_after (
		.din(new_net_6877),
		.dout(new_net_6878)
	);

	bfr new_net_6879_bfr_after (
		.din(new_net_6878),
		.dout(new_net_6879)
	);

	bfr new_net_6880_bfr_after (
		.din(new_net_6879),
		.dout(new_net_6880)
	);

	bfr new_net_6881_bfr_after (
		.din(new_net_6880),
		.dout(new_net_6881)
	);

	bfr new_net_6882_bfr_after (
		.din(new_net_6881),
		.dout(new_net_6882)
	);

	bfr new_net_6883_bfr_after (
		.din(new_net_6882),
		.dout(new_net_6883)
	);

	bfr new_net_6884_bfr_after (
		.din(new_net_6883),
		.dout(new_net_6884)
	);

	bfr new_net_6885_bfr_after (
		.din(new_net_6884),
		.dout(new_net_6885)
	);

	bfr new_net_6886_bfr_after (
		.din(new_net_6885),
		.dout(new_net_6886)
	);

	bfr new_net_6887_bfr_after (
		.din(new_net_6886),
		.dout(new_net_6887)
	);

	bfr new_net_6888_bfr_after (
		.din(new_net_6887),
		.dout(new_net_6888)
	);

	bfr new_net_6889_bfr_after (
		.din(new_net_6888),
		.dout(new_net_6889)
	);

	bfr new_net_6890_bfr_after (
		.din(new_net_6889),
		.dout(new_net_6890)
	);

	bfr new_net_6891_bfr_after (
		.din(new_net_6890),
		.dout(new_net_6891)
	);

	bfr new_net_2338_bfr_after (
		.din(new_net_6891),
		.dout(new_net_2338)
	);

	bfr new_net_6892_bfr_after (
		.din(G110),
		.dout(new_net_6892)
	);

	bfr new_net_2128_bfr_after (
		.din(new_net_6892),
		.dout(new_net_2128)
	);

	bfr new_net_2149_bfr_after (
		.din(_0750_),
		.dout(new_net_2149)
	);

	bfr new_net_6893_bfr_after (
		.din(G52),
		.dout(new_net_6893)
	);

	bfr new_net_6894_bfr_after (
		.din(new_net_6893),
		.dout(new_net_6894)
	);

	bfr new_net_6895_bfr_after (
		.din(new_net_6894),
		.dout(new_net_6895)
	);

	bfr new_net_6896_bfr_after (
		.din(new_net_6895),
		.dout(new_net_6896)
	);

	bfr new_net_2170_bfr_after (
		.din(new_net_6896),
		.dout(new_net_2170)
	);

	bfr new_net_6897_bfr_after (
		.din(_0987_),
		.dout(new_net_6897)
	);

	bfr new_net_6898_bfr_after (
		.din(new_net_6897),
		.dout(new_net_6898)
	);

	bfr new_net_6899_bfr_after (
		.din(new_net_6898),
		.dout(new_net_6899)
	);

	bfr new_net_6900_bfr_after (
		.din(new_net_6899),
		.dout(new_net_6900)
	);

	bfr new_net_6901_bfr_after (
		.din(new_net_6900),
		.dout(new_net_6901)
	);

	bfr new_net_6902_bfr_after (
		.din(new_net_6901),
		.dout(new_net_6902)
	);

	bfr new_net_6903_bfr_after (
		.din(new_net_6902),
		.dout(new_net_6903)
	);

	bfr new_net_6904_bfr_after (
		.din(new_net_6903),
		.dout(new_net_6904)
	);

	bfr new_net_6905_bfr_after (
		.din(new_net_6904),
		.dout(new_net_6905)
	);

	bfr new_net_6906_bfr_after (
		.din(new_net_6905),
		.dout(new_net_6906)
	);

	bfr new_net_6907_bfr_after (
		.din(new_net_6906),
		.dout(new_net_6907)
	);

	bfr new_net_6908_bfr_after (
		.din(new_net_6907),
		.dout(new_net_6908)
	);

	bfr new_net_6909_bfr_after (
		.din(new_net_6908),
		.dout(new_net_6909)
	);

	bfr new_net_6910_bfr_after (
		.din(new_net_6909),
		.dout(new_net_6910)
	);

	bfr new_net_6911_bfr_after (
		.din(new_net_6910),
		.dout(new_net_6911)
	);

	bfr new_net_6912_bfr_after (
		.din(new_net_6911),
		.dout(new_net_6912)
	);

	bfr new_net_6913_bfr_after (
		.din(new_net_6912),
		.dout(new_net_6913)
	);

	bfr new_net_6914_bfr_after (
		.din(new_net_6913),
		.dout(new_net_6914)
	);

	bfr new_net_6915_bfr_after (
		.din(new_net_6914),
		.dout(new_net_6915)
	);

	bfr new_net_6916_bfr_after (
		.din(new_net_6915),
		.dout(new_net_6916)
	);

	bfr new_net_2191_bfr_after (
		.din(new_net_6916),
		.dout(new_net_2191)
	);

	bfr new_net_6917_bfr_after (
		.din(_0371_),
		.dout(new_net_6917)
	);

	bfr new_net_6918_bfr_after (
		.din(new_net_6917),
		.dout(new_net_6918)
	);

	bfr new_net_6919_bfr_after (
		.din(new_net_6918),
		.dout(new_net_6919)
	);

	bfr new_net_6920_bfr_after (
		.din(new_net_6919),
		.dout(new_net_6920)
	);

	bfr new_net_6921_bfr_after (
		.din(new_net_6920),
		.dout(new_net_6921)
	);

	bfr new_net_6922_bfr_after (
		.din(new_net_6921),
		.dout(new_net_6922)
	);

	bfr new_net_6923_bfr_after (
		.din(new_net_6922),
		.dout(new_net_6923)
	);

	bfr new_net_6924_bfr_after (
		.din(new_net_6923),
		.dout(new_net_6924)
	);

	bfr new_net_6925_bfr_after (
		.din(new_net_6924),
		.dout(new_net_6925)
	);

	bfr new_net_6926_bfr_after (
		.din(new_net_6925),
		.dout(new_net_6926)
	);

	bfr new_net_6927_bfr_after (
		.din(new_net_6926),
		.dout(new_net_6927)
	);

	bfr new_net_6928_bfr_after (
		.din(new_net_6927),
		.dout(new_net_6928)
	);

	bfr new_net_6929_bfr_after (
		.din(new_net_6928),
		.dout(new_net_6929)
	);

	bfr new_net_6930_bfr_after (
		.din(new_net_6929),
		.dout(new_net_6930)
	);

	bfr new_net_6931_bfr_after (
		.din(new_net_6930),
		.dout(new_net_6931)
	);

	bfr new_net_6932_bfr_after (
		.din(new_net_6931),
		.dout(new_net_6932)
	);

	bfr new_net_6933_bfr_after (
		.din(new_net_6932),
		.dout(new_net_6933)
	);

	bfr new_net_6934_bfr_after (
		.din(new_net_6933),
		.dout(new_net_6934)
	);

	bfr new_net_2296_bfr_after (
		.din(new_net_6934),
		.dout(new_net_2296)
	);

	bfr new_net_6935_bfr_after (
		.din(new_net_2481),
		.dout(new_net_6935)
	);

	bfr new_net_6936_bfr_after (
		.din(new_net_6935),
		.dout(new_net_6936)
	);

	bfr new_net_6937_bfr_after (
		.din(new_net_6936),
		.dout(new_net_6937)
	);

	bfr new_net_6938_bfr_after (
		.din(new_net_6937),
		.dout(new_net_6938)
	);

	bfr new_net_6939_bfr_after (
		.din(new_net_6938),
		.dout(new_net_6939)
	);

	bfr new_net_6940_bfr_after (
		.din(new_net_6939),
		.dout(new_net_6940)
	);

	bfr new_net_6941_bfr_after (
		.din(new_net_6940),
		.dout(new_net_6941)
	);

	bfr new_net_6942_bfr_after (
		.din(new_net_6941),
		.dout(new_net_6942)
	);

	bfr new_net_6943_bfr_after (
		.din(new_net_6942),
		.dout(new_net_6943)
	);

	bfr new_net_6944_bfr_after (
		.din(new_net_6943),
		.dout(new_net_6944)
	);

	bfr new_net_6945_bfr_after (
		.din(new_net_6944),
		.dout(new_net_6945)
	);

	bfr G5273_bfr_after (
		.din(new_net_6945),
		.dout(G5273)
	);

	bfr new_net_6946_bfr_after (
		.din(new_net_2501),
		.dout(new_net_6946)
	);

	bfr new_net_6947_bfr_after (
		.din(new_net_6946),
		.dout(new_net_6947)
	);

	bfr new_net_6948_bfr_after (
		.din(new_net_6947),
		.dout(new_net_6948)
	);

	bfr new_net_6949_bfr_after (
		.din(new_net_6948),
		.dout(new_net_6949)
	);

	bfr new_net_6950_bfr_after (
		.din(new_net_6949),
		.dout(new_net_6950)
	);

	bfr new_net_6951_bfr_after (
		.din(new_net_6950),
		.dout(new_net_6951)
	);

	bfr new_net_6952_bfr_after (
		.din(new_net_6951),
		.dout(new_net_6952)
	);

	bfr new_net_6953_bfr_after (
		.din(new_net_6952),
		.dout(new_net_6953)
	);

	bfr new_net_6954_bfr_after (
		.din(new_net_6953),
		.dout(new_net_6954)
	);

	bfr new_net_6955_bfr_after (
		.din(new_net_6954),
		.dout(new_net_6955)
	);

	bfr new_net_6956_bfr_after (
		.din(new_net_6955),
		.dout(new_net_6956)
	);

	bfr G5268_bfr_after (
		.din(new_net_6956),
		.dout(G5268)
	);

	bfr new_net_2228_bfr_after (
		.din(_0080_),
		.dout(new_net_2228)
	);

	bfr new_net_6957_bfr_after (
		.din(_0220_),
		.dout(new_net_6957)
	);

	bfr new_net_2249_bfr_after (
		.din(new_net_6957),
		.dout(new_net_2249)
	);

	bfr new_net_6958_bfr_after (
		.din(_0438_),
		.dout(new_net_6958)
	);

	bfr new_net_6959_bfr_after (
		.din(new_net_6958),
		.dout(new_net_6959)
	);

	bfr new_net_6960_bfr_after (
		.din(new_net_6959),
		.dout(new_net_6960)
	);

	bfr new_net_6961_bfr_after (
		.din(new_net_6960),
		.dout(new_net_6961)
	);

	bfr new_net_6962_bfr_after (
		.din(new_net_6961),
		.dout(new_net_6962)
	);

	bfr new_net_6963_bfr_after (
		.din(new_net_6962),
		.dout(new_net_6963)
	);

	bfr new_net_6964_bfr_after (
		.din(new_net_6963),
		.dout(new_net_6964)
	);

	bfr new_net_6965_bfr_after (
		.din(new_net_6964),
		.dout(new_net_6965)
	);

	bfr new_net_6966_bfr_after (
		.din(new_net_6965),
		.dout(new_net_6966)
	);

	bfr new_net_2312_bfr_after (
		.din(new_net_6966),
		.dout(new_net_2312)
	);

	bfr new_net_6967_bfr_after (
		.din(_0278_),
		.dout(new_net_6967)
	);

	bfr new_net_2270_bfr_after (
		.din(new_net_6967),
		.dout(new_net_2270)
	);

	bfr new_net_6968_bfr_after (
		.din(_0524_),
		.dout(new_net_6968)
	);

	bfr new_net_6969_bfr_after (
		.din(new_net_6968),
		.dout(new_net_6969)
	);

	bfr new_net_6970_bfr_after (
		.din(new_net_6969),
		.dout(new_net_6970)
	);

	bfr new_net_6971_bfr_after (
		.din(new_net_6970),
		.dout(new_net_6971)
	);

	bfr new_net_6972_bfr_after (
		.din(new_net_6971),
		.dout(new_net_6972)
	);

	bfr new_net_6973_bfr_after (
		.din(new_net_6972),
		.dout(new_net_6973)
	);

	bfr new_net_6974_bfr_after (
		.din(new_net_6973),
		.dout(new_net_6974)
	);

	bfr new_net_6975_bfr_after (
		.din(new_net_6974),
		.dout(new_net_6975)
	);

	bfr new_net_6976_bfr_after (
		.din(new_net_6975),
		.dout(new_net_6976)
	);

	bfr new_net_6977_bfr_after (
		.din(new_net_6976),
		.dout(new_net_6977)
	);

	bfr new_net_6978_bfr_after (
		.din(new_net_6977),
		.dout(new_net_6978)
	);

	bfr new_net_6979_bfr_after (
		.din(new_net_6978),
		.dout(new_net_6979)
	);

	bfr new_net_6980_bfr_after (
		.din(new_net_6979),
		.dout(new_net_6980)
	);

	bfr new_net_6981_bfr_after (
		.din(new_net_6980),
		.dout(new_net_6981)
	);

	bfr new_net_6982_bfr_after (
		.din(new_net_6981),
		.dout(new_net_6982)
	);

	bfr new_net_6983_bfr_after (
		.din(new_net_6982),
		.dout(new_net_6983)
	);

	bfr new_net_2333_bfr_after (
		.din(new_net_6983),
		.dout(new_net_2333)
	);

	bfr new_net_2123_bfr_after (
		.din(_0611_),
		.dout(new_net_2123)
	);

	bfr new_net_6984_bfr_after (
		.din(G53),
		.dout(new_net_6984)
	);

	bfr new_net_6985_bfr_after (
		.din(new_net_6984),
		.dout(new_net_6985)
	);

	bfr new_net_6986_bfr_after (
		.din(new_net_6985),
		.dout(new_net_6986)
	);

	bfr new_net_6987_bfr_after (
		.din(new_net_6986),
		.dout(new_net_6987)
	);

	bfr new_net_2144_bfr_after (
		.din(new_net_6987),
		.dout(new_net_2144)
	);

	bfr new_net_2165_bfr_after (
		.din(_0835_),
		.dout(new_net_2165)
	);

	bfr new_net_6988_bfr_after (
		.din(G93),
		.dout(new_net_6988)
	);

	bfr new_net_2186_bfr_after (
		.din(new_net_6988),
		.dout(new_net_2186)
	);

	bfr new_net_6989_bfr_after (
		.din(_1048_),
		.dout(new_net_6989)
	);

	bfr new_net_6990_bfr_after (
		.din(new_net_6989),
		.dout(new_net_6990)
	);

	bfr new_net_6991_bfr_after (
		.din(new_net_6990),
		.dout(new_net_6991)
	);

	bfr new_net_6992_bfr_after (
		.din(new_net_6991),
		.dout(new_net_6992)
	);

	bfr new_net_2204_bfr_after (
		.din(new_net_6992),
		.dout(new_net_2204)
	);

	bfr new_net_6993_bfr_after (
		.din(_0349_),
		.dout(new_net_6993)
	);

	bfr new_net_6994_bfr_after (
		.din(new_net_6993),
		.dout(new_net_6994)
	);

	bfr new_net_6995_bfr_after (
		.din(new_net_6994),
		.dout(new_net_6995)
	);

	bfr new_net_6996_bfr_after (
		.din(new_net_6995),
		.dout(new_net_6996)
	);

	bfr new_net_6997_bfr_after (
		.din(new_net_6996),
		.dout(new_net_6997)
	);

	bfr new_net_6998_bfr_after (
		.din(new_net_6997),
		.dout(new_net_6998)
	);

	bfr new_net_6999_bfr_after (
		.din(new_net_6998),
		.dout(new_net_6999)
	);

	bfr new_net_7000_bfr_after (
		.din(new_net_6999),
		.dout(new_net_7000)
	);

	bfr new_net_7001_bfr_after (
		.din(new_net_7000),
		.dout(new_net_7001)
	);

	bfr new_net_7002_bfr_after (
		.din(new_net_7001),
		.dout(new_net_7002)
	);

	bfr new_net_7003_bfr_after (
		.din(new_net_7002),
		.dout(new_net_7003)
	);

	bfr new_net_7004_bfr_after (
		.din(new_net_7003),
		.dout(new_net_7004)
	);

	bfr new_net_7005_bfr_after (
		.din(new_net_7004),
		.dout(new_net_7005)
	);

	bfr new_net_7006_bfr_after (
		.din(new_net_7005),
		.dout(new_net_7006)
	);

	bfr new_net_7007_bfr_after (
		.din(new_net_7006),
		.dout(new_net_7007)
	);

	bfr new_net_7008_bfr_after (
		.din(new_net_7007),
		.dout(new_net_7008)
	);

	bfr new_net_7009_bfr_after (
		.din(new_net_7008),
		.dout(new_net_7009)
	);

	bfr new_net_7010_bfr_after (
		.din(new_net_7009),
		.dout(new_net_7010)
	);

	bfr new_net_7011_bfr_after (
		.din(new_net_7010),
		.dout(new_net_7011)
	);

	bfr new_net_7012_bfr_after (
		.din(new_net_7011),
		.dout(new_net_7012)
	);

	bfr new_net_7013_bfr_after (
		.din(new_net_7012),
		.dout(new_net_7013)
	);

	bfr new_net_7014_bfr_after (
		.din(new_net_7013),
		.dout(new_net_7014)
	);

	bfr new_net_2291_bfr_after (
		.din(new_net_7014),
		.dout(new_net_2291)
	);

	bfr new_net_7015_bfr_after (
		.din(new_net_2355),
		.dout(new_net_7015)
	);

	bfr new_net_7016_bfr_after (
		.din(new_net_7015),
		.dout(new_net_7016)
	);

	bfr G5296_bfr_after (
		.din(new_net_7016),
		.dout(G5296)
	);

	bfr new_net_2223_bfr_after (
		.din(_0010_),
		.dout(new_net_2223)
	);

	bfr new_net_7017_bfr_after (
		.din(_0419_),
		.dout(new_net_7017)
	);

	bfr new_net_7018_bfr_after (
		.din(new_net_7017),
		.dout(new_net_7018)
	);

	bfr new_net_7019_bfr_after (
		.din(new_net_7018),
		.dout(new_net_7019)
	);

	bfr new_net_7020_bfr_after (
		.din(new_net_7019),
		.dout(new_net_7020)
	);

	bfr new_net_7021_bfr_after (
		.din(new_net_7020),
		.dout(new_net_7021)
	);

	bfr new_net_7022_bfr_after (
		.din(new_net_7021),
		.dout(new_net_7022)
	);

	bfr new_net_7023_bfr_after (
		.din(new_net_7022),
		.dout(new_net_7023)
	);

	bfr new_net_7024_bfr_after (
		.din(new_net_7023),
		.dout(new_net_7024)
	);

	bfr new_net_7025_bfr_after (
		.din(new_net_7024),
		.dout(new_net_7025)
	);

	bfr new_net_7026_bfr_after (
		.din(new_net_7025),
		.dout(new_net_7026)
	);

	bfr new_net_7027_bfr_after (
		.din(new_net_7026),
		.dout(new_net_7027)
	);

	bfr new_net_7028_bfr_after (
		.din(new_net_7027),
		.dout(new_net_7028)
	);

	bfr new_net_7029_bfr_after (
		.din(new_net_7028),
		.dout(new_net_7029)
	);

	bfr new_net_7030_bfr_after (
		.din(new_net_7029),
		.dout(new_net_7030)
	);

	bfr new_net_7031_bfr_after (
		.din(new_net_7030),
		.dout(new_net_7031)
	);

	bfr new_net_7032_bfr_after (
		.din(new_net_7031),
		.dout(new_net_7032)
	);

	bfr new_net_7033_bfr_after (
		.din(new_net_7032),
		.dout(new_net_7033)
	);

	bfr new_net_7034_bfr_after (
		.din(new_net_7033),
		.dout(new_net_7034)
	);

	bfr new_net_7035_bfr_after (
		.din(new_net_7034),
		.dout(new_net_7035)
	);

	bfr new_net_7036_bfr_after (
		.din(new_net_7035),
		.dout(new_net_7036)
	);

	bfr new_net_7037_bfr_after (
		.din(new_net_7036),
		.dout(new_net_7037)
	);

	bfr new_net_7038_bfr_after (
		.din(new_net_7037),
		.dout(new_net_7038)
	);

	bfr new_net_2307_bfr_after (
		.din(new_net_7038),
		.dout(new_net_2307)
	);

	bfr new_net_7039_bfr_after (
		.din(new_net_2417),
		.dout(new_net_7039)
	);

	bfr new_net_7040_bfr_after (
		.din(new_net_7039),
		.dout(new_net_7040)
	);

	bfr new_net_7041_bfr_after (
		.din(new_net_7040),
		.dout(new_net_7041)
	);

	bfr new_net_7042_bfr_after (
		.din(new_net_7041),
		.dout(new_net_7042)
	);

	bfr new_net_7043_bfr_after (
		.din(new_net_7042),
		.dout(new_net_7043)
	);

	bfr new_net_7044_bfr_after (
		.din(new_net_7043),
		.dout(new_net_7044)
	);

	bfr new_net_7045_bfr_after (
		.din(new_net_7044),
		.dout(new_net_7045)
	);

	bfr new_net_7046_bfr_after (
		.din(new_net_7045),
		.dout(new_net_7046)
	);

	bfr new_net_7047_bfr_after (
		.din(new_net_7046),
		.dout(new_net_7047)
	);

	bfr G5263_bfr_after (
		.din(new_net_7047),
		.dout(G5263)
	);

	bfr new_net_2244_bfr_after (
		.din(_0217_),
		.dout(new_net_2244)
	);

	bfr new_net_7048_bfr_after (
		.din(_0504_),
		.dout(new_net_7048)
	);

	bfr new_net_7049_bfr_after (
		.din(new_net_7048),
		.dout(new_net_7049)
	);

	bfr new_net_7050_bfr_after (
		.din(new_net_7049),
		.dout(new_net_7050)
	);

	bfr new_net_7051_bfr_after (
		.din(new_net_7050),
		.dout(new_net_7051)
	);

	bfr new_net_7052_bfr_after (
		.din(new_net_7051),
		.dout(new_net_7052)
	);

	bfr new_net_7053_bfr_after (
		.din(new_net_7052),
		.dout(new_net_7053)
	);

	bfr new_net_7054_bfr_after (
		.din(new_net_7053),
		.dout(new_net_7054)
	);

	bfr new_net_7055_bfr_after (
		.din(new_net_7054),
		.dout(new_net_7055)
	);

	bfr new_net_7056_bfr_after (
		.din(new_net_7055),
		.dout(new_net_7056)
	);

	bfr new_net_7057_bfr_after (
		.din(new_net_7056),
		.dout(new_net_7057)
	);

	bfr new_net_7058_bfr_after (
		.din(new_net_7057),
		.dout(new_net_7058)
	);

	bfr new_net_7059_bfr_after (
		.din(new_net_7058),
		.dout(new_net_7059)
	);

	bfr new_net_7060_bfr_after (
		.din(new_net_7059),
		.dout(new_net_7060)
	);

	bfr new_net_7061_bfr_after (
		.din(new_net_7060),
		.dout(new_net_7061)
	);

	bfr new_net_7062_bfr_after (
		.din(new_net_7061),
		.dout(new_net_7062)
	);

	bfr new_net_7063_bfr_after (
		.din(new_net_7062),
		.dout(new_net_7063)
	);

	bfr new_net_7064_bfr_after (
		.din(new_net_7063),
		.dout(new_net_7064)
	);

	bfr new_net_7065_bfr_after (
		.din(new_net_7064),
		.dout(new_net_7065)
	);

	bfr new_net_7066_bfr_after (
		.din(new_net_7065),
		.dout(new_net_7066)
	);

	bfr new_net_7067_bfr_after (
		.din(new_net_7066),
		.dout(new_net_7067)
	);

	bfr new_net_7068_bfr_after (
		.din(new_net_7067),
		.dout(new_net_7068)
	);

	bfr new_net_7069_bfr_after (
		.din(new_net_7068),
		.dout(new_net_7069)
	);

	bfr new_net_7070_bfr_after (
		.din(new_net_7069),
		.dout(new_net_7070)
	);

	bfr new_net_7071_bfr_after (
		.din(new_net_7070),
		.dout(new_net_7071)
	);

	bfr new_net_7072_bfr_after (
		.din(new_net_7071),
		.dout(new_net_7072)
	);

	bfr new_net_7073_bfr_after (
		.din(new_net_7072),
		.dout(new_net_7073)
	);

	bfr new_net_7074_bfr_after (
		.din(new_net_7073),
		.dout(new_net_7074)
	);

	bfr new_net_7075_bfr_after (
		.din(new_net_7074),
		.dout(new_net_7075)
	);

	bfr new_net_2328_bfr_after (
		.din(new_net_7075),
		.dout(new_net_2328)
	);

	bfr new_net_7076_bfr_after (
		.din(_0264_),
		.dout(new_net_7076)
	);

	bfr new_net_7077_bfr_after (
		.din(new_net_7076),
		.dout(new_net_7077)
	);

	bfr new_net_2265_bfr_after (
		.din(new_net_7077),
		.dout(new_net_2265)
	);

	bfr new_net_7078_bfr_after (
		.din(_0712_),
		.dout(new_net_7078)
	);

	bfr new_net_7079_bfr_after (
		.din(new_net_7078),
		.dout(new_net_7079)
	);

	bfr new_net_7080_bfr_after (
		.din(new_net_7079),
		.dout(new_net_7080)
	);

	bfr new_net_7081_bfr_after (
		.din(new_net_7080),
		.dout(new_net_7081)
	);

	bfr new_net_7082_bfr_after (
		.din(new_net_7081),
		.dout(new_net_7082)
	);

	bfr new_net_7083_bfr_after (
		.din(new_net_7082),
		.dout(new_net_7083)
	);

	bfr new_net_7084_bfr_after (
		.din(new_net_7083),
		.dout(new_net_7084)
	);

	bfr new_net_7085_bfr_after (
		.din(new_net_7084),
		.dout(new_net_7085)
	);

	bfr new_net_7086_bfr_after (
		.din(new_net_7085),
		.dout(new_net_7086)
	);

	bfr new_net_7087_bfr_after (
		.din(new_net_7086),
		.dout(new_net_7087)
	);

	bfr new_net_7088_bfr_after (
		.din(new_net_7087),
		.dout(new_net_7088)
	);

	bfr new_net_7089_bfr_after (
		.din(new_net_7088),
		.dout(new_net_7089)
	);

	bfr new_net_7090_bfr_after (
		.din(new_net_7089),
		.dout(new_net_7090)
	);

	bfr new_net_2139_bfr_after (
		.din(new_net_7090),
		.dout(new_net_2139)
	);

	bfr new_net_7091_bfr_after (
		.din(G56),
		.dout(new_net_7091)
	);

	bfr new_net_7092_bfr_after (
		.din(new_net_7091),
		.dout(new_net_7092)
	);

	bfr new_net_7093_bfr_after (
		.din(new_net_7092),
		.dout(new_net_7093)
	);

	bfr new_net_7094_bfr_after (
		.din(new_net_7093),
		.dout(new_net_7094)
	);

	bfr new_net_2160_bfr_after (
		.din(new_net_7094),
		.dout(new_net_2160)
	);

	bfr new_net_7095_bfr_after (
		.din(_0911_),
		.dout(new_net_7095)
	);

	bfr new_net_7096_bfr_after (
		.din(new_net_7095),
		.dout(new_net_7096)
	);

	bfr new_net_7097_bfr_after (
		.din(new_net_7096),
		.dout(new_net_7097)
	);

	bfr new_net_7098_bfr_after (
		.din(new_net_7097),
		.dout(new_net_7098)
	);

	bfr new_net_7099_bfr_after (
		.din(new_net_7098),
		.dout(new_net_7099)
	);

	bfr new_net_7100_bfr_after (
		.din(new_net_7099),
		.dout(new_net_7100)
	);

	bfr new_net_7101_bfr_after (
		.din(new_net_7100),
		.dout(new_net_7101)
	);

	bfr new_net_7102_bfr_after (
		.din(new_net_7101),
		.dout(new_net_7102)
	);

	bfr new_net_7103_bfr_after (
		.din(new_net_7102),
		.dout(new_net_7103)
	);

	bfr new_net_7104_bfr_after (
		.din(new_net_7103),
		.dout(new_net_7104)
	);

	bfr new_net_7105_bfr_after (
		.din(new_net_7104),
		.dout(new_net_7105)
	);

	bfr new_net_7106_bfr_after (
		.din(new_net_7105),
		.dout(new_net_7106)
	);

	bfr new_net_7107_bfr_after (
		.din(new_net_7106),
		.dout(new_net_7107)
	);

	bfr new_net_7108_bfr_after (
		.din(new_net_7107),
		.dout(new_net_7108)
	);

	bfr new_net_7109_bfr_after (
		.din(new_net_7108),
		.dout(new_net_7109)
	);

	bfr new_net_7110_bfr_after (
		.din(new_net_7109),
		.dout(new_net_7110)
	);

	bfr new_net_7111_bfr_after (
		.din(new_net_7110),
		.dout(new_net_7111)
	);

	bfr new_net_7112_bfr_after (
		.din(new_net_7111),
		.dout(new_net_7112)
	);

	bfr new_net_7113_bfr_after (
		.din(new_net_7112),
		.dout(new_net_7113)
	);

	bfr new_net_7114_bfr_after (
		.din(new_net_7113),
		.dout(new_net_7114)
	);

	bfr new_net_7115_bfr_after (
		.din(new_net_7114),
		.dout(new_net_7115)
	);

	bfr new_net_2181_bfr_after (
		.din(new_net_7115),
		.dout(new_net_2181)
	);

	bfr new_net_7116_bfr_after (
		.din(G32),
		.dout(new_net_7116)
	);

	bfr new_net_7117_bfr_after (
		.din(new_net_7116),
		.dout(new_net_7117)
	);

	bfr new_net_7118_bfr_after (
		.din(new_net_7117),
		.dout(new_net_7118)
	);

	bfr new_net_2118_bfr_after (
		.din(new_net_7118),
		.dout(new_net_2118)
	);

	bfr new_net_7119_bfr_after (
		.din(new_net_2435),
		.dout(new_net_7119)
	);

	bfr new_net_7120_bfr_after (
		.din(new_net_7119),
		.dout(new_net_7120)
	);

	bfr new_net_7121_bfr_after (
		.din(new_net_7120),
		.dout(new_net_7121)
	);

	bfr new_net_7122_bfr_after (
		.din(new_net_7121),
		.dout(new_net_7122)
	);

	bfr new_net_7123_bfr_after (
		.din(new_net_7122),
		.dout(new_net_7123)
	);

	bfr new_net_7124_bfr_after (
		.din(new_net_7123),
		.dout(new_net_7124)
	);

	bfr new_net_7125_bfr_after (
		.din(new_net_7124),
		.dout(new_net_7125)
	);

	bfr new_net_7126_bfr_after (
		.din(new_net_7125),
		.dout(new_net_7126)
	);

	bfr new_net_7127_bfr_after (
		.din(new_net_7126),
		.dout(new_net_7127)
	);

	bfr new_net_7128_bfr_after (
		.din(new_net_7127),
		.dout(new_net_7128)
	);

	bfr new_net_7129_bfr_after (
		.din(new_net_7128),
		.dout(new_net_7129)
	);

	bfr new_net_7130_bfr_after (
		.din(new_net_7129),
		.dout(new_net_7130)
	);

	bfr new_net_7131_bfr_after (
		.din(new_net_7130),
		.dout(new_net_7131)
	);

	bfr new_net_7132_bfr_after (
		.din(new_net_7131),
		.dout(new_net_7132)
	);

	bfr new_net_7133_bfr_after (
		.din(new_net_7132),
		.dout(new_net_7133)
	);

	bfr new_net_7134_bfr_after (
		.din(new_net_7133),
		.dout(new_net_7134)
	);

	bfr new_net_7135_bfr_after (
		.din(new_net_7134),
		.dout(new_net_7135)
	);

	bfr new_net_7136_bfr_after (
		.din(new_net_7135),
		.dout(new_net_7136)
	);

	bfr new_net_7137_bfr_after (
		.din(new_net_7136),
		.dout(new_net_7137)
	);

	bfr new_net_7138_bfr_after (
		.din(new_net_7137),
		.dout(new_net_7138)
	);

	bfr new_net_7139_bfr_after (
		.din(new_net_7138),
		.dout(new_net_7139)
	);

	bfr new_net_7140_bfr_after (
		.din(new_net_7139),
		.dout(new_net_7140)
	);

	bfr new_net_7141_bfr_after (
		.din(new_net_7140),
		.dout(new_net_7141)
	);

	bfr new_net_7142_bfr_after (
		.din(new_net_7141),
		.dout(new_net_7142)
	);

	bfr new_net_7143_bfr_after (
		.din(new_net_7142),
		.dout(new_net_7143)
	);

	bfr new_net_7144_bfr_after (
		.din(new_net_7143),
		.dout(new_net_7144)
	);

	bfr new_net_7145_bfr_after (
		.din(new_net_7144),
		.dout(new_net_7145)
	);

	bfr new_net_7146_bfr_after (
		.din(new_net_7145),
		.dout(new_net_7146)
	);

	bfr new_net_7147_bfr_after (
		.din(new_net_7146),
		.dout(new_net_7147)
	);

	bfr new_net_7148_bfr_after (
		.din(new_net_7147),
		.dout(new_net_7148)
	);

	bfr new_net_7149_bfr_after (
		.din(new_net_7148),
		.dout(new_net_7149)
	);

	bfr new_net_7150_bfr_after (
		.din(new_net_7149),
		.dout(new_net_7150)
	);

	bfr new_net_7151_bfr_after (
		.din(new_net_7150),
		.dout(new_net_7151)
	);

	bfr new_net_7152_bfr_after (
		.din(new_net_7151),
		.dout(new_net_7152)
	);

	bfr new_net_7153_bfr_after (
		.din(new_net_7152),
		.dout(new_net_7153)
	);

	bfr new_net_7154_bfr_after (
		.din(new_net_7153),
		.dout(new_net_7154)
	);

	bfr new_net_7155_bfr_after (
		.din(new_net_7154),
		.dout(new_net_7155)
	);

	bfr new_net_7156_bfr_after (
		.din(new_net_7155),
		.dout(new_net_7156)
	);

	bfr new_net_7157_bfr_after (
		.din(new_net_7156),
		.dout(new_net_7157)
	);

	bfr G5210_bfr_after (
		.din(new_net_7157),
		.dout(G5210)
	);

	bfr new_net_7158_bfr_after (
		.din(_0470_),
		.dout(new_net_7158)
	);

	bfr new_net_2322_bfr_after (
		.din(new_net_7158),
		.dout(new_net_2322)
	);

	bfr new_net_7159_bfr_after (
		.din(new_net_2415),
		.dout(new_net_7159)
	);

	bfr new_net_7160_bfr_after (
		.din(new_net_7159),
		.dout(new_net_7160)
	);

	bfr new_net_7161_bfr_after (
		.din(new_net_7160),
		.dout(new_net_7161)
	);

	bfr new_net_7162_bfr_after (
		.din(new_net_7161),
		.dout(new_net_7162)
	);

	bfr new_net_7163_bfr_after (
		.din(new_net_7162),
		.dout(new_net_7163)
	);

	bfr new_net_7164_bfr_after (
		.din(new_net_7163),
		.dout(new_net_7164)
	);

	bfr new_net_7165_bfr_after (
		.din(new_net_7164),
		.dout(new_net_7165)
	);

	bfr new_net_7166_bfr_after (
		.din(new_net_7165),
		.dout(new_net_7166)
	);

	bfr new_net_7167_bfr_after (
		.din(new_net_7166),
		.dout(new_net_7167)
	);

	bfr new_net_7168_bfr_after (
		.din(new_net_7167),
		.dout(new_net_7168)
	);

	bfr new_net_7169_bfr_after (
		.din(new_net_7168),
		.dout(new_net_7169)
	);

	bfr new_net_7170_bfr_after (
		.din(new_net_7169),
		.dout(new_net_7170)
	);

	bfr new_net_7171_bfr_after (
		.din(new_net_7170),
		.dout(new_net_7171)
	);

	bfr new_net_7172_bfr_after (
		.din(new_net_7171),
		.dout(new_net_7172)
	);

	bfr new_net_7173_bfr_after (
		.din(new_net_7172),
		.dout(new_net_7173)
	);

	bfr new_net_7174_bfr_after (
		.din(new_net_7173),
		.dout(new_net_7174)
	);

	bfr new_net_7175_bfr_after (
		.din(new_net_7174),
		.dout(new_net_7175)
	);

	bfr new_net_7176_bfr_after (
		.din(new_net_7175),
		.dout(new_net_7176)
	);

	bfr new_net_7177_bfr_after (
		.din(new_net_7176),
		.dout(new_net_7177)
	);

	bfr new_net_7178_bfr_after (
		.din(new_net_7177),
		.dout(new_net_7178)
	);

	bfr new_net_7179_bfr_after (
		.din(new_net_7178),
		.dout(new_net_7179)
	);

	bfr new_net_7180_bfr_after (
		.din(new_net_7179),
		.dout(new_net_7180)
	);

	bfr new_net_7181_bfr_after (
		.din(new_net_7180),
		.dout(new_net_7181)
	);

	bfr new_net_7182_bfr_after (
		.din(new_net_7181),
		.dout(new_net_7182)
	);

	bfr new_net_7183_bfr_after (
		.din(new_net_7182),
		.dout(new_net_7183)
	);

	bfr new_net_7184_bfr_after (
		.din(new_net_7183),
		.dout(new_net_7184)
	);

	bfr new_net_7185_bfr_after (
		.din(new_net_7184),
		.dout(new_net_7185)
	);

	bfr new_net_7186_bfr_after (
		.din(new_net_7185),
		.dout(new_net_7186)
	);

	bfr new_net_7187_bfr_after (
		.din(new_net_7186),
		.dout(new_net_7187)
	);

	bfr new_net_7188_bfr_after (
		.din(new_net_7187),
		.dout(new_net_7188)
	);

	bfr new_net_7189_bfr_after (
		.din(new_net_7188),
		.dout(new_net_7189)
	);

	bfr new_net_7190_bfr_after (
		.din(new_net_7189),
		.dout(new_net_7190)
	);

	bfr new_net_7191_bfr_after (
		.din(new_net_7190),
		.dout(new_net_7191)
	);

	bfr new_net_7192_bfr_after (
		.din(new_net_7191),
		.dout(new_net_7192)
	);

	bfr new_net_7193_bfr_after (
		.din(new_net_7192),
		.dout(new_net_7193)
	);

	bfr new_net_7194_bfr_after (
		.din(new_net_7193),
		.dout(new_net_7194)
	);

	bfr new_net_7195_bfr_after (
		.din(new_net_7194),
		.dout(new_net_7195)
	);

	bfr new_net_7196_bfr_after (
		.din(new_net_7195),
		.dout(new_net_7196)
	);

	bfr new_net_7197_bfr_after (
		.din(new_net_7196),
		.dout(new_net_7197)
	);

	bfr G5195_bfr_after (
		.din(new_net_7197),
		.dout(G5195)
	);

	bfr new_net_7198_bfr_after (
		.din(G31),
		.dout(new_net_7198)
	);

	bfr new_net_2255_bfr_after (
		.din(new_net_7198),
		.dout(new_net_2255)
	);

	bfr new_net_7199_bfr_after (
		.din(_0456_),
		.dout(new_net_7199)
	);

	bfr new_net_2318_bfr_after (
		.din(new_net_7199),
		.dout(new_net_2318)
	);

	bfr new_net_7200_bfr_after (
		.din(_1008_),
		.dout(new_net_7200)
	);

	bfr new_net_7201_bfr_after (
		.din(new_net_7200),
		.dout(new_net_7201)
	);

	bfr new_net_7202_bfr_after (
		.din(new_net_7201),
		.dout(new_net_7202)
	);

	bfr new_net_7203_bfr_after (
		.din(new_net_7202),
		.dout(new_net_7203)
	);

	bfr new_net_7204_bfr_after (
		.din(new_net_7203),
		.dout(new_net_7204)
	);

	bfr new_net_7205_bfr_after (
		.din(new_net_7204),
		.dout(new_net_7205)
	);

	bfr new_net_7206_bfr_after (
		.din(new_net_7205),
		.dout(new_net_7206)
	);

	bfr new_net_7207_bfr_after (
		.din(new_net_7206),
		.dout(new_net_7207)
	);

	bfr new_net_7208_bfr_after (
		.din(new_net_7207),
		.dout(new_net_7208)
	);

	bfr new_net_7209_bfr_after (
		.din(new_net_7208),
		.dout(new_net_7209)
	);

	bfr new_net_7210_bfr_after (
		.din(new_net_7209),
		.dout(new_net_7210)
	);

	bfr new_net_7211_bfr_after (
		.din(new_net_7210),
		.dout(new_net_7211)
	);

	bfr new_net_7212_bfr_after (
		.din(new_net_7211),
		.dout(new_net_7212)
	);

	bfr new_net_7213_bfr_after (
		.din(new_net_7212),
		.dout(new_net_7213)
	);

	bfr new_net_7214_bfr_after (
		.din(new_net_7213),
		.dout(new_net_7214)
	);

	bfr new_net_7215_bfr_after (
		.din(new_net_7214),
		.dout(new_net_7215)
	);

	bfr new_net_7216_bfr_after (
		.din(new_net_7215),
		.dout(new_net_7216)
	);

	bfr new_net_7217_bfr_after (
		.din(new_net_7216),
		.dout(new_net_7217)
	);

	bfr new_net_7218_bfr_after (
		.din(new_net_7217),
		.dout(new_net_7218)
	);

	bfr new_net_7219_bfr_after (
		.din(new_net_7218),
		.dout(new_net_7219)
	);

	bfr new_net_7220_bfr_after (
		.din(new_net_7219),
		.dout(new_net_7220)
	);

	bfr new_net_7221_bfr_after (
		.din(new_net_7220),
		.dout(new_net_7221)
	);

	bfr new_net_7222_bfr_after (
		.din(new_net_7221),
		.dout(new_net_7222)
	);

	bfr new_net_7223_bfr_after (
		.din(new_net_7222),
		.dout(new_net_7223)
	);

	bfr new_net_7224_bfr_after (
		.din(new_net_7223),
		.dout(new_net_7224)
	);

	bfr new_net_2198_bfr_after (
		.din(new_net_7224),
		.dout(new_net_2198)
	);

	bfr new_net_7225_bfr_after (
		.din(_0345_),
		.dout(new_net_7225)
	);

	bfr new_net_7226_bfr_after (
		.din(new_net_7225),
		.dout(new_net_7226)
	);

	bfr new_net_2290_bfr_after (
		.din(new_net_7226),
		.dout(new_net_2290)
	);

	bfr new_net_7227_bfr_after (
		.din(new_net_2433),
		.dout(new_net_7227)
	);

	bfr new_net_7228_bfr_after (
		.din(new_net_7227),
		.dout(new_net_7228)
	);

	bfr new_net_7229_bfr_after (
		.din(new_net_7228),
		.dout(new_net_7229)
	);

	bfr new_net_7230_bfr_after (
		.din(new_net_7229),
		.dout(new_net_7230)
	);

	bfr new_net_7231_bfr_after (
		.din(new_net_7230),
		.dout(new_net_7231)
	);

	bfr new_net_7232_bfr_after (
		.din(new_net_7231),
		.dout(new_net_7232)
	);

	bfr new_net_7233_bfr_after (
		.din(new_net_7232),
		.dout(new_net_7233)
	);

	bfr new_net_7234_bfr_after (
		.din(new_net_7233),
		.dout(new_net_7234)
	);

	bfr new_net_7235_bfr_after (
		.din(new_net_7234),
		.dout(new_net_7235)
	);

	bfr new_net_7236_bfr_after (
		.din(new_net_7235),
		.dout(new_net_7236)
	);

	bfr new_net_7237_bfr_after (
		.din(new_net_7236),
		.dout(new_net_7237)
	);

	bfr new_net_7238_bfr_after (
		.din(new_net_7237),
		.dout(new_net_7238)
	);

	bfr new_net_7239_bfr_after (
		.din(new_net_7238),
		.dout(new_net_7239)
	);

	bfr new_net_7240_bfr_after (
		.din(new_net_7239),
		.dout(new_net_7240)
	);

	bfr new_net_7241_bfr_after (
		.din(new_net_7240),
		.dout(new_net_7241)
	);

	bfr new_net_7242_bfr_after (
		.din(new_net_7241),
		.dout(new_net_7242)
	);

	bfr new_net_7243_bfr_after (
		.din(new_net_7242),
		.dout(new_net_7243)
	);

	bfr new_net_7244_bfr_after (
		.din(new_net_7243),
		.dout(new_net_7244)
	);

	bfr new_net_7245_bfr_after (
		.din(new_net_7244),
		.dout(new_net_7245)
	);

	bfr new_net_7246_bfr_after (
		.din(new_net_7245),
		.dout(new_net_7246)
	);

	bfr new_net_7247_bfr_after (
		.din(new_net_7246),
		.dout(new_net_7247)
	);

	bfr new_net_7248_bfr_after (
		.din(new_net_7247),
		.dout(new_net_7248)
	);

	bfr new_net_7249_bfr_after (
		.din(new_net_7248),
		.dout(new_net_7249)
	);

	bfr G5240_bfr_after (
		.din(new_net_7249),
		.dout(G5240)
	);

	bfr new_net_7250_bfr_after (
		.din(new_net_2447),
		.dout(new_net_7250)
	);

	bfr new_net_7251_bfr_after (
		.din(new_net_7250),
		.dout(new_net_7251)
	);

	bfr new_net_7252_bfr_after (
		.din(new_net_7251),
		.dout(new_net_7252)
	);

	bfr new_net_7253_bfr_after (
		.din(new_net_7252),
		.dout(new_net_7253)
	);

	bfr new_net_7254_bfr_after (
		.din(new_net_7253),
		.dout(new_net_7254)
	);

	bfr new_net_7255_bfr_after (
		.din(new_net_7254),
		.dout(new_net_7255)
	);

	bfr new_net_7256_bfr_after (
		.din(new_net_7255),
		.dout(new_net_7256)
	);

	bfr new_net_7257_bfr_after (
		.din(new_net_7256),
		.dout(new_net_7257)
	);

	bfr new_net_7258_bfr_after (
		.din(new_net_7257),
		.dout(new_net_7258)
	);

	bfr new_net_7259_bfr_after (
		.din(new_net_7258),
		.dout(new_net_7259)
	);

	bfr new_net_7260_bfr_after (
		.din(new_net_7259),
		.dout(new_net_7260)
	);

	bfr new_net_7261_bfr_after (
		.din(new_net_7260),
		.dout(new_net_7261)
	);

	bfr new_net_7262_bfr_after (
		.din(new_net_7261),
		.dout(new_net_7262)
	);

	bfr new_net_7263_bfr_after (
		.din(new_net_7262),
		.dout(new_net_7263)
	);

	bfr new_net_7264_bfr_after (
		.din(new_net_7263),
		.dout(new_net_7264)
	);

	bfr new_net_7265_bfr_after (
		.din(new_net_7264),
		.dout(new_net_7265)
	);

	bfr new_net_7266_bfr_after (
		.din(new_net_7265),
		.dout(new_net_7266)
	);

	bfr new_net_7267_bfr_after (
		.din(new_net_7266),
		.dout(new_net_7267)
	);

	bfr new_net_7268_bfr_after (
		.din(new_net_7267),
		.dout(new_net_7268)
	);

	bfr new_net_7269_bfr_after (
		.din(new_net_7268),
		.dout(new_net_7269)
	);

	bfr new_net_7270_bfr_after (
		.din(new_net_7269),
		.dout(new_net_7270)
	);

	bfr new_net_7271_bfr_after (
		.din(new_net_7270),
		.dout(new_net_7271)
	);

	bfr new_net_7272_bfr_after (
		.din(new_net_7271),
		.dout(new_net_7272)
	);

	bfr new_net_7273_bfr_after (
		.din(new_net_7272),
		.dout(new_net_7273)
	);

	bfr new_net_7274_bfr_after (
		.din(new_net_7273),
		.dout(new_net_7274)
	);

	bfr new_net_7275_bfr_after (
		.din(new_net_7274),
		.dout(new_net_7275)
	);

	bfr new_net_7276_bfr_after (
		.din(new_net_7275),
		.dout(new_net_7276)
	);

	bfr new_net_7277_bfr_after (
		.din(new_net_7276),
		.dout(new_net_7277)
	);

	bfr new_net_7278_bfr_after (
		.din(new_net_7277),
		.dout(new_net_7278)
	);

	bfr G5236_bfr_after (
		.din(new_net_7278),
		.dout(G5236)
	);

	bfr new_net_7279_bfr_after (
		.din(new_net_2459),
		.dout(new_net_7279)
	);

	bfr new_net_7280_bfr_after (
		.din(new_net_7279),
		.dout(new_net_7280)
	);

	bfr new_net_7281_bfr_after (
		.din(new_net_7280),
		.dout(new_net_7281)
	);

	bfr new_net_7282_bfr_after (
		.din(new_net_7281),
		.dout(new_net_7282)
	);

	bfr new_net_7283_bfr_after (
		.din(new_net_7282),
		.dout(new_net_7283)
	);

	bfr new_net_7284_bfr_after (
		.din(new_net_7283),
		.dout(new_net_7284)
	);

	bfr new_net_7285_bfr_after (
		.din(new_net_7284),
		.dout(new_net_7285)
	);

	bfr new_net_7286_bfr_after (
		.din(new_net_7285),
		.dout(new_net_7286)
	);

	bfr new_net_7287_bfr_after (
		.din(new_net_7286),
		.dout(new_net_7287)
	);

	bfr new_net_7288_bfr_after (
		.din(new_net_7287),
		.dout(new_net_7288)
	);

	bfr new_net_7289_bfr_after (
		.din(new_net_7288),
		.dout(new_net_7289)
	);

	bfr new_net_7290_bfr_after (
		.din(new_net_7289),
		.dout(new_net_7290)
	);

	bfr new_net_7291_bfr_after (
		.din(new_net_7290),
		.dout(new_net_7291)
	);

	bfr new_net_7292_bfr_after (
		.din(new_net_7291),
		.dout(new_net_7292)
	);

	bfr new_net_7293_bfr_after (
		.din(new_net_7292),
		.dout(new_net_7293)
	);

	bfr new_net_7294_bfr_after (
		.din(new_net_7293),
		.dout(new_net_7294)
	);

	bfr new_net_7295_bfr_after (
		.din(new_net_7294),
		.dout(new_net_7295)
	);

	bfr new_net_7296_bfr_after (
		.din(new_net_7295),
		.dout(new_net_7296)
	);

	bfr new_net_7297_bfr_after (
		.din(new_net_7296),
		.dout(new_net_7297)
	);

	bfr new_net_7298_bfr_after (
		.din(new_net_7297),
		.dout(new_net_7298)
	);

	bfr new_net_7299_bfr_after (
		.din(new_net_7298),
		.dout(new_net_7299)
	);

	bfr new_net_7300_bfr_after (
		.din(new_net_7299),
		.dout(new_net_7300)
	);

	bfr new_net_7301_bfr_after (
		.din(new_net_7300),
		.dout(new_net_7301)
	);

	bfr new_net_7302_bfr_after (
		.din(new_net_7301),
		.dout(new_net_7302)
	);

	bfr new_net_7303_bfr_after (
		.din(new_net_7302),
		.dout(new_net_7303)
	);

	bfr new_net_7304_bfr_after (
		.din(new_net_7303),
		.dout(new_net_7304)
	);

	bfr new_net_7305_bfr_after (
		.din(new_net_7304),
		.dout(new_net_7305)
	);

	bfr new_net_7306_bfr_after (
		.din(new_net_7305),
		.dout(new_net_7306)
	);

	bfr new_net_7307_bfr_after (
		.din(new_net_7306),
		.dout(new_net_7307)
	);

	bfr new_net_7308_bfr_after (
		.din(new_net_7307),
		.dout(new_net_7308)
	);

	bfr new_net_7309_bfr_after (
		.din(new_net_7308),
		.dout(new_net_7309)
	);

	bfr new_net_7310_bfr_after (
		.din(new_net_7309),
		.dout(new_net_7310)
	);

	bfr new_net_7311_bfr_after (
		.din(new_net_7310),
		.dout(new_net_7311)
	);

	bfr new_net_7312_bfr_after (
		.din(new_net_7311),
		.dout(new_net_7312)
	);

	bfr G5234_bfr_after (
		.din(new_net_7312),
		.dout(G5234)
	);

	bfr new_net_7313_bfr_after (
		.din(new_net_2471),
		.dout(new_net_7313)
	);

	bfr new_net_7314_bfr_after (
		.din(new_net_7313),
		.dout(new_net_7314)
	);

	bfr new_net_7315_bfr_after (
		.din(new_net_7314),
		.dout(new_net_7315)
	);

	bfr new_net_7316_bfr_after (
		.din(new_net_7315),
		.dout(new_net_7316)
	);

	bfr new_net_7317_bfr_after (
		.din(new_net_7316),
		.dout(new_net_7317)
	);

	bfr new_net_7318_bfr_after (
		.din(new_net_7317),
		.dout(new_net_7318)
	);

	bfr new_net_7319_bfr_after (
		.din(new_net_7318),
		.dout(new_net_7319)
	);

	bfr new_net_7320_bfr_after (
		.din(new_net_7319),
		.dout(new_net_7320)
	);

	bfr new_net_7321_bfr_after (
		.din(new_net_7320),
		.dout(new_net_7321)
	);

	bfr new_net_7322_bfr_after (
		.din(new_net_7321),
		.dout(new_net_7322)
	);

	bfr G5282_bfr_after (
		.din(new_net_7322),
		.dout(G5282)
	);

	bfr new_net_7323_bfr_after (
		.din(new_net_2483),
		.dout(new_net_7323)
	);

	bfr new_net_7324_bfr_after (
		.din(new_net_7323),
		.dout(new_net_7324)
	);

	bfr new_net_7325_bfr_after (
		.din(new_net_7324),
		.dout(new_net_7325)
	);

	bfr new_net_7326_bfr_after (
		.din(new_net_7325),
		.dout(new_net_7326)
	);

	bfr new_net_7327_bfr_after (
		.din(new_net_7326),
		.dout(new_net_7327)
	);

	bfr G5298_bfr_after (
		.din(new_net_7327),
		.dout(G5298)
	);

	bfr new_net_7328_bfr_after (
		.din(new_net_2495),
		.dout(new_net_7328)
	);

	bfr new_net_7329_bfr_after (
		.din(new_net_7328),
		.dout(new_net_7329)
	);

	bfr new_net_7330_bfr_after (
		.din(new_net_7329),
		.dout(new_net_7330)
	);

	bfr new_net_7331_bfr_after (
		.din(new_net_7330),
		.dout(new_net_7331)
	);

	bfr new_net_7332_bfr_after (
		.din(new_net_7331),
		.dout(new_net_7332)
	);

	bfr new_net_7333_bfr_after (
		.din(new_net_7332),
		.dout(new_net_7333)
	);

	bfr new_net_7334_bfr_after (
		.din(new_net_7333),
		.dout(new_net_7334)
	);

	bfr new_net_7335_bfr_after (
		.din(new_net_7334),
		.dout(new_net_7335)
	);

	bfr new_net_7336_bfr_after (
		.din(new_net_7335),
		.dout(new_net_7336)
	);

	bfr new_net_7337_bfr_after (
		.din(new_net_7336),
		.dout(new_net_7337)
	);

	bfr new_net_7338_bfr_after (
		.din(new_net_7337),
		.dout(new_net_7338)
	);

	bfr new_net_7339_bfr_after (
		.din(new_net_7338),
		.dout(new_net_7339)
	);

	bfr new_net_7340_bfr_after (
		.din(new_net_7339),
		.dout(new_net_7340)
	);

	bfr new_net_7341_bfr_after (
		.din(new_net_7340),
		.dout(new_net_7341)
	);

	bfr new_net_7342_bfr_after (
		.din(new_net_7341),
		.dout(new_net_7342)
	);

	bfr new_net_7343_bfr_after (
		.din(new_net_7342),
		.dout(new_net_7343)
	);

	bfr new_net_7344_bfr_after (
		.din(new_net_7343),
		.dout(new_net_7344)
	);

	bfr new_net_7345_bfr_after (
		.din(new_net_7344),
		.dout(new_net_7345)
	);

	bfr new_net_7346_bfr_after (
		.din(new_net_7345),
		.dout(new_net_7346)
	);

	bfr new_net_7347_bfr_after (
		.din(new_net_7346),
		.dout(new_net_7347)
	);

	bfr new_net_7348_bfr_after (
		.din(new_net_7347),
		.dout(new_net_7348)
	);

	bfr new_net_7349_bfr_after (
		.din(new_net_7348),
		.dout(new_net_7349)
	);

	bfr new_net_7350_bfr_after (
		.din(new_net_7349),
		.dout(new_net_7350)
	);

	bfr new_net_7351_bfr_after (
		.din(new_net_7350),
		.dout(new_net_7351)
	);

	bfr new_net_7352_bfr_after (
		.din(new_net_7351),
		.dout(new_net_7352)
	);

	bfr new_net_7353_bfr_after (
		.din(new_net_7352),
		.dout(new_net_7353)
	);

	bfr new_net_7354_bfr_after (
		.din(new_net_7353),
		.dout(new_net_7354)
	);

	bfr new_net_7355_bfr_after (
		.din(new_net_7354),
		.dout(new_net_7355)
	);

	bfr new_net_7356_bfr_after (
		.din(new_net_7355),
		.dout(new_net_7356)
	);

	bfr new_net_7357_bfr_after (
		.din(new_net_7356),
		.dout(new_net_7357)
	);

	bfr new_net_7358_bfr_after (
		.din(new_net_7357),
		.dout(new_net_7358)
	);

	bfr new_net_7359_bfr_after (
		.din(new_net_7358),
		.dout(new_net_7359)
	);

	bfr new_net_7360_bfr_after (
		.din(new_net_7359),
		.dout(new_net_7360)
	);

	bfr new_net_7361_bfr_after (
		.din(new_net_7360),
		.dout(new_net_7361)
	);

	bfr new_net_7362_bfr_after (
		.din(new_net_7361),
		.dout(new_net_7362)
	);

	bfr new_net_7363_bfr_after (
		.din(new_net_7362),
		.dout(new_net_7363)
	);

	bfr G5231_bfr_after (
		.din(new_net_7363),
		.dout(G5231)
	);

	bfr new_net_7364_bfr_after (
		.din(new_net_2507),
		.dout(new_net_7364)
	);

	bfr new_net_7365_bfr_after (
		.din(new_net_7364),
		.dout(new_net_7365)
	);

	bfr new_net_7366_bfr_after (
		.din(new_net_7365),
		.dout(new_net_7366)
	);

	bfr new_net_7367_bfr_after (
		.din(new_net_7366),
		.dout(new_net_7367)
	);

	bfr new_net_7368_bfr_after (
		.din(new_net_7367),
		.dout(new_net_7368)
	);

	bfr new_net_7369_bfr_after (
		.din(new_net_7368),
		.dout(new_net_7369)
	);

	bfr new_net_7370_bfr_after (
		.din(new_net_7369),
		.dout(new_net_7370)
	);

	bfr new_net_7371_bfr_after (
		.din(new_net_7370),
		.dout(new_net_7371)
	);

	bfr new_net_7372_bfr_after (
		.din(new_net_7371),
		.dout(new_net_7372)
	);

	bfr new_net_7373_bfr_after (
		.din(new_net_7372),
		.dout(new_net_7373)
	);

	bfr new_net_7374_bfr_after (
		.din(new_net_7373),
		.dout(new_net_7374)
	);

	bfr new_net_7375_bfr_after (
		.din(new_net_7374),
		.dout(new_net_7375)
	);

	bfr new_net_7376_bfr_after (
		.din(new_net_7375),
		.dout(new_net_7376)
	);

	bfr new_net_7377_bfr_after (
		.din(new_net_7376),
		.dout(new_net_7377)
	);

	bfr new_net_7378_bfr_after (
		.din(new_net_7377),
		.dout(new_net_7378)
	);

	bfr new_net_7379_bfr_after (
		.din(new_net_7378),
		.dout(new_net_7379)
	);

	bfr new_net_7380_bfr_after (
		.din(new_net_7379),
		.dout(new_net_7380)
	);

	bfr new_net_7381_bfr_after (
		.din(new_net_7380),
		.dout(new_net_7381)
	);

	bfr new_net_7382_bfr_after (
		.din(new_net_7381),
		.dout(new_net_7382)
	);

	bfr new_net_7383_bfr_after (
		.din(new_net_7382),
		.dout(new_net_7383)
	);

	bfr new_net_7384_bfr_after (
		.din(new_net_7383),
		.dout(new_net_7384)
	);

	bfr new_net_7385_bfr_after (
		.din(new_net_7384),
		.dout(new_net_7385)
	);

	bfr new_net_7386_bfr_after (
		.din(new_net_7385),
		.dout(new_net_7386)
	);

	bfr new_net_7387_bfr_after (
		.din(new_net_7386),
		.dout(new_net_7387)
	);

	bfr new_net_7388_bfr_after (
		.din(new_net_7387),
		.dout(new_net_7388)
	);

	bfr new_net_7389_bfr_after (
		.din(new_net_7388),
		.dout(new_net_7389)
	);

	bfr new_net_7390_bfr_after (
		.din(new_net_7389),
		.dout(new_net_7390)
	);

	bfr new_net_7391_bfr_after (
		.din(new_net_7390),
		.dout(new_net_7391)
	);

	bfr new_net_7392_bfr_after (
		.din(new_net_7391),
		.dout(new_net_7392)
	);

	bfr new_net_7393_bfr_after (
		.din(new_net_7392),
		.dout(new_net_7393)
	);

	bfr new_net_7394_bfr_after (
		.din(new_net_7393),
		.dout(new_net_7394)
	);

	bfr new_net_7395_bfr_after (
		.din(new_net_7394),
		.dout(new_net_7395)
	);

	bfr new_net_7396_bfr_after (
		.din(new_net_7395),
		.dout(new_net_7396)
	);

	bfr new_net_7397_bfr_after (
		.din(new_net_7396),
		.dout(new_net_7397)
	);

	bfr new_net_7398_bfr_after (
		.din(new_net_7397),
		.dout(new_net_7398)
	);

	bfr G5228_bfr_after (
		.din(new_net_7398),
		.dout(G5228)
	);

	bfr new_net_7399_bfr_after (
		.din(_0328_),
		.dout(new_net_7399)
	);

	bfr new_net_7400_bfr_after (
		.din(new_net_7399),
		.dout(new_net_7400)
	);

	bfr new_net_7401_bfr_after (
		.din(new_net_7400),
		.dout(new_net_7401)
	);

	bfr new_net_7402_bfr_after (
		.din(new_net_7401),
		.dout(new_net_7402)
	);

	bfr new_net_7403_bfr_after (
		.din(new_net_7402),
		.dout(new_net_7403)
	);

	bfr new_net_7404_bfr_after (
		.din(new_net_7403),
		.dout(new_net_7404)
	);

	bfr new_net_7405_bfr_after (
		.din(new_net_7404),
		.dout(new_net_7405)
	);

	bfr new_net_7406_bfr_after (
		.din(new_net_7405),
		.dout(new_net_7406)
	);

	bfr new_net_7407_bfr_after (
		.din(new_net_7406),
		.dout(new_net_7407)
	);

	bfr new_net_7408_bfr_after (
		.din(new_net_7407),
		.dout(new_net_7408)
	);

	bfr new_net_7409_bfr_after (
		.din(new_net_7408),
		.dout(new_net_7409)
	);

	bfr new_net_7410_bfr_after (
		.din(new_net_7409),
		.dout(new_net_7410)
	);

	bfr new_net_7411_bfr_after (
		.din(new_net_7410),
		.dout(new_net_7411)
	);

	bfr new_net_7412_bfr_after (
		.din(new_net_7411),
		.dout(new_net_7412)
	);

	bfr new_net_7413_bfr_after (
		.din(new_net_7412),
		.dout(new_net_7413)
	);

	bfr new_net_7414_bfr_after (
		.din(new_net_7413),
		.dout(new_net_7414)
	);

	bfr new_net_7415_bfr_after (
		.din(new_net_7414),
		.dout(new_net_7415)
	);

	bfr new_net_7416_bfr_after (
		.din(new_net_7415),
		.dout(new_net_7416)
	);

	bfr new_net_2286_bfr_after (
		.din(new_net_7416),
		.dout(new_net_2286)
	);

	bfr new_net_7417_bfr_after (
		.din(_0084_),
		.dout(new_net_7417)
	);

	bfr new_net_7418_bfr_after (
		.din(new_net_7417),
		.dout(new_net_7418)
	);

	bfr new_net_7419_bfr_after (
		.din(new_net_7418),
		.dout(new_net_7419)
	);

	bfr new_net_7420_bfr_after (
		.din(new_net_7419),
		.dout(new_net_7420)
	);

	bfr new_net_7421_bfr_after (
		.din(new_net_7420),
		.dout(new_net_7421)
	);

	bfr new_net_7422_bfr_after (
		.din(new_net_7421),
		.dout(new_net_7422)
	);

	bfr new_net_7423_bfr_after (
		.din(new_net_7422),
		.dout(new_net_7423)
	);

	bfr new_net_7424_bfr_after (
		.din(new_net_7423),
		.dout(new_net_7424)
	);

	bfr new_net_7425_bfr_after (
		.din(new_net_7424),
		.dout(new_net_7425)
	);

	bfr new_net_2229_bfr_after (
		.din(new_net_7425),
		.dout(new_net_2229)
	);

	bfr new_net_7426_bfr_after (
		.din(new_net_2367),
		.dout(new_net_7426)
	);

	bfr new_net_7427_bfr_after (
		.din(new_net_7426),
		.dout(new_net_7427)
	);

	bfr new_net_7428_bfr_after (
		.din(new_net_7427),
		.dout(new_net_7428)
	);

	bfr new_net_7429_bfr_after (
		.din(new_net_7428),
		.dout(new_net_7429)
	);

	bfr new_net_7430_bfr_after (
		.din(new_net_7429),
		.dout(new_net_7430)
	);

	bfr new_net_7431_bfr_after (
		.din(new_net_7430),
		.dout(new_net_7431)
	);

	bfr new_net_7432_bfr_after (
		.din(new_net_7431),
		.dout(new_net_7432)
	);

	bfr new_net_7433_bfr_after (
		.din(new_net_7432),
		.dout(new_net_7433)
	);

	bfr new_net_7434_bfr_after (
		.din(new_net_7433),
		.dout(new_net_7434)
	);

	bfr new_net_7435_bfr_after (
		.din(new_net_7434),
		.dout(new_net_7435)
	);

	bfr new_net_7436_bfr_after (
		.din(new_net_7435),
		.dout(new_net_7436)
	);

	bfr new_net_7437_bfr_after (
		.din(new_net_7436),
		.dout(new_net_7437)
	);

	bfr new_net_7438_bfr_after (
		.din(new_net_7437),
		.dout(new_net_7438)
	);

	bfr new_net_7439_bfr_after (
		.din(new_net_7438),
		.dout(new_net_7439)
	);

	bfr new_net_7440_bfr_after (
		.din(new_net_7439),
		.dout(new_net_7440)
	);

	bfr new_net_7441_bfr_after (
		.din(new_net_7440),
		.dout(new_net_7441)
	);

	bfr new_net_7442_bfr_after (
		.din(new_net_7441),
		.dout(new_net_7442)
	);

	bfr new_net_7443_bfr_after (
		.din(new_net_7442),
		.dout(new_net_7443)
	);

	bfr new_net_7444_bfr_after (
		.din(new_net_7443),
		.dout(new_net_7444)
	);

	bfr new_net_7445_bfr_after (
		.din(new_net_7444),
		.dout(new_net_7445)
	);

	bfr new_net_7446_bfr_after (
		.din(new_net_7445),
		.dout(new_net_7446)
	);

	bfr new_net_7447_bfr_after (
		.din(new_net_7446),
		.dout(new_net_7447)
	);

	bfr new_net_7448_bfr_after (
		.din(new_net_7447),
		.dout(new_net_7448)
	);

	bfr new_net_7449_bfr_after (
		.din(new_net_7448),
		.dout(new_net_7449)
	);

	bfr new_net_7450_bfr_after (
		.din(new_net_7449),
		.dout(new_net_7450)
	);

	bfr new_net_7451_bfr_after (
		.din(new_net_7450),
		.dout(new_net_7451)
	);

	bfr new_net_7452_bfr_after (
		.din(new_net_7451),
		.dout(new_net_7452)
	);

	bfr new_net_7453_bfr_after (
		.din(new_net_7452),
		.dout(new_net_7453)
	);

	bfr new_net_7454_bfr_after (
		.din(new_net_7453),
		.dout(new_net_7454)
	);

	bfr new_net_7455_bfr_after (
		.din(new_net_7454),
		.dout(new_net_7455)
	);

	bfr new_net_7456_bfr_after (
		.din(new_net_7455),
		.dout(new_net_7456)
	);

	bfr new_net_7457_bfr_after (
		.din(new_net_7456),
		.dout(new_net_7457)
	);

	bfr new_net_7458_bfr_after (
		.din(new_net_7457),
		.dout(new_net_7458)
	);

	bfr new_net_7459_bfr_after (
		.din(new_net_7458),
		.dout(new_net_7459)
	);

	bfr new_net_7460_bfr_after (
		.din(new_net_7459),
		.dout(new_net_7460)
	);

	bfr new_net_7461_bfr_after (
		.din(new_net_7460),
		.dout(new_net_7461)
	);

	bfr new_net_7462_bfr_after (
		.din(new_net_7461),
		.dout(new_net_7462)
	);

	bfr new_net_7463_bfr_after (
		.din(new_net_7462),
		.dout(new_net_7463)
	);

	bfr new_net_7464_bfr_after (
		.din(new_net_7463),
		.dout(new_net_7464)
	);

	bfr G5205_bfr_after (
		.din(new_net_7464),
		.dout(G5205)
	);

	bfr new_net_2281_bfr_after (
		.din(_0310_),
		.dout(new_net_2281)
	);

	bfr new_net_7465_bfr_after (
		.din(_0563_),
		.dout(new_net_7465)
	);

	bfr new_net_7466_bfr_after (
		.din(new_net_7465),
		.dout(new_net_7466)
	);

	bfr new_net_7467_bfr_after (
		.din(new_net_7466),
		.dout(new_net_7467)
	);

	bfr new_net_7468_bfr_after (
		.din(new_net_7467),
		.dout(new_net_7468)
	);

	bfr new_net_7469_bfr_after (
		.din(new_net_7468),
		.dout(new_net_7469)
	);

	bfr new_net_7470_bfr_after (
		.din(new_net_7469),
		.dout(new_net_7470)
	);

	bfr new_net_7471_bfr_after (
		.din(new_net_7470),
		.dout(new_net_7471)
	);

	bfr new_net_7472_bfr_after (
		.din(new_net_7471),
		.dout(new_net_7472)
	);

	bfr new_net_7473_bfr_after (
		.din(new_net_7472),
		.dout(new_net_7473)
	);

	bfr new_net_7474_bfr_after (
		.din(new_net_7473),
		.dout(new_net_7474)
	);

	bfr new_net_7475_bfr_after (
		.din(new_net_7474),
		.dout(new_net_7475)
	);

	bfr new_net_7476_bfr_after (
		.din(new_net_7475),
		.dout(new_net_7476)
	);

	bfr new_net_7477_bfr_after (
		.din(new_net_7476),
		.dout(new_net_7477)
	);

	bfr new_net_7478_bfr_after (
		.din(new_net_7477),
		.dout(new_net_7478)
	);

	bfr new_net_7479_bfr_after (
		.din(new_net_7478),
		.dout(new_net_7479)
	);

	bfr new_net_7480_bfr_after (
		.din(new_net_7479),
		.dout(new_net_7480)
	);

	bfr new_net_7481_bfr_after (
		.din(new_net_7480),
		.dout(new_net_7481)
	);

	bfr new_net_7482_bfr_after (
		.din(new_net_7481),
		.dout(new_net_7482)
	);

	bfr new_net_7483_bfr_after (
		.din(new_net_7482),
		.dout(new_net_7483)
	);

	bfr new_net_7484_bfr_after (
		.din(new_net_7483),
		.dout(new_net_7484)
	);

	bfr new_net_7485_bfr_after (
		.din(new_net_7484),
		.dout(new_net_7485)
	);

	bfr new_net_7486_bfr_after (
		.din(new_net_7485),
		.dout(new_net_7486)
	);

	bfr new_net_7487_bfr_after (
		.din(new_net_7486),
		.dout(new_net_7487)
	);

	bfr new_net_7488_bfr_after (
		.din(new_net_7487),
		.dout(new_net_7488)
	);

	bfr new_net_7489_bfr_after (
		.din(new_net_7488),
		.dout(new_net_7489)
	);

	bfr new_net_7490_bfr_after (
		.din(new_net_7489),
		.dout(new_net_7490)
	);

	bfr new_net_7491_bfr_after (
		.din(new_net_7490),
		.dout(new_net_7491)
	);

	bfr new_net_7492_bfr_after (
		.din(new_net_7491),
		.dout(new_net_7492)
	);

	bfr new_net_2344_bfr_after (
		.din(new_net_7492),
		.dout(new_net_2344)
	);

	bfr new_net_2218_bfr_after (
		.din(_1232_),
		.dout(new_net_2218)
	);

	bfr new_net_7493_bfr_after (
		.din(_0399_),
		.dout(new_net_7493)
	);

	bfr new_net_2302_bfr_after (
		.din(new_net_7493),
		.dout(new_net_2302)
	);

	bfr new_net_7494_bfr_after (
		.din(new_net_2441),
		.dout(new_net_7494)
	);

	bfr new_net_7495_bfr_after (
		.din(new_net_7494),
		.dout(new_net_7495)
	);

	bfr new_net_7496_bfr_after (
		.din(new_net_7495),
		.dout(new_net_7496)
	);

	bfr new_net_7497_bfr_after (
		.din(new_net_7496),
		.dout(new_net_7497)
	);

	bfr new_net_7498_bfr_after (
		.din(new_net_7497),
		.dout(new_net_7498)
	);

	bfr new_net_7499_bfr_after (
		.din(new_net_7498),
		.dout(new_net_7499)
	);

	bfr new_net_7500_bfr_after (
		.din(new_net_7499),
		.dout(new_net_7500)
	);

	bfr new_net_7501_bfr_after (
		.din(new_net_7500),
		.dout(new_net_7501)
	);

	bfr new_net_7502_bfr_after (
		.din(new_net_7501),
		.dout(new_net_7502)
	);

	bfr new_net_7503_bfr_after (
		.din(new_net_7502),
		.dout(new_net_7503)
	);

	bfr new_net_7504_bfr_after (
		.din(new_net_7503),
		.dout(new_net_7504)
	);

	bfr new_net_7505_bfr_after (
		.din(new_net_7504),
		.dout(new_net_7505)
	);

	bfr new_net_7506_bfr_after (
		.din(new_net_7505),
		.dout(new_net_7506)
	);

	bfr new_net_7507_bfr_after (
		.din(new_net_7506),
		.dout(new_net_7507)
	);

	bfr new_net_7508_bfr_after (
		.din(new_net_7507),
		.dout(new_net_7508)
	);

	bfr new_net_7509_bfr_after (
		.din(new_net_7508),
		.dout(new_net_7509)
	);

	bfr new_net_7510_bfr_after (
		.din(new_net_7509),
		.dout(new_net_7510)
	);

	bfr new_net_7511_bfr_after (
		.din(new_net_7510),
		.dout(new_net_7511)
	);

	bfr new_net_7512_bfr_after (
		.din(new_net_7511),
		.dout(new_net_7512)
	);

	bfr new_net_7513_bfr_after (
		.din(new_net_7512),
		.dout(new_net_7513)
	);

	bfr new_net_7514_bfr_after (
		.din(new_net_7513),
		.dout(new_net_7514)
	);

	bfr new_net_7515_bfr_after (
		.din(new_net_7514),
		.dout(new_net_7515)
	);

	bfr new_net_7516_bfr_after (
		.din(new_net_7515),
		.dout(new_net_7516)
	);

	bfr new_net_7517_bfr_after (
		.din(new_net_7516),
		.dout(new_net_7517)
	);

	bfr new_net_7518_bfr_after (
		.din(new_net_7517),
		.dout(new_net_7518)
	);

	bfr new_net_7519_bfr_after (
		.din(new_net_7518),
		.dout(new_net_7519)
	);

	bfr new_net_7520_bfr_after (
		.din(new_net_7519),
		.dout(new_net_7520)
	);

	bfr new_net_7521_bfr_after (
		.din(new_net_7520),
		.dout(new_net_7521)
	);

	bfr new_net_7522_bfr_after (
		.din(new_net_7521),
		.dout(new_net_7522)
	);

	bfr new_net_7523_bfr_after (
		.din(new_net_7522),
		.dout(new_net_7523)
	);

	bfr new_net_7524_bfr_after (
		.din(new_net_7523),
		.dout(new_net_7524)
	);

	bfr new_net_7525_bfr_after (
		.din(new_net_7524),
		.dout(new_net_7525)
	);

	bfr new_net_7526_bfr_after (
		.din(new_net_7525),
		.dout(new_net_7526)
	);

	bfr new_net_7527_bfr_after (
		.din(new_net_7526),
		.dout(new_net_7527)
	);

	bfr new_net_7528_bfr_after (
		.din(new_net_7527),
		.dout(new_net_7528)
	);

	bfr new_net_7529_bfr_after (
		.din(new_net_7528),
		.dout(new_net_7529)
	);

	bfr new_net_7530_bfr_after (
		.din(new_net_7529),
		.dout(new_net_7530)
	);

	bfr new_net_7531_bfr_after (
		.din(new_net_7530),
		.dout(new_net_7531)
	);

	bfr new_net_7532_bfr_after (
		.din(new_net_7531),
		.dout(new_net_7532)
	);

	bfr G5206_bfr_after (
		.din(new_net_7532),
		.dout(G5206)
	);

	bfr G5314_bfr_after (
		.din(new_net_2453),
		.dout(G5314)
	);

	bfr new_net_7533_bfr_after (
		.din(new_net_2477),
		.dout(new_net_7533)
	);

	bfr new_net_7534_bfr_after (
		.din(new_net_7533),
		.dout(new_net_7534)
	);

	bfr new_net_7535_bfr_after (
		.din(new_net_7534),
		.dout(new_net_7535)
	);

	bfr new_net_7536_bfr_after (
		.din(new_net_7535),
		.dout(new_net_7536)
	);

	bfr new_net_7537_bfr_after (
		.din(new_net_7536),
		.dout(new_net_7537)
	);

	bfr new_net_7538_bfr_after (
		.din(new_net_7537),
		.dout(new_net_7538)
	);

	bfr new_net_7539_bfr_after (
		.din(new_net_7538),
		.dout(new_net_7539)
	);

	bfr new_net_7540_bfr_after (
		.din(new_net_7539),
		.dout(new_net_7540)
	);

	bfr new_net_7541_bfr_after (
		.din(new_net_7540),
		.dout(new_net_7541)
	);

	bfr new_net_7542_bfr_after (
		.din(new_net_7541),
		.dout(new_net_7542)
	);

	bfr new_net_7543_bfr_after (
		.din(new_net_7542),
		.dout(new_net_7543)
	);

	bfr new_net_7544_bfr_after (
		.din(new_net_7543),
		.dout(new_net_7544)
	);

	bfr new_net_7545_bfr_after (
		.din(new_net_7544),
		.dout(new_net_7545)
	);

	bfr new_net_7546_bfr_after (
		.din(new_net_7545),
		.dout(new_net_7546)
	);

	bfr new_net_7547_bfr_after (
		.din(new_net_7546),
		.dout(new_net_7547)
	);

	bfr new_net_7548_bfr_after (
		.din(new_net_7547),
		.dout(new_net_7548)
	);

	bfr new_net_7549_bfr_after (
		.din(new_net_7548),
		.dout(new_net_7549)
	);

	bfr new_net_7550_bfr_after (
		.din(new_net_7549),
		.dout(new_net_7550)
	);

	bfr new_net_7551_bfr_after (
		.din(new_net_7550),
		.dout(new_net_7551)
	);

	bfr new_net_7552_bfr_after (
		.din(new_net_7551),
		.dout(new_net_7552)
	);

	bfr new_net_7553_bfr_after (
		.din(new_net_7552),
		.dout(new_net_7553)
	);

	bfr new_net_7554_bfr_after (
		.din(new_net_7553),
		.dout(new_net_7554)
	);

	bfr new_net_7555_bfr_after (
		.din(new_net_7554),
		.dout(new_net_7555)
	);

	bfr new_net_7556_bfr_after (
		.din(new_net_7555),
		.dout(new_net_7556)
	);

	bfr new_net_7557_bfr_after (
		.din(new_net_7556),
		.dout(new_net_7557)
	);

	bfr new_net_7558_bfr_after (
		.din(new_net_7557),
		.dout(new_net_7558)
	);

	bfr new_net_7559_bfr_after (
		.din(new_net_7558),
		.dout(new_net_7559)
	);

	bfr new_net_7560_bfr_after (
		.din(new_net_7559),
		.dout(new_net_7560)
	);

	bfr new_net_7561_bfr_after (
		.din(new_net_7560),
		.dout(new_net_7561)
	);

	bfr new_net_7562_bfr_after (
		.din(new_net_7561),
		.dout(new_net_7562)
	);

	bfr new_net_7563_bfr_after (
		.din(new_net_7562),
		.dout(new_net_7563)
	);

	bfr new_net_7564_bfr_after (
		.din(new_net_7563),
		.dout(new_net_7564)
	);

	bfr new_net_7565_bfr_after (
		.din(new_net_7564),
		.dout(new_net_7565)
	);

	bfr new_net_7566_bfr_after (
		.din(new_net_7565),
		.dout(new_net_7566)
	);

	bfr G5235_bfr_after (
		.din(new_net_7566),
		.dout(G5235)
	);

	bfr new_net_7567_bfr_after (
		.din(G112),
		.dout(new_net_7567)
	);

	bfr new_net_2239_bfr_after (
		.din(new_net_7567),
		.dout(new_net_2239)
	);

	bfr new_net_7568_bfr_after (
		.din(_0476_),
		.dout(new_net_7568)
	);

	bfr new_net_7569_bfr_after (
		.din(new_net_7568),
		.dout(new_net_7569)
	);

	bfr new_net_7570_bfr_after (
		.din(new_net_7569),
		.dout(new_net_7570)
	);

	bfr new_net_7571_bfr_after (
		.din(new_net_7570),
		.dout(new_net_7571)
	);

	bfr new_net_7572_bfr_after (
		.din(new_net_7571),
		.dout(new_net_7572)
	);

	bfr new_net_7573_bfr_after (
		.din(new_net_7572),
		.dout(new_net_7573)
	);

	bfr new_net_7574_bfr_after (
		.din(new_net_7573),
		.dout(new_net_7574)
	);

	bfr new_net_7575_bfr_after (
		.din(new_net_7574),
		.dout(new_net_7575)
	);

	bfr new_net_7576_bfr_after (
		.din(new_net_7575),
		.dout(new_net_7576)
	);

	bfr new_net_7577_bfr_after (
		.din(new_net_7576),
		.dout(new_net_7577)
	);

	bfr new_net_7578_bfr_after (
		.din(new_net_7577),
		.dout(new_net_7578)
	);

	bfr new_net_7579_bfr_after (
		.din(new_net_7578),
		.dout(new_net_7579)
	);

	bfr new_net_7580_bfr_after (
		.din(new_net_7579),
		.dout(new_net_7580)
	);

	bfr new_net_7581_bfr_after (
		.din(new_net_7580),
		.dout(new_net_7581)
	);

	bfr new_net_7582_bfr_after (
		.din(new_net_7581),
		.dout(new_net_7582)
	);

	bfr new_net_7583_bfr_after (
		.din(new_net_7582),
		.dout(new_net_7583)
	);

	bfr new_net_7584_bfr_after (
		.din(new_net_7583),
		.dout(new_net_7584)
	);

	bfr new_net_7585_bfr_after (
		.din(new_net_7584),
		.dout(new_net_7585)
	);

	bfr new_net_7586_bfr_after (
		.din(new_net_7585),
		.dout(new_net_7586)
	);

	bfr new_net_7587_bfr_after (
		.din(new_net_7586),
		.dout(new_net_7587)
	);

	bfr new_net_7588_bfr_after (
		.din(new_net_7587),
		.dout(new_net_7588)
	);

	bfr new_net_7589_bfr_after (
		.din(new_net_7588),
		.dout(new_net_7589)
	);

	bfr new_net_7590_bfr_after (
		.din(new_net_7589),
		.dout(new_net_7590)
	);

	bfr new_net_7591_bfr_after (
		.din(new_net_7590),
		.dout(new_net_7591)
	);

	bfr new_net_7592_bfr_after (
		.din(new_net_7591),
		.dout(new_net_7592)
	);

	bfr new_net_7593_bfr_after (
		.din(new_net_7592),
		.dout(new_net_7593)
	);

	bfr new_net_7594_bfr_after (
		.din(new_net_7593),
		.dout(new_net_7594)
	);

	bfr new_net_7595_bfr_after (
		.din(new_net_7594),
		.dout(new_net_7595)
	);

	bfr new_net_2323_bfr_after (
		.din(new_net_7595),
		.dout(new_net_2323)
	);

	bfr new_net_2260_bfr_after (
		.din(_0239_),
		.dout(new_net_2260)
	);

	bfr new_net_7596_bfr_after (
		.din(new_net_2387),
		.dout(new_net_7596)
	);

	bfr new_net_7597_bfr_after (
		.din(new_net_7596),
		.dout(new_net_7597)
	);

	bfr new_net_7598_bfr_after (
		.din(new_net_7597),
		.dout(new_net_7598)
	);

	bfr new_net_7599_bfr_after (
		.din(new_net_7598),
		.dout(new_net_7599)
	);

	bfr new_net_7600_bfr_after (
		.din(new_net_7599),
		.dout(new_net_7600)
	);

	bfr new_net_7601_bfr_after (
		.din(new_net_7600),
		.dout(new_net_7601)
	);

	bfr new_net_7602_bfr_after (
		.din(new_net_7601),
		.dout(new_net_7602)
	);

	bfr new_net_7603_bfr_after (
		.din(new_net_7602),
		.dout(new_net_7603)
	);

	bfr new_net_7604_bfr_after (
		.din(new_net_7603),
		.dout(new_net_7604)
	);

	bfr new_net_7605_bfr_after (
		.din(new_net_7604),
		.dout(new_net_7605)
	);

	bfr G5278_bfr_after (
		.din(new_net_7605),
		.dout(G5278)
	);

	bfr new_net_7606_bfr_after (
		.din(_0677_),
		.dout(new_net_7606)
	);

	bfr new_net_7607_bfr_after (
		.din(new_net_7606),
		.dout(new_net_7607)
	);

	bfr new_net_2134_bfr_after (
		.din(new_net_7607),
		.dout(new_net_2134)
	);

	bfr new_net_7608_bfr_after (
		.din(_1027_),
		.dout(new_net_7608)
	);

	bfr new_net_7609_bfr_after (
		.din(new_net_7608),
		.dout(new_net_7609)
	);

	bfr new_net_7610_bfr_after (
		.din(new_net_7609),
		.dout(new_net_7610)
	);

	bfr new_net_7611_bfr_after (
		.din(new_net_7610),
		.dout(new_net_7611)
	);

	bfr new_net_7612_bfr_after (
		.din(new_net_7611),
		.dout(new_net_7612)
	);

	bfr new_net_7613_bfr_after (
		.din(new_net_7612),
		.dout(new_net_7613)
	);

	bfr new_net_7614_bfr_after (
		.din(new_net_7613),
		.dout(new_net_7614)
	);

	bfr new_net_7615_bfr_after (
		.din(new_net_7614),
		.dout(new_net_7615)
	);

	bfr new_net_7616_bfr_after (
		.din(new_net_7615),
		.dout(new_net_7616)
	);

	bfr new_net_7617_bfr_after (
		.din(new_net_7616),
		.dout(new_net_7617)
	);

	bfr new_net_7618_bfr_after (
		.din(new_net_7617),
		.dout(new_net_7618)
	);

	bfr new_net_7619_bfr_after (
		.din(new_net_7618),
		.dout(new_net_7619)
	);

	bfr new_net_7620_bfr_after (
		.din(new_net_7619),
		.dout(new_net_7620)
	);

	bfr new_net_7621_bfr_after (
		.din(new_net_7620),
		.dout(new_net_7621)
	);

	bfr new_net_7622_bfr_after (
		.din(new_net_7621),
		.dout(new_net_7622)
	);

	bfr new_net_7623_bfr_after (
		.din(new_net_7622),
		.dout(new_net_7623)
	);

	bfr new_net_7624_bfr_after (
		.din(new_net_7623),
		.dout(new_net_7624)
	);

	bfr new_net_7625_bfr_after (
		.din(new_net_7624),
		.dout(new_net_7625)
	);

	bfr new_net_7626_bfr_after (
		.din(new_net_7625),
		.dout(new_net_7626)
	);

	bfr new_net_7627_bfr_after (
		.din(new_net_7626),
		.dout(new_net_7627)
	);

	bfr new_net_2197_bfr_after (
		.din(new_net_7627),
		.dout(new_net_2197)
	);

	bfr new_net_7628_bfr_after (
		.din(_0287_),
		.dout(new_net_7628)
	);

	bfr new_net_7629_bfr_after (
		.din(new_net_7628),
		.dout(new_net_7629)
	);

	bfr new_net_2276_bfr_after (
		.din(new_net_7629),
		.dout(new_net_2276)
	);

	bfr new_net_7630_bfr_after (
		.din(_0556_),
		.dout(new_net_7630)
	);

	bfr new_net_7631_bfr_after (
		.din(new_net_7630),
		.dout(new_net_7631)
	);

	bfr new_net_7632_bfr_after (
		.din(new_net_7631),
		.dout(new_net_7632)
	);

	bfr new_net_7633_bfr_after (
		.din(new_net_7632),
		.dout(new_net_7633)
	);

	bfr new_net_7634_bfr_after (
		.din(new_net_7633),
		.dout(new_net_7634)
	);

	bfr new_net_7635_bfr_after (
		.din(new_net_7634),
		.dout(new_net_7635)
	);

	bfr new_net_7636_bfr_after (
		.din(new_net_7635),
		.dout(new_net_7636)
	);

	bfr new_net_7637_bfr_after (
		.din(new_net_7636),
		.dout(new_net_7637)
	);

	bfr new_net_7638_bfr_after (
		.din(new_net_7637),
		.dout(new_net_7638)
	);

	bfr new_net_7639_bfr_after (
		.din(new_net_7638),
		.dout(new_net_7639)
	);

	bfr new_net_7640_bfr_after (
		.din(new_net_7639),
		.dout(new_net_7640)
	);

	bfr new_net_7641_bfr_after (
		.din(new_net_7640),
		.dout(new_net_7641)
	);

	bfr new_net_7642_bfr_after (
		.din(new_net_7641),
		.dout(new_net_7642)
	);

	bfr new_net_7643_bfr_after (
		.din(new_net_7642),
		.dout(new_net_7643)
	);

	bfr new_net_7644_bfr_after (
		.din(new_net_7643),
		.dout(new_net_7644)
	);

	bfr new_net_7645_bfr_after (
		.din(new_net_7644),
		.dout(new_net_7645)
	);

	bfr new_net_2339_bfr_after (
		.din(new_net_7645),
		.dout(new_net_2339)
	);

	bfr new_net_2129_bfr_after (
		.din(_0636_),
		.dout(new_net_2129)
	);

	bfr new_net_7646_bfr_after (
		.din(G104),
		.dout(new_net_7646)
	);

	bfr new_net_2150_bfr_after (
		.din(new_net_7646),
		.dout(new_net_2150)
	);

	bfr new_net_7647_bfr_after (
		.din(G118),
		.dout(new_net_7647)
	);

	bfr new_net_7648_bfr_after (
		.din(new_net_7647),
		.dout(new_net_7648)
	);

	bfr new_net_2171_bfr_after (
		.din(new_net_7648),
		.dout(new_net_2171)
	);

	bfr new_net_2108_bfr_after (
		.din(_0585_),
		.dout(new_net_2108)
	);

	bfr new_net_7649_bfr_after (
		.din(_0928_),
		.dout(new_net_7649)
	);

	bfr new_net_7650_bfr_after (
		.din(new_net_7649),
		.dout(new_net_7650)
	);

	bfr new_net_7651_bfr_after (
		.din(new_net_7650),
		.dout(new_net_7651)
	);

	bfr new_net_7652_bfr_after (
		.din(new_net_7651),
		.dout(new_net_7652)
	);

	bfr new_net_7653_bfr_after (
		.din(new_net_7652),
		.dout(new_net_7653)
	);

	bfr new_net_7654_bfr_after (
		.din(new_net_7653),
		.dout(new_net_7654)
	);

	bfr new_net_7655_bfr_after (
		.din(new_net_7654),
		.dout(new_net_7655)
	);

	bfr new_net_7656_bfr_after (
		.din(new_net_7655),
		.dout(new_net_7656)
	);

	bfr new_net_7657_bfr_after (
		.din(new_net_7656),
		.dout(new_net_7657)
	);

	bfr new_net_7658_bfr_after (
		.din(new_net_7657),
		.dout(new_net_7658)
	);

	bfr new_net_7659_bfr_after (
		.din(new_net_7658),
		.dout(new_net_7659)
	);

	bfr new_net_7660_bfr_after (
		.din(new_net_7659),
		.dout(new_net_7660)
	);

	bfr new_net_7661_bfr_after (
		.din(new_net_7660),
		.dout(new_net_7661)
	);

	bfr new_net_7662_bfr_after (
		.din(new_net_7661),
		.dout(new_net_7662)
	);

	bfr new_net_7663_bfr_after (
		.din(new_net_7662),
		.dout(new_net_7663)
	);

	bfr new_net_7664_bfr_after (
		.din(new_net_7663),
		.dout(new_net_7664)
	);

	bfr new_net_7665_bfr_after (
		.din(new_net_7664),
		.dout(new_net_7665)
	);

	bfr new_net_7666_bfr_after (
		.din(new_net_7665),
		.dout(new_net_7666)
	);

	bfr new_net_7667_bfr_after (
		.din(new_net_7666),
		.dout(new_net_7667)
	);

	bfr new_net_7668_bfr_after (
		.din(new_net_7667),
		.dout(new_net_7668)
	);

	bfr new_net_7669_bfr_after (
		.din(new_net_7668),
		.dout(new_net_7669)
	);

	bfr new_net_7670_bfr_after (
		.din(new_net_7669),
		.dout(new_net_7670)
	);

	bfr new_net_7671_bfr_after (
		.din(new_net_7670),
		.dout(new_net_7671)
	);

	bfr new_net_7672_bfr_after (
		.din(new_net_7671),
		.dout(new_net_7672)
	);

	bfr new_net_7673_bfr_after (
		.din(new_net_7672),
		.dout(new_net_7673)
	);

	bfr new_net_2192_bfr_after (
		.din(new_net_7673),
		.dout(new_net_2192)
	);

	bfr new_net_7674_bfr_after (
		.din(_0375_),
		.dout(new_net_7674)
	);

	bfr new_net_7675_bfr_after (
		.din(new_net_7674),
		.dout(new_net_7675)
	);

	bfr new_net_2297_bfr_after (
		.din(new_net_7675),
		.dout(new_net_2297)
	);

	bfr new_net_2213_bfr_after (
		.din(_1122_),
		.dout(new_net_2213)
	);

	bfr new_net_7676_bfr_after (
		.din(_0101_),
		.dout(new_net_7676)
	);

	bfr new_net_7677_bfr_after (
		.din(new_net_7676),
		.dout(new_net_7677)
	);

	bfr new_net_2234_bfr_after (
		.din(new_net_7677),
		.dout(new_net_2234)
	);

	bfr new_net_7678_bfr_after (
		.din(new_net_2425),
		.dout(new_net_7678)
	);

	bfr new_net_7679_bfr_after (
		.din(new_net_7678),
		.dout(new_net_7679)
	);

	bfr new_net_7680_bfr_after (
		.din(new_net_7679),
		.dout(new_net_7680)
	);

	bfr new_net_7681_bfr_after (
		.din(new_net_7680),
		.dout(new_net_7681)
	);

	bfr new_net_7682_bfr_after (
		.din(new_net_7681),
		.dout(new_net_7682)
	);

	bfr new_net_7683_bfr_after (
		.din(new_net_7682),
		.dout(new_net_7683)
	);

	bfr new_net_7684_bfr_after (
		.din(new_net_7683),
		.dout(new_net_7684)
	);

	bfr new_net_7685_bfr_after (
		.din(new_net_7684),
		.dout(new_net_7685)
	);

	bfr new_net_7686_bfr_after (
		.din(new_net_7685),
		.dout(new_net_7686)
	);

	bfr new_net_7687_bfr_after (
		.din(new_net_7686),
		.dout(new_net_7687)
	);

	bfr new_net_7688_bfr_after (
		.din(new_net_7687),
		.dout(new_net_7688)
	);

	bfr new_net_7689_bfr_after (
		.din(new_net_7688),
		.dout(new_net_7689)
	);

	bfr new_net_7690_bfr_after (
		.din(new_net_7689),
		.dout(new_net_7690)
	);

	bfr new_net_7691_bfr_after (
		.din(new_net_7690),
		.dout(new_net_7691)
	);

	bfr new_net_7692_bfr_after (
		.din(new_net_7691),
		.dout(new_net_7692)
	);

	bfr new_net_7693_bfr_after (
		.din(new_net_7692),
		.dout(new_net_7693)
	);

	bfr new_net_7694_bfr_after (
		.din(new_net_7693),
		.dout(new_net_7694)
	);

	bfr new_net_7695_bfr_after (
		.din(new_net_7694),
		.dout(new_net_7695)
	);

	bfr new_net_7696_bfr_after (
		.din(new_net_7695),
		.dout(new_net_7696)
	);

	bfr new_net_7697_bfr_after (
		.din(new_net_7696),
		.dout(new_net_7697)
	);

	bfr new_net_7698_bfr_after (
		.din(new_net_7697),
		.dout(new_net_7698)
	);

	bfr new_net_7699_bfr_after (
		.din(new_net_7698),
		.dout(new_net_7699)
	);

	bfr new_net_7700_bfr_after (
		.din(new_net_7699),
		.dout(new_net_7700)
	);

	bfr G5239_bfr_after (
		.din(new_net_7700),
		.dout(G5239)
	);

	bfr new_net_7701_bfr_after (
		.din(new_net_2493),
		.dout(new_net_7701)
	);

	bfr new_net_7702_bfr_after (
		.din(new_net_7701),
		.dout(new_net_7702)
	);

	bfr G5307_bfr_after (
		.din(new_net_7702),
		.dout(G5307)
	);

	bfr new_net_7703_bfr_after (
		.din(new_net_2349),
		.dout(new_net_7703)
	);

	bfr G5313_bfr_after (
		.din(new_net_7703),
		.dout(G5313)
	);

	bfr new_net_7704_bfr_after (
		.din(new_net_2361),
		.dout(new_net_7704)
	);

	bfr new_net_7705_bfr_after (
		.din(new_net_7704),
		.dout(new_net_7705)
	);

	bfr new_net_7706_bfr_after (
		.din(new_net_7705),
		.dout(new_net_7706)
	);

	bfr new_net_7707_bfr_after (
		.din(new_net_7706),
		.dout(new_net_7707)
	);

	bfr G5302_bfr_after (
		.din(new_net_7707),
		.dout(G5302)
	);

	bfr new_net_7708_bfr_after (
		.din(new_net_2373),
		.dout(new_net_7708)
	);

	bfr new_net_7709_bfr_after (
		.din(new_net_7708),
		.dout(new_net_7709)
	);

	bfr new_net_7710_bfr_after (
		.din(new_net_7709),
		.dout(new_net_7710)
	);

	bfr new_net_7711_bfr_after (
		.din(new_net_7710),
		.dout(new_net_7711)
	);

	bfr new_net_7712_bfr_after (
		.din(new_net_7711),
		.dout(new_net_7712)
	);

	bfr new_net_7713_bfr_after (
		.din(new_net_7712),
		.dout(new_net_7713)
	);

	bfr new_net_7714_bfr_after (
		.din(new_net_7713),
		.dout(new_net_7714)
	);

	bfr new_net_7715_bfr_after (
		.din(new_net_7714),
		.dout(new_net_7715)
	);

	bfr new_net_7716_bfr_after (
		.din(new_net_7715),
		.dout(new_net_7716)
	);

	bfr new_net_7717_bfr_after (
		.din(new_net_7716),
		.dout(new_net_7717)
	);

	bfr new_net_7718_bfr_after (
		.din(new_net_7717),
		.dout(new_net_7718)
	);

	bfr new_net_7719_bfr_after (
		.din(new_net_7718),
		.dout(new_net_7719)
	);

	bfr new_net_7720_bfr_after (
		.din(new_net_7719),
		.dout(new_net_7720)
	);

	bfr new_net_7721_bfr_after (
		.din(new_net_7720),
		.dout(new_net_7721)
	);

	bfr new_net_7722_bfr_after (
		.din(new_net_7721),
		.dout(new_net_7722)
	);

	bfr new_net_7723_bfr_after (
		.din(new_net_7722),
		.dout(new_net_7723)
	);

	bfr new_net_7724_bfr_after (
		.din(new_net_7723),
		.dout(new_net_7724)
	);

	bfr new_net_7725_bfr_after (
		.din(new_net_7724),
		.dout(new_net_7725)
	);

	bfr new_net_7726_bfr_after (
		.din(new_net_7725),
		.dout(new_net_7726)
	);

	bfr new_net_7727_bfr_after (
		.din(new_net_7726),
		.dout(new_net_7727)
	);

	bfr new_net_7728_bfr_after (
		.din(new_net_7727),
		.dout(new_net_7728)
	);

	bfr G5244_bfr_after (
		.din(new_net_7728),
		.dout(G5244)
	);

	bfr new_net_7729_bfr_after (
		.din(new_net_2385),
		.dout(new_net_7729)
	);

	bfr new_net_7730_bfr_after (
		.din(new_net_7729),
		.dout(new_net_7730)
	);

	bfr new_net_7731_bfr_after (
		.din(new_net_7730),
		.dout(new_net_7731)
	);

	bfr new_net_7732_bfr_after (
		.din(new_net_7731),
		.dout(new_net_7732)
	);

	bfr new_net_7733_bfr_after (
		.din(new_net_7732),
		.dout(new_net_7733)
	);

	bfr new_net_7734_bfr_after (
		.din(new_net_7733),
		.dout(new_net_7734)
	);

	bfr new_net_7735_bfr_after (
		.din(new_net_7734),
		.dout(new_net_7735)
	);

	bfr new_net_7736_bfr_after (
		.din(new_net_7735),
		.dout(new_net_7736)
	);

	bfr new_net_7737_bfr_after (
		.din(new_net_7736),
		.dout(new_net_7737)
	);

	bfr new_net_7738_bfr_after (
		.din(new_net_7737),
		.dout(new_net_7738)
	);

	bfr new_net_7739_bfr_after (
		.din(new_net_7738),
		.dout(new_net_7739)
	);

	bfr new_net_7740_bfr_after (
		.din(new_net_7739),
		.dout(new_net_7740)
	);

	bfr new_net_7741_bfr_after (
		.din(new_net_7740),
		.dout(new_net_7741)
	);

	bfr new_net_7742_bfr_after (
		.din(new_net_7741),
		.dout(new_net_7742)
	);

	bfr new_net_7743_bfr_after (
		.din(new_net_7742),
		.dout(new_net_7743)
	);

	bfr new_net_7744_bfr_after (
		.din(new_net_7743),
		.dout(new_net_7744)
	);

	bfr new_net_7745_bfr_after (
		.din(new_net_7744),
		.dout(new_net_7745)
	);

	bfr new_net_7746_bfr_after (
		.din(new_net_7745),
		.dout(new_net_7746)
	);

	bfr new_net_7747_bfr_after (
		.din(new_net_7746),
		.dout(new_net_7747)
	);

	bfr new_net_7748_bfr_after (
		.din(new_net_7747),
		.dout(new_net_7748)
	);

	bfr new_net_7749_bfr_after (
		.din(new_net_7748),
		.dout(new_net_7749)
	);

	bfr G5246_bfr_after (
		.din(new_net_7749),
		.dout(G5246)
	);

	bfr new_net_7750_bfr_after (
		.din(new_net_2397),
		.dout(new_net_7750)
	);

	bfr new_net_7751_bfr_after (
		.din(new_net_7750),
		.dout(new_net_7751)
	);

	bfr new_net_7752_bfr_after (
		.din(new_net_7751),
		.dout(new_net_7752)
	);

	bfr new_net_7753_bfr_after (
		.din(new_net_7752),
		.dout(new_net_7753)
	);

	bfr new_net_7754_bfr_after (
		.din(new_net_7753),
		.dout(new_net_7754)
	);

	bfr new_net_7755_bfr_after (
		.din(new_net_7754),
		.dout(new_net_7755)
	);

	bfr new_net_7756_bfr_after (
		.din(new_net_7755),
		.dout(new_net_7756)
	);

	bfr new_net_7757_bfr_after (
		.din(new_net_7756),
		.dout(new_net_7757)
	);

	bfr new_net_7758_bfr_after (
		.din(new_net_7757),
		.dout(new_net_7758)
	);

	bfr new_net_7759_bfr_after (
		.din(new_net_7758),
		.dout(new_net_7759)
	);

	bfr new_net_7760_bfr_after (
		.din(new_net_7759),
		.dout(new_net_7760)
	);

	bfr new_net_7761_bfr_after (
		.din(new_net_7760),
		.dout(new_net_7761)
	);

	bfr new_net_7762_bfr_after (
		.din(new_net_7761),
		.dout(new_net_7762)
	);

	bfr new_net_7763_bfr_after (
		.din(new_net_7762),
		.dout(new_net_7763)
	);

	bfr new_net_7764_bfr_after (
		.din(new_net_7763),
		.dout(new_net_7764)
	);

	bfr new_net_7765_bfr_after (
		.din(new_net_7764),
		.dout(new_net_7765)
	);

	bfr new_net_7766_bfr_after (
		.din(new_net_7765),
		.dout(new_net_7766)
	);

	bfr new_net_7767_bfr_after (
		.din(new_net_7766),
		.dout(new_net_7767)
	);

	bfr G5266_bfr_after (
		.din(new_net_7767),
		.dout(G5266)
	);

	bfr new_net_7768_bfr_after (
		.din(new_net_2409),
		.dout(new_net_7768)
	);

	bfr new_net_7769_bfr_after (
		.din(new_net_7768),
		.dout(new_net_7769)
	);

	bfr new_net_7770_bfr_after (
		.din(new_net_7769),
		.dout(new_net_7770)
	);

	bfr new_net_7771_bfr_after (
		.din(new_net_7770),
		.dout(new_net_7771)
	);

	bfr new_net_7772_bfr_after (
		.din(new_net_7771),
		.dout(new_net_7772)
	);

	bfr G5311_bfr_after (
		.din(new_net_7772),
		.dout(G5311)
	);

	bfr new_net_7773_bfr_after (
		.din(_0279_),
		.dout(new_net_7773)
	);

	bfr new_net_2271_bfr_after (
		.din(new_net_7773),
		.dout(new_net_2271)
	);

	bfr new_net_7774_bfr_after (
		.din(_0528_),
		.dout(new_net_7774)
	);

	bfr new_net_7775_bfr_after (
		.din(new_net_7774),
		.dout(new_net_7775)
	);

	bfr new_net_7776_bfr_after (
		.din(new_net_7775),
		.dout(new_net_7776)
	);

	bfr new_net_7777_bfr_after (
		.din(new_net_7776),
		.dout(new_net_7777)
	);

	bfr new_net_7778_bfr_after (
		.din(new_net_7777),
		.dout(new_net_7778)
	);

	bfr new_net_7779_bfr_after (
		.din(new_net_7778),
		.dout(new_net_7779)
	);

	bfr new_net_7780_bfr_after (
		.din(new_net_7779),
		.dout(new_net_7780)
	);

	bfr new_net_7781_bfr_after (
		.din(new_net_7780),
		.dout(new_net_7781)
	);

	bfr new_net_7782_bfr_after (
		.din(new_net_7781),
		.dout(new_net_7782)
	);

	bfr new_net_7783_bfr_after (
		.din(new_net_7782),
		.dout(new_net_7783)
	);

	bfr new_net_7784_bfr_after (
		.din(new_net_7783),
		.dout(new_net_7784)
	);

	bfr new_net_7785_bfr_after (
		.din(new_net_7784),
		.dout(new_net_7785)
	);

	bfr new_net_7786_bfr_after (
		.din(new_net_7785),
		.dout(new_net_7786)
	);

	bfr new_net_7787_bfr_after (
		.din(new_net_7786),
		.dout(new_net_7787)
	);

	bfr new_net_7788_bfr_after (
		.din(new_net_7787),
		.dout(new_net_7788)
	);

	bfr new_net_7789_bfr_after (
		.din(new_net_7788),
		.dout(new_net_7789)
	);

	bfr new_net_7790_bfr_after (
		.din(new_net_7789),
		.dout(new_net_7790)
	);

	bfr new_net_7791_bfr_after (
		.din(new_net_7790),
		.dout(new_net_7791)
	);

	bfr new_net_7792_bfr_after (
		.din(new_net_7791),
		.dout(new_net_7792)
	);

	bfr new_net_7793_bfr_after (
		.din(new_net_7792),
		.dout(new_net_7793)
	);

	bfr new_net_7794_bfr_after (
		.din(new_net_7793),
		.dout(new_net_7794)
	);

	bfr new_net_7795_bfr_after (
		.din(new_net_7794),
		.dout(new_net_7795)
	);

	bfr new_net_7796_bfr_after (
		.din(new_net_7795),
		.dout(new_net_7796)
	);

	bfr new_net_7797_bfr_after (
		.din(new_net_7796),
		.dout(new_net_7797)
	);

	bfr new_net_7798_bfr_after (
		.din(new_net_7797),
		.dout(new_net_7798)
	);

	bfr new_net_7799_bfr_after (
		.din(new_net_7798),
		.dout(new_net_7799)
	);

	bfr new_net_7800_bfr_after (
		.din(new_net_7799),
		.dout(new_net_7800)
	);

	bfr new_net_7801_bfr_after (
		.din(new_net_7800),
		.dout(new_net_7801)
	);

	bfr new_net_7802_bfr_after (
		.din(new_net_7801),
		.dout(new_net_7802)
	);

	bfr new_net_7803_bfr_after (
		.din(new_net_7802),
		.dout(new_net_7803)
	);

	bfr new_net_2334_bfr_after (
		.din(new_net_7803),
		.dout(new_net_2334)
	);

	bfr new_net_7804_bfr_after (
		.din(new_net_2391),
		.dout(new_net_7804)
	);

	bfr new_net_7805_bfr_after (
		.din(new_net_7804),
		.dout(new_net_7805)
	);

	bfr G5309_bfr_after (
		.din(new_net_7805),
		.dout(G5309)
	);

	bfr new_net_7806_bfr_after (
		.din(_0617_),
		.dout(new_net_7806)
	);

	bfr new_net_2124_bfr_after (
		.din(new_net_7806),
		.dout(new_net_2124)
	);

	bfr new_net_7807_bfr_after (
		.din(G97),
		.dout(new_net_7807)
	);

	bfr new_net_2145_bfr_after (
		.din(new_net_7807),
		.dout(new_net_2145)
	);

	bfr new_net_2187_bfr_after (
		.din(_0945_),
		.dout(new_net_2187)
	);

	bfr new_net_7808_bfr_after (
		.din(_0352_),
		.dout(new_net_7808)
	);

	bfr new_net_2292_bfr_after (
		.din(new_net_7808),
		.dout(new_net_2292)
	);

	bfr new_net_7809_bfr_after (
		.din(new_net_2379),
		.dout(new_net_7809)
	);

	bfr new_net_7810_bfr_after (
		.din(new_net_7809),
		.dout(new_net_7810)
	);

	bfr new_net_7811_bfr_after (
		.din(new_net_7810),
		.dout(new_net_7811)
	);

	bfr new_net_7812_bfr_after (
		.din(new_net_7811),
		.dout(new_net_7812)
	);

	bfr new_net_7813_bfr_after (
		.din(new_net_7812),
		.dout(new_net_7813)
	);

	bfr new_net_7814_bfr_after (
		.din(new_net_7813),
		.dout(new_net_7814)
	);

	bfr new_net_7815_bfr_after (
		.din(new_net_7814),
		.dout(new_net_7815)
	);

	bfr new_net_7816_bfr_after (
		.din(new_net_7815),
		.dout(new_net_7816)
	);

	bfr new_net_7817_bfr_after (
		.din(new_net_7816),
		.dout(new_net_7817)
	);

	bfr new_net_7818_bfr_after (
		.din(new_net_7817),
		.dout(new_net_7818)
	);

	bfr new_net_7819_bfr_after (
		.din(new_net_7818),
		.dout(new_net_7819)
	);

	bfr new_net_7820_bfr_after (
		.din(new_net_7819),
		.dout(new_net_7820)
	);

	bfr new_net_7821_bfr_after (
		.din(new_net_7820),
		.dout(new_net_7821)
	);

	bfr new_net_7822_bfr_after (
		.din(new_net_7821),
		.dout(new_net_7822)
	);

	bfr new_net_7823_bfr_after (
		.din(new_net_7822),
		.dout(new_net_7823)
	);

	bfr new_net_7824_bfr_after (
		.din(new_net_7823),
		.dout(new_net_7824)
	);

	bfr new_net_7825_bfr_after (
		.din(new_net_7824),
		.dout(new_net_7825)
	);

	bfr new_net_7826_bfr_after (
		.din(new_net_7825),
		.dout(new_net_7826)
	);

	bfr new_net_7827_bfr_after (
		.din(new_net_7826),
		.dout(new_net_7827)
	);

	bfr new_net_7828_bfr_after (
		.din(new_net_7827),
		.dout(new_net_7828)
	);

	bfr new_net_7829_bfr_after (
		.din(new_net_7828),
		.dout(new_net_7829)
	);

	bfr new_net_7830_bfr_after (
		.din(new_net_7829),
		.dout(new_net_7830)
	);

	bfr new_net_7831_bfr_after (
		.din(new_net_7830),
		.dout(new_net_7831)
	);

	bfr new_net_7832_bfr_after (
		.din(new_net_7831),
		.dout(new_net_7832)
	);

	bfr new_net_7833_bfr_after (
		.din(new_net_7832),
		.dout(new_net_7833)
	);

	bfr new_net_7834_bfr_after (
		.din(new_net_7833),
		.dout(new_net_7834)
	);

	bfr new_net_7835_bfr_after (
		.din(new_net_7834),
		.dout(new_net_7835)
	);

	bfr new_net_7836_bfr_after (
		.din(new_net_7835),
		.dout(new_net_7836)
	);

	bfr new_net_7837_bfr_after (
		.din(new_net_7836),
		.dout(new_net_7837)
	);

	bfr new_net_7838_bfr_after (
		.din(new_net_7837),
		.dout(new_net_7838)
	);

	bfr new_net_7839_bfr_after (
		.din(new_net_7838),
		.dout(new_net_7839)
	);

	bfr new_net_7840_bfr_after (
		.din(new_net_7839),
		.dout(new_net_7840)
	);

	bfr new_net_7841_bfr_after (
		.din(new_net_7840),
		.dout(new_net_7841)
	);

	bfr new_net_7842_bfr_after (
		.din(new_net_7841),
		.dout(new_net_7842)
	);

	bfr new_net_7843_bfr_after (
		.din(new_net_7842),
		.dout(new_net_7843)
	);

	bfr new_net_7844_bfr_after (
		.din(new_net_7843),
		.dout(new_net_7844)
	);

	bfr new_net_7845_bfr_after (
		.din(new_net_7844),
		.dout(new_net_7845)
	);

	bfr new_net_7846_bfr_after (
		.din(new_net_7845),
		.dout(new_net_7846)
	);

	bfr new_net_7847_bfr_after (
		.din(new_net_7846),
		.dout(new_net_7847)
	);

	bfr G5193_bfr_after (
		.din(new_net_7847),
		.dout(G5193)
	);

	bfr new_net_7848_bfr_after (
		.din(_0848_),
		.dout(new_net_7848)
	);

	bfr new_net_7849_bfr_after (
		.din(new_net_7848),
		.dout(new_net_7849)
	);

	bfr new_net_7850_bfr_after (
		.din(new_net_7849),
		.dout(new_net_7850)
	);

	bfr new_net_7851_bfr_after (
		.din(new_net_7850),
		.dout(new_net_7851)
	);

	bfr new_net_7852_bfr_after (
		.din(new_net_7851),
		.dout(new_net_7852)
	);

	bfr new_net_7853_bfr_after (
		.din(new_net_7852),
		.dout(new_net_7853)
	);

	bfr new_net_7854_bfr_after (
		.din(new_net_7853),
		.dout(new_net_7854)
	);

	bfr new_net_7855_bfr_after (
		.din(new_net_7854),
		.dout(new_net_7855)
	);

	bfr new_net_2166_bfr_after (
		.din(new_net_7855),
		.dout(new_net_2166)
	);

	bfr new_net_2208_bfr_after (
		.din(_1097_),
		.dout(new_net_2208)
	);

	bfr new_net_7856_bfr_after (
		.din(_0791_),
		.dout(new_net_7856)
	);

	bfr new_net_7857_bfr_after (
		.din(new_net_7856),
		.dout(new_net_7857)
	);

	bfr new_net_7858_bfr_after (
		.din(new_net_7857),
		.dout(new_net_7858)
	);

	bfr new_net_7859_bfr_after (
		.din(new_net_7858),
		.dout(new_net_7859)
	);

	bfr new_net_7860_bfr_after (
		.din(new_net_7859),
		.dout(new_net_7860)
	);

	bfr new_net_7861_bfr_after (
		.din(new_net_7860),
		.dout(new_net_7861)
	);

	bfr new_net_7862_bfr_after (
		.din(new_net_7861),
		.dout(new_net_7862)
	);

	bfr new_net_7863_bfr_after (
		.din(new_net_7862),
		.dout(new_net_7863)
	);

	bfr new_net_7864_bfr_after (
		.din(new_net_7863),
		.dout(new_net_7864)
	);

	bfr new_net_7865_bfr_after (
		.din(new_net_7864),
		.dout(new_net_7865)
	);

	bfr new_net_7866_bfr_after (
		.din(new_net_7865),
		.dout(new_net_7866)
	);

	bfr new_net_7867_bfr_after (
		.din(new_net_7866),
		.dout(new_net_7867)
	);

	bfr new_net_7868_bfr_after (
		.din(new_net_7867),
		.dout(new_net_7868)
	);

	bfr new_net_7869_bfr_after (
		.din(new_net_7868),
		.dout(new_net_7869)
	);

	bfr new_net_7870_bfr_after (
		.din(new_net_7869),
		.dout(new_net_7870)
	);

	bfr new_net_7871_bfr_after (
		.din(new_net_7870),
		.dout(new_net_7871)
	);

	bfr new_net_7872_bfr_after (
		.din(new_net_7871),
		.dout(new_net_7872)
	);

	bfr new_net_2159_bfr_after (
		.din(new_net_7872),
		.dout(new_net_2159)
	);

	bfr new_net_7873_bfr_after (
		.din(G60),
		.dout(new_net_7873)
	);

	bfr new_net_7874_bfr_after (
		.din(new_net_7873),
		.dout(new_net_7874)
	);

	bfr new_net_7875_bfr_after (
		.din(new_net_7874),
		.dout(new_net_7875)
	);

	bfr new_net_7876_bfr_after (
		.din(new_net_7875),
		.dout(new_net_7876)
	);

	bfr new_net_2119_bfr_after (
		.din(new_net_7876),
		.dout(new_net_2119)
	);

	bfr new_net_7877_bfr_after (
		.din(_0216_),
		.dout(new_net_7877)
	);

	bfr new_net_2245_bfr_after (
		.din(new_net_7877),
		.dout(new_net_2245)
	);

	bfr new_net_7878_bfr_after (
		.din(_0506_),
		.dout(new_net_7878)
	);

	bfr new_net_2329_bfr_after (
		.din(new_net_7878),
		.dout(new_net_2329)
	);

	bfr new_net_7879_bfr_after (
		.din(_0270_),
		.dout(new_net_7879)
	);

	bfr new_net_7880_bfr_after (
		.din(new_net_7879),
		.dout(new_net_7880)
	);

	bfr new_net_7881_bfr_after (
		.din(new_net_7880),
		.dout(new_net_7881)
	);

	bfr new_net_7882_bfr_after (
		.din(new_net_7881),
		.dout(new_net_7882)
	);

	bfr new_net_7883_bfr_after (
		.din(new_net_7882),
		.dout(new_net_7883)
	);

	bfr new_net_7884_bfr_after (
		.din(new_net_7883),
		.dout(new_net_7884)
	);

	bfr new_net_7885_bfr_after (
		.din(new_net_7884),
		.dout(new_net_7885)
	);

	bfr new_net_7886_bfr_after (
		.din(new_net_7885),
		.dout(new_net_7886)
	);

	bfr new_net_7887_bfr_after (
		.din(new_net_7886),
		.dout(new_net_7887)
	);

	bfr new_net_7888_bfr_after (
		.din(new_net_7887),
		.dout(new_net_7888)
	);

	bfr new_net_7889_bfr_after (
		.din(new_net_7888),
		.dout(new_net_7889)
	);

	bfr new_net_7890_bfr_after (
		.din(new_net_7889),
		.dout(new_net_7890)
	);

	bfr new_net_7891_bfr_after (
		.din(new_net_7890),
		.dout(new_net_7891)
	);

	bfr new_net_7892_bfr_after (
		.din(new_net_7891),
		.dout(new_net_7892)
	);

	bfr new_net_2266_bfr_after (
		.din(new_net_7892),
		.dout(new_net_2266)
	);

	bfr new_net_7893_bfr_after (
		.din(_0702_),
		.dout(new_net_7893)
	);

	bfr new_net_7894_bfr_after (
		.din(new_net_7893),
		.dout(new_net_7894)
	);

	bfr new_net_7895_bfr_after (
		.din(new_net_7894),
		.dout(new_net_7895)
	);

	bfr new_net_7896_bfr_after (
		.din(new_net_7895),
		.dout(new_net_7896)
	);

	bfr new_net_7897_bfr_after (
		.din(new_net_7896),
		.dout(new_net_7897)
	);

	bfr new_net_7898_bfr_after (
		.din(new_net_7897),
		.dout(new_net_7898)
	);

	bfr new_net_7899_bfr_after (
		.din(new_net_7898),
		.dout(new_net_7899)
	);

	bfr new_net_7900_bfr_after (
		.din(new_net_7899),
		.dout(new_net_7900)
	);

	bfr new_net_7901_bfr_after (
		.din(new_net_7900),
		.dout(new_net_7901)
	);

	bfr new_net_7902_bfr_after (
		.din(new_net_7901),
		.dout(new_net_7902)
	);

	bfr new_net_7903_bfr_after (
		.din(new_net_7902),
		.dout(new_net_7903)
	);

	bfr new_net_7904_bfr_after (
		.din(new_net_7903),
		.dout(new_net_7904)
	);

	bfr new_net_7905_bfr_after (
		.din(new_net_7904),
		.dout(new_net_7905)
	);

	bfr new_net_7906_bfr_after (
		.din(new_net_7905),
		.dout(new_net_7906)
	);

	bfr new_net_7907_bfr_after (
		.din(new_net_7906),
		.dout(new_net_7907)
	);

	bfr new_net_2140_bfr_after (
		.din(new_net_7907),
		.dout(new_net_2140)
	);

	bfr new_net_2161_bfr_after (
		.din(_0826_),
		.dout(new_net_2161)
	);

	bfr new_net_7908_bfr_after (
		.din(G46),
		.dout(new_net_7908)
	);

	bfr new_net_7909_bfr_after (
		.din(new_net_7908),
		.dout(new_net_7909)
	);

	bfr new_net_7910_bfr_after (
		.din(new_net_7909),
		.dout(new_net_7910)
	);

	bfr new_net_7911_bfr_after (
		.din(new_net_7910),
		.dout(new_net_7911)
	);

	bfr new_net_2182_bfr_after (
		.din(new_net_7911),
		.dout(new_net_2182)
	);

	bfr new_net_7912_bfr_after (
		.din(_1052_),
		.dout(new_net_7912)
	);

	bfr new_net_7913_bfr_after (
		.din(new_net_7912),
		.dout(new_net_7913)
	);

	bfr new_net_7914_bfr_after (
		.din(new_net_7913),
		.dout(new_net_7914)
	);

	bfr new_net_2203_bfr_after (
		.din(new_net_7914),
		.dout(new_net_2203)
	);

	bfr new_net_7915_bfr_after (
		.din(_0335_),
		.dout(new_net_7915)
	);

	bfr new_net_7916_bfr_after (
		.din(new_net_7915),
		.dout(new_net_7916)
	);

	bfr new_net_7917_bfr_after (
		.din(new_net_7916),
		.dout(new_net_7917)
	);

	bfr new_net_7918_bfr_after (
		.din(new_net_7917),
		.dout(new_net_7918)
	);

	bfr new_net_7919_bfr_after (
		.din(new_net_7918),
		.dout(new_net_7919)
	);

	bfr new_net_7920_bfr_after (
		.din(new_net_7919),
		.dout(new_net_7920)
	);

	bfr new_net_7921_bfr_after (
		.din(new_net_7920),
		.dout(new_net_7921)
	);

	bfr new_net_7922_bfr_after (
		.din(new_net_7921),
		.dout(new_net_7922)
	);

	bfr new_net_7923_bfr_after (
		.din(new_net_7922),
		.dout(new_net_7923)
	);

	bfr new_net_7924_bfr_after (
		.din(new_net_7923),
		.dout(new_net_7924)
	);

	bfr new_net_7925_bfr_after (
		.din(new_net_7924),
		.dout(new_net_7925)
	);

	bfr new_net_7926_bfr_after (
		.din(new_net_7925),
		.dout(new_net_7926)
	);

	bfr new_net_7927_bfr_after (
		.din(new_net_7926),
		.dout(new_net_7927)
	);

	bfr new_net_7928_bfr_after (
		.din(new_net_7927),
		.dout(new_net_7928)
	);

	bfr new_net_7929_bfr_after (
		.din(new_net_7928),
		.dout(new_net_7929)
	);

	bfr new_net_7930_bfr_after (
		.din(new_net_7929),
		.dout(new_net_7930)
	);

	bfr new_net_7931_bfr_after (
		.din(new_net_7930),
		.dout(new_net_7931)
	);

	bfr new_net_7932_bfr_after (
		.din(new_net_7931),
		.dout(new_net_7932)
	);

	bfr new_net_7933_bfr_after (
		.din(new_net_7932),
		.dout(new_net_7933)
	);

	bfr new_net_7934_bfr_after (
		.din(new_net_7933),
		.dout(new_net_7934)
	);

	bfr new_net_7935_bfr_after (
		.din(new_net_7934),
		.dout(new_net_7935)
	);

	bfr new_net_7936_bfr_after (
		.din(new_net_7935),
		.dout(new_net_7936)
	);

	bfr new_net_7937_bfr_after (
		.din(new_net_7936),
		.dout(new_net_7937)
	);

	bfr new_net_2287_bfr_after (
		.din(new_net_7937),
		.dout(new_net_2287)
	);

	bfr new_net_7938_bfr_after (
		.din(_0009_),
		.dout(new_net_7938)
	);

	bfr new_net_2224_bfr_after (
		.din(new_net_7938),
		.dout(new_net_2224)
	);

	bfr new_net_7939_bfr_after (
		.din(new_net_2461),
		.dout(new_net_7939)
	);

	bfr new_net_7940_bfr_after (
		.din(new_net_7939),
		.dout(new_net_7940)
	);

	bfr new_net_7941_bfr_after (
		.din(new_net_7940),
		.dout(new_net_7941)
	);

	bfr new_net_7942_bfr_after (
		.din(new_net_7941),
		.dout(new_net_7942)
	);

	bfr new_net_7943_bfr_after (
		.din(new_net_7942),
		.dout(new_net_7943)
	);

	bfr new_net_7944_bfr_after (
		.din(new_net_7943),
		.dout(new_net_7944)
	);

	bfr new_net_7945_bfr_after (
		.din(new_net_7944),
		.dout(new_net_7945)
	);

	bfr new_net_7946_bfr_after (
		.din(new_net_7945),
		.dout(new_net_7946)
	);

	bfr new_net_7947_bfr_after (
		.din(new_net_7946),
		.dout(new_net_7947)
	);

	bfr G5275_bfr_after (
		.din(new_net_7947),
		.dout(G5275)
	);

	bfr new_net_7948_bfr_after (
		.din(_1230_),
		.dout(new_net_7948)
	);

	bfr new_net_7949_bfr_after (
		.din(new_net_7948),
		.dout(new_net_7949)
	);

	bfr new_net_2219_bfr_after (
		.din(new_net_7949),
		.dout(new_net_2219)
	);

	bfr new_net_7950_bfr_after (
		.din(_0403_),
		.dout(new_net_7950)
	);

	bfr new_net_7951_bfr_after (
		.din(new_net_7950),
		.dout(new_net_7951)
	);

	bfr new_net_7952_bfr_after (
		.din(new_net_7951),
		.dout(new_net_7952)
	);

	bfr new_net_7953_bfr_after (
		.din(new_net_7952),
		.dout(new_net_7953)
	);

	bfr new_net_7954_bfr_after (
		.din(new_net_7953),
		.dout(new_net_7954)
	);

	bfr new_net_7955_bfr_after (
		.din(new_net_7954),
		.dout(new_net_7955)
	);

	bfr new_net_7956_bfr_after (
		.din(new_net_7955),
		.dout(new_net_7956)
	);

	bfr new_net_7957_bfr_after (
		.din(new_net_7956),
		.dout(new_net_7957)
	);

	bfr new_net_7958_bfr_after (
		.din(new_net_7957),
		.dout(new_net_7958)
	);

	bfr new_net_7959_bfr_after (
		.din(new_net_7958),
		.dout(new_net_7959)
	);

	bfr new_net_7960_bfr_after (
		.din(new_net_7959),
		.dout(new_net_7960)
	);

	bfr new_net_7961_bfr_after (
		.din(new_net_7960),
		.dout(new_net_7961)
	);

	bfr new_net_7962_bfr_after (
		.din(new_net_7961),
		.dout(new_net_7962)
	);

	bfr new_net_7963_bfr_after (
		.din(new_net_7962),
		.dout(new_net_7963)
	);

	bfr new_net_7964_bfr_after (
		.din(new_net_7963),
		.dout(new_net_7964)
	);

	bfr new_net_7965_bfr_after (
		.din(new_net_7964),
		.dout(new_net_7965)
	);

	bfr new_net_7966_bfr_after (
		.din(new_net_7965),
		.dout(new_net_7966)
	);

	bfr new_net_7967_bfr_after (
		.din(new_net_7966),
		.dout(new_net_7967)
	);

	bfr new_net_2303_bfr_after (
		.din(new_net_7967),
		.dout(new_net_2303)
	);

	bfr new_net_2240_bfr_after (
		.din(G67),
		.dout(new_net_2240)
	);

	bfr new_net_7968_bfr_after (
		.din(_0483_),
		.dout(new_net_7968)
	);

	bfr new_net_7969_bfr_after (
		.din(new_net_7968),
		.dout(new_net_7969)
	);

	bfr new_net_7970_bfr_after (
		.din(new_net_7969),
		.dout(new_net_7970)
	);

	bfr new_net_7971_bfr_after (
		.din(new_net_7970),
		.dout(new_net_7971)
	);

	bfr new_net_7972_bfr_after (
		.din(new_net_7971),
		.dout(new_net_7972)
	);

	bfr new_net_7973_bfr_after (
		.din(new_net_7972),
		.dout(new_net_7973)
	);

	bfr new_net_7974_bfr_after (
		.din(new_net_7973),
		.dout(new_net_7974)
	);

	bfr new_net_7975_bfr_after (
		.din(new_net_7974),
		.dout(new_net_7975)
	);

	bfr new_net_7976_bfr_after (
		.din(new_net_7975),
		.dout(new_net_7976)
	);

	bfr new_net_7977_bfr_after (
		.din(new_net_7976),
		.dout(new_net_7977)
	);

	bfr new_net_7978_bfr_after (
		.din(new_net_7977),
		.dout(new_net_7978)
	);

	bfr new_net_7979_bfr_after (
		.din(new_net_7978),
		.dout(new_net_7979)
	);

	bfr new_net_7980_bfr_after (
		.din(new_net_7979),
		.dout(new_net_7980)
	);

	bfr new_net_7981_bfr_after (
		.din(new_net_7980),
		.dout(new_net_7981)
	);

	bfr new_net_7982_bfr_after (
		.din(new_net_7981),
		.dout(new_net_7982)
	);

	bfr new_net_7983_bfr_after (
		.din(new_net_7982),
		.dout(new_net_7983)
	);

	bfr new_net_7984_bfr_after (
		.din(new_net_7983),
		.dout(new_net_7984)
	);

	bfr new_net_7985_bfr_after (
		.din(new_net_7984),
		.dout(new_net_7985)
	);

	bfr new_net_7986_bfr_after (
		.din(new_net_7985),
		.dout(new_net_7986)
	);

	bfr new_net_7987_bfr_after (
		.din(new_net_7986),
		.dout(new_net_7987)
	);

	bfr new_net_7988_bfr_after (
		.din(new_net_7987),
		.dout(new_net_7988)
	);

	bfr new_net_7989_bfr_after (
		.din(new_net_7988),
		.dout(new_net_7989)
	);

	bfr new_net_7990_bfr_after (
		.din(new_net_7989),
		.dout(new_net_7990)
	);

	bfr new_net_7991_bfr_after (
		.din(new_net_7990),
		.dout(new_net_7991)
	);

	bfr new_net_7992_bfr_after (
		.din(new_net_7991),
		.dout(new_net_7992)
	);

	bfr new_net_7993_bfr_after (
		.din(new_net_7992),
		.dout(new_net_7993)
	);

	bfr new_net_7994_bfr_after (
		.din(new_net_7993),
		.dout(new_net_7994)
	);

	bfr new_net_7995_bfr_after (
		.din(new_net_7994),
		.dout(new_net_7995)
	);

	bfr new_net_7996_bfr_after (
		.din(new_net_7995),
		.dout(new_net_7996)
	);

	bfr new_net_7997_bfr_after (
		.din(new_net_7996),
		.dout(new_net_7997)
	);

	bfr new_net_2324_bfr_after (
		.din(new_net_7997),
		.dout(new_net_2324)
	);

	bfr new_net_2261_bfr_after (
		.din(_0238_),
		.dout(new_net_2261)
	);

	bfr new_net_7998_bfr_after (
		.din(_0566_),
		.dout(new_net_7998)
	);

	bfr new_net_7999_bfr_after (
		.din(new_net_7998),
		.dout(new_net_7999)
	);

	bfr new_net_2345_bfr_after (
		.din(new_net_7999),
		.dout(new_net_2345)
	);

	bfr new_net_8000_bfr_after (
		.din(G122),
		.dout(new_net_8000)
	);

	bfr new_net_8001_bfr_after (
		.din(new_net_8000),
		.dout(new_net_8001)
	);

	bfr new_net_2135_bfr_after (
		.din(new_net_8001),
		.dout(new_net_2135)
	);

	bfr new_net_8002_bfr_after (
		.din(G57),
		.dout(new_net_8002)
	);

	bfr new_net_8003_bfr_after (
		.din(new_net_8002),
		.dout(new_net_8003)
	);

	bfr new_net_8004_bfr_after (
		.din(new_net_8003),
		.dout(new_net_8004)
	);

	bfr new_net_8005_bfr_after (
		.din(new_net_8004),
		.dout(new_net_8005)
	);

	bfr new_net_2156_bfr_after (
		.din(new_net_8005),
		.dout(new_net_2156)
	);

	bfr new_net_8006_bfr_after (
		.din(_0908_),
		.dout(new_net_8006)
	);

	bfr new_net_8007_bfr_after (
		.din(new_net_8006),
		.dout(new_net_8007)
	);

	bfr new_net_8008_bfr_after (
		.din(new_net_8007),
		.dout(new_net_8008)
	);

	bfr new_net_8009_bfr_after (
		.din(new_net_8008),
		.dout(new_net_8009)
	);

	bfr new_net_8010_bfr_after (
		.din(new_net_8009),
		.dout(new_net_8010)
	);

	bfr new_net_8011_bfr_after (
		.din(new_net_8010),
		.dout(new_net_8011)
	);

	bfr new_net_8012_bfr_after (
		.din(new_net_8011),
		.dout(new_net_8012)
	);

	bfr new_net_8013_bfr_after (
		.din(new_net_8012),
		.dout(new_net_8013)
	);

	bfr new_net_8014_bfr_after (
		.din(new_net_8013),
		.dout(new_net_8014)
	);

	bfr new_net_8015_bfr_after (
		.din(new_net_8014),
		.dout(new_net_8015)
	);

	bfr new_net_8016_bfr_after (
		.din(new_net_8015),
		.dout(new_net_8016)
	);

	bfr new_net_8017_bfr_after (
		.din(new_net_8016),
		.dout(new_net_8017)
	);

	bfr new_net_8018_bfr_after (
		.din(new_net_8017),
		.dout(new_net_8018)
	);

	bfr new_net_8019_bfr_after (
		.din(new_net_8018),
		.dout(new_net_8019)
	);

	bfr new_net_8020_bfr_after (
		.din(new_net_8019),
		.dout(new_net_8020)
	);

	bfr new_net_8021_bfr_after (
		.din(new_net_8020),
		.dout(new_net_8021)
	);

	bfr new_net_8022_bfr_after (
		.din(new_net_8021),
		.dout(new_net_8022)
	);

	bfr new_net_8023_bfr_after (
		.din(new_net_8022),
		.dout(new_net_8023)
	);

	bfr new_net_8024_bfr_after (
		.din(new_net_8023),
		.dout(new_net_8024)
	);

	bfr new_net_8025_bfr_after (
		.din(new_net_8024),
		.dout(new_net_8025)
	);

	bfr new_net_2177_bfr_after (
		.din(new_net_8025),
		.dout(new_net_2177)
	);

	bfr new_net_2114_bfr_after (
		.din(_0588_),
		.dout(new_net_2114)
	);

	bfr new_net_8026_bfr_after (
		.din(_0961_),
		.dout(new_net_8026)
	);

	bfr new_net_8027_bfr_after (
		.din(new_net_8026),
		.dout(new_net_8027)
	);

	bfr new_net_8028_bfr_after (
		.din(new_net_8027),
		.dout(new_net_8028)
	);

	bfr new_net_8029_bfr_after (
		.din(new_net_8028),
		.dout(new_net_8029)
	);

	bfr new_net_2190_bfr_after (
		.din(new_net_8029),
		.dout(new_net_2190)
	);

	bfr new_net_8030_bfr_after (
		.din(new_net_2505),
		.dout(new_net_8030)
	);

	bfr new_net_8031_bfr_after (
		.din(new_net_8030),
		.dout(new_net_8031)
	);

	bfr new_net_8032_bfr_after (
		.din(new_net_8031),
		.dout(new_net_8032)
	);

	bfr new_net_8033_bfr_after (
		.din(new_net_8032),
		.dout(new_net_8033)
	);

	bfr new_net_8034_bfr_after (
		.din(new_net_8033),
		.dout(new_net_8034)
	);

	bfr new_net_8035_bfr_after (
		.din(new_net_8034),
		.dout(new_net_8035)
	);

	bfr new_net_8036_bfr_after (
		.din(new_net_8035),
		.dout(new_net_8036)
	);

	bfr new_net_8037_bfr_after (
		.din(new_net_8036),
		.dout(new_net_8037)
	);

	bfr new_net_8038_bfr_after (
		.din(new_net_8037),
		.dout(new_net_8038)
	);

	bfr new_net_8039_bfr_after (
		.din(new_net_8038),
		.dout(new_net_8039)
	);

	bfr new_net_8040_bfr_after (
		.din(new_net_8039),
		.dout(new_net_8040)
	);

	bfr new_net_8041_bfr_after (
		.din(new_net_8040),
		.dout(new_net_8041)
	);

	bfr new_net_8042_bfr_after (
		.din(new_net_8041),
		.dout(new_net_8042)
	);

	bfr new_net_8043_bfr_after (
		.din(new_net_8042),
		.dout(new_net_8043)
	);

	bfr new_net_8044_bfr_after (
		.din(new_net_8043),
		.dout(new_net_8044)
	);

	bfr new_net_8045_bfr_after (
		.din(new_net_8044),
		.dout(new_net_8045)
	);

	bfr new_net_8046_bfr_after (
		.din(new_net_8045),
		.dout(new_net_8046)
	);

	bfr new_net_8047_bfr_after (
		.din(new_net_8046),
		.dout(new_net_8047)
	);

	bfr new_net_8048_bfr_after (
		.din(new_net_8047),
		.dout(new_net_8048)
	);

	bfr new_net_8049_bfr_after (
		.din(new_net_8048),
		.dout(new_net_8049)
	);

	bfr new_net_8050_bfr_after (
		.din(new_net_8049),
		.dout(new_net_8050)
	);

	bfr G5261_bfr_after (
		.din(new_net_8050),
		.dout(G5261)
	);

	bfr new_net_8051_bfr_after (
		.din(_0314_),
		.dout(new_net_8051)
	);

	bfr new_net_8052_bfr_after (
		.din(new_net_8051),
		.dout(new_net_8052)
	);

	bfr new_net_8053_bfr_after (
		.din(new_net_8052),
		.dout(new_net_8053)
	);

	bfr new_net_8054_bfr_after (
		.din(new_net_8053),
		.dout(new_net_8054)
	);

	bfr new_net_8055_bfr_after (
		.din(new_net_8054),
		.dout(new_net_8055)
	);

	bfr new_net_8056_bfr_after (
		.din(new_net_8055),
		.dout(new_net_8056)
	);

	bfr new_net_8057_bfr_after (
		.din(new_net_8056),
		.dout(new_net_8057)
	);

	bfr new_net_8058_bfr_after (
		.din(new_net_8057),
		.dout(new_net_8058)
	);

	bfr new_net_8059_bfr_after (
		.din(new_net_8058),
		.dout(new_net_8059)
	);

	bfr new_net_8060_bfr_after (
		.din(new_net_8059),
		.dout(new_net_8060)
	);

	bfr new_net_8061_bfr_after (
		.din(new_net_8060),
		.dout(new_net_8061)
	);

	bfr new_net_8062_bfr_after (
		.din(new_net_8061),
		.dout(new_net_8062)
	);

	bfr new_net_8063_bfr_after (
		.din(new_net_8062),
		.dout(new_net_8063)
	);

	bfr new_net_8064_bfr_after (
		.din(new_net_8063),
		.dout(new_net_8064)
	);

	bfr new_net_8065_bfr_after (
		.din(new_net_8064),
		.dout(new_net_8065)
	);

	bfr new_net_8066_bfr_after (
		.din(new_net_8065),
		.dout(new_net_8066)
	);

	bfr new_net_8067_bfr_after (
		.din(new_net_8066),
		.dout(new_net_8067)
	);

	bfr new_net_8068_bfr_after (
		.din(new_net_8067),
		.dout(new_net_8068)
	);

	bfr new_net_8069_bfr_after (
		.din(new_net_8068),
		.dout(new_net_8069)
	);

	bfr new_net_8070_bfr_after (
		.din(new_net_8069),
		.dout(new_net_8070)
	);

	bfr new_net_8071_bfr_after (
		.din(new_net_8070),
		.dout(new_net_8071)
	);

	bfr new_net_8072_bfr_after (
		.din(new_net_8071),
		.dout(new_net_8072)
	);

	bfr new_net_2282_bfr_after (
		.din(new_net_8072),
		.dout(new_net_2282)
	);

	bfr new_net_8073_bfr_after (
		.din(G45),
		.dout(new_net_8073)
	);

	bfr new_net_8074_bfr_after (
		.din(new_net_8073),
		.dout(new_net_8074)
	);

	bfr new_net_8075_bfr_after (
		.din(new_net_8074),
		.dout(new_net_8075)
	);

	bfr new_net_8076_bfr_after (
		.din(new_net_8075),
		.dout(new_net_8076)
	);

	bfr new_net_2193_bfr_after (
		.din(new_net_8076),
		.dout(new_net_2193)
	);

	bfr new_net_8077_bfr_after (
		.din(_0379_),
		.dout(new_net_8077)
	);

	bfr new_net_8078_bfr_after (
		.din(new_net_8077),
		.dout(new_net_8078)
	);

	bfr new_net_8079_bfr_after (
		.din(new_net_8078),
		.dout(new_net_8079)
	);

	bfr new_net_8080_bfr_after (
		.din(new_net_8079),
		.dout(new_net_8080)
	);

	bfr new_net_8081_bfr_after (
		.din(new_net_8080),
		.dout(new_net_8081)
	);

	bfr new_net_8082_bfr_after (
		.din(new_net_8081),
		.dout(new_net_8082)
	);

	bfr new_net_8083_bfr_after (
		.din(new_net_8082),
		.dout(new_net_8083)
	);

	bfr new_net_8084_bfr_after (
		.din(new_net_8083),
		.dout(new_net_8084)
	);

	bfr new_net_8085_bfr_after (
		.din(new_net_8084),
		.dout(new_net_8085)
	);

	bfr new_net_8086_bfr_after (
		.din(new_net_8085),
		.dout(new_net_8086)
	);

	bfr new_net_8087_bfr_after (
		.din(new_net_8086),
		.dout(new_net_8087)
	);

	bfr new_net_8088_bfr_after (
		.din(new_net_8087),
		.dout(new_net_8088)
	);

	bfr new_net_8089_bfr_after (
		.din(new_net_8088),
		.dout(new_net_8089)
	);

	bfr new_net_8090_bfr_after (
		.din(new_net_8089),
		.dout(new_net_8090)
	);

	bfr new_net_8091_bfr_after (
		.din(new_net_8090),
		.dout(new_net_8091)
	);

	bfr new_net_8092_bfr_after (
		.din(new_net_8091),
		.dout(new_net_8092)
	);

	bfr new_net_8093_bfr_after (
		.din(new_net_8092),
		.dout(new_net_8093)
	);

	bfr new_net_8094_bfr_after (
		.din(new_net_8093),
		.dout(new_net_8094)
	);

	bfr new_net_8095_bfr_after (
		.din(new_net_8094),
		.dout(new_net_8095)
	);

	bfr new_net_8096_bfr_after (
		.din(new_net_8095),
		.dout(new_net_8096)
	);

	bfr new_net_8097_bfr_after (
		.din(new_net_8096),
		.dout(new_net_8097)
	);

	bfr new_net_8098_bfr_after (
		.din(new_net_8097),
		.dout(new_net_8098)
	);

	bfr new_net_2298_bfr_after (
		.din(new_net_8098),
		.dout(new_net_2298)
	);

	bfr new_net_2214_bfr_after (
		.din(_1219_),
		.dout(new_net_2214)
	);

	bfr new_net_8099_bfr_after (
		.din(_0462_),
		.dout(new_net_8099)
	);

	bfr new_net_8100_bfr_after (
		.din(new_net_8099),
		.dout(new_net_8100)
	);

	bfr new_net_8101_bfr_after (
		.din(new_net_8100),
		.dout(new_net_8101)
	);

	bfr new_net_8102_bfr_after (
		.din(new_net_8101),
		.dout(new_net_8102)
	);

	bfr new_net_8103_bfr_after (
		.din(new_net_8102),
		.dout(new_net_8103)
	);

	bfr new_net_8104_bfr_after (
		.din(new_net_8103),
		.dout(new_net_8104)
	);

	bfr new_net_8105_bfr_after (
		.din(new_net_8104),
		.dout(new_net_8105)
	);

	bfr new_net_8106_bfr_after (
		.din(new_net_8105),
		.dout(new_net_8106)
	);

	bfr new_net_8107_bfr_after (
		.din(new_net_8106),
		.dout(new_net_8107)
	);

	bfr new_net_8108_bfr_after (
		.din(new_net_8107),
		.dout(new_net_8108)
	);

	bfr new_net_8109_bfr_after (
		.din(new_net_8108),
		.dout(new_net_8109)
	);

	bfr new_net_8110_bfr_after (
		.din(new_net_8109),
		.dout(new_net_8110)
	);

	bfr new_net_8111_bfr_after (
		.din(new_net_8110),
		.dout(new_net_8111)
	);

	bfr new_net_8112_bfr_after (
		.din(new_net_8111),
		.dout(new_net_8112)
	);

	bfr new_net_8113_bfr_after (
		.din(new_net_8112),
		.dout(new_net_8113)
	);

	bfr new_net_8114_bfr_after (
		.din(new_net_8113),
		.dout(new_net_8114)
	);

	bfr new_net_8115_bfr_after (
		.din(new_net_8114),
		.dout(new_net_8115)
	);

	bfr new_net_8116_bfr_after (
		.din(new_net_8115),
		.dout(new_net_8116)
	);

	bfr new_net_8117_bfr_after (
		.din(new_net_8116),
		.dout(new_net_8117)
	);

	bfr new_net_8118_bfr_after (
		.din(new_net_8117),
		.dout(new_net_8118)
	);

	bfr new_net_8119_bfr_after (
		.din(new_net_8118),
		.dout(new_net_8119)
	);

	bfr new_net_8120_bfr_after (
		.din(new_net_8119),
		.dout(new_net_8120)
	);

	bfr new_net_8121_bfr_after (
		.din(new_net_8120),
		.dout(new_net_8121)
	);

	bfr new_net_8122_bfr_after (
		.din(new_net_8121),
		.dout(new_net_8122)
	);

	bfr new_net_8123_bfr_after (
		.din(new_net_8122),
		.dout(new_net_8123)
	);

	bfr new_net_8124_bfr_after (
		.din(new_net_8123),
		.dout(new_net_8124)
	);

	bfr new_net_8125_bfr_after (
		.din(new_net_8124),
		.dout(new_net_8125)
	);

	bfr new_net_8126_bfr_after (
		.din(new_net_8125),
		.dout(new_net_8126)
	);

	bfr new_net_8127_bfr_after (
		.din(new_net_8126),
		.dout(new_net_8127)
	);

	bfr new_net_8128_bfr_after (
		.din(new_net_8127),
		.dout(new_net_8128)
	);

	bfr new_net_8129_bfr_after (
		.din(new_net_8128),
		.dout(new_net_8129)
	);

	bfr new_net_2319_bfr_after (
		.din(new_net_8129),
		.dout(new_net_2319)
	);

	bfr new_net_8130_bfr_after (
		.din(_0107_),
		.dout(new_net_8130)
	);

	bfr new_net_8131_bfr_after (
		.din(new_net_8130),
		.dout(new_net_8131)
	);

	bfr new_net_8132_bfr_after (
		.din(new_net_8131),
		.dout(new_net_8132)
	);

	bfr new_net_8133_bfr_after (
		.din(new_net_8132),
		.dout(new_net_8133)
	);

	bfr new_net_8134_bfr_after (
		.din(new_net_8133),
		.dout(new_net_8134)
	);

	bfr new_net_8135_bfr_after (
		.din(new_net_8134),
		.dout(new_net_8135)
	);

	bfr new_net_8136_bfr_after (
		.din(new_net_8135),
		.dout(new_net_8136)
	);

	bfr new_net_8137_bfr_after (
		.din(new_net_8136),
		.dout(new_net_8137)
	);

	bfr new_net_8138_bfr_after (
		.din(new_net_8137),
		.dout(new_net_8138)
	);

	bfr new_net_8139_bfr_after (
		.din(new_net_8138),
		.dout(new_net_8139)
	);

	bfr new_net_8140_bfr_after (
		.din(new_net_8139),
		.dout(new_net_8140)
	);

	bfr new_net_8141_bfr_after (
		.din(new_net_8140),
		.dout(new_net_8141)
	);

	bfr new_net_8142_bfr_after (
		.din(new_net_8141),
		.dout(new_net_8142)
	);

	bfr new_net_8143_bfr_after (
		.din(new_net_8142),
		.dout(new_net_8143)
	);

	bfr new_net_8144_bfr_after (
		.din(new_net_8143),
		.dout(new_net_8144)
	);

	bfr new_net_8145_bfr_after (
		.din(new_net_8144),
		.dout(new_net_8145)
	);

	bfr new_net_8146_bfr_after (
		.din(new_net_8145),
		.dout(new_net_8146)
	);

	bfr new_net_8147_bfr_after (
		.din(new_net_8146),
		.dout(new_net_8147)
	);

	bfr new_net_8148_bfr_after (
		.din(new_net_8147),
		.dout(new_net_8148)
	);

	bfr new_net_8149_bfr_after (
		.din(new_net_8148),
		.dout(new_net_8149)
	);

	bfr new_net_8150_bfr_after (
		.din(new_net_8149),
		.dout(new_net_8150)
	);

	bfr new_net_8151_bfr_after (
		.din(new_net_8150),
		.dout(new_net_8151)
	);

	bfr new_net_8152_bfr_after (
		.din(new_net_8151),
		.dout(new_net_8152)
	);

	bfr new_net_8153_bfr_after (
		.din(new_net_8152),
		.dout(new_net_8153)
	);

	bfr new_net_8154_bfr_after (
		.din(new_net_8153),
		.dout(new_net_8154)
	);

	bfr new_net_8155_bfr_after (
		.din(new_net_8154),
		.dout(new_net_8155)
	);

	bfr new_net_8156_bfr_after (
		.din(new_net_8155),
		.dout(new_net_8156)
	);

	bfr new_net_8157_bfr_after (
		.din(new_net_8156),
		.dout(new_net_8157)
	);

	bfr new_net_8158_bfr_after (
		.din(new_net_8157),
		.dout(new_net_8158)
	);

	bfr new_net_8159_bfr_after (
		.din(new_net_8158),
		.dout(new_net_8159)
	);

	bfr new_net_8160_bfr_after (
		.din(new_net_8159),
		.dout(new_net_8160)
	);

	bfr new_net_8161_bfr_after (
		.din(new_net_8160),
		.dout(new_net_8161)
	);

	bfr new_net_2235_bfr_after (
		.din(new_net_8161),
		.dout(new_net_2235)
	);

	bfr new_net_2256_bfr_after (
		.din(_0229_),
		.dout(new_net_2256)
	);

	bfr new_net_8162_bfr_after (
		.din(_0291_),
		.dout(new_net_8162)
	);

	bfr new_net_8163_bfr_after (
		.din(new_net_8162),
		.dout(new_net_8163)
	);

	bfr new_net_8164_bfr_after (
		.din(new_net_8163),
		.dout(new_net_8164)
	);

	bfr new_net_8165_bfr_after (
		.din(new_net_8164),
		.dout(new_net_8165)
	);

	bfr new_net_8166_bfr_after (
		.din(new_net_8165),
		.dout(new_net_8166)
	);

	bfr new_net_8167_bfr_after (
		.din(new_net_8166),
		.dout(new_net_8167)
	);

	bfr new_net_8168_bfr_after (
		.din(new_net_8167),
		.dout(new_net_8168)
	);

	bfr new_net_8169_bfr_after (
		.din(new_net_8168),
		.dout(new_net_8169)
	);

	bfr new_net_8170_bfr_after (
		.din(new_net_8169),
		.dout(new_net_8170)
	);

	bfr new_net_8171_bfr_after (
		.din(new_net_8170),
		.dout(new_net_8171)
	);

	bfr new_net_8172_bfr_after (
		.din(new_net_8171),
		.dout(new_net_8172)
	);

	bfr new_net_8173_bfr_after (
		.din(new_net_8172),
		.dout(new_net_8173)
	);

	bfr new_net_8174_bfr_after (
		.din(new_net_8173),
		.dout(new_net_8174)
	);

	bfr new_net_8175_bfr_after (
		.din(new_net_8174),
		.dout(new_net_8175)
	);

	bfr new_net_2277_bfr_after (
		.din(new_net_8175),
		.dout(new_net_2277)
	);

	bfr new_net_8176_bfr_after (
		.din(_0560_),
		.dout(new_net_8176)
	);

	bfr new_net_8177_bfr_after (
		.din(new_net_8176),
		.dout(new_net_8177)
	);

	bfr new_net_8178_bfr_after (
		.din(new_net_8177),
		.dout(new_net_8178)
	);

	bfr new_net_8179_bfr_after (
		.din(new_net_8178),
		.dout(new_net_8179)
	);

	bfr new_net_8180_bfr_after (
		.din(new_net_8179),
		.dout(new_net_8180)
	);

	bfr new_net_8181_bfr_after (
		.din(new_net_8180),
		.dout(new_net_8181)
	);

	bfr new_net_8182_bfr_after (
		.din(new_net_8181),
		.dout(new_net_8182)
	);

	bfr new_net_8183_bfr_after (
		.din(new_net_8182),
		.dout(new_net_8183)
	);

	bfr new_net_8184_bfr_after (
		.din(new_net_8183),
		.dout(new_net_8184)
	);

	bfr new_net_8185_bfr_after (
		.din(new_net_8184),
		.dout(new_net_8185)
	);

	bfr new_net_8186_bfr_after (
		.din(new_net_8185),
		.dout(new_net_8186)
	);

	bfr new_net_8187_bfr_after (
		.din(new_net_8186),
		.dout(new_net_8187)
	);

	bfr new_net_8188_bfr_after (
		.din(new_net_8187),
		.dout(new_net_8188)
	);

	bfr new_net_8189_bfr_after (
		.din(new_net_8188),
		.dout(new_net_8189)
	);

	bfr new_net_8190_bfr_after (
		.din(new_net_8189),
		.dout(new_net_8190)
	);

	bfr new_net_8191_bfr_after (
		.din(new_net_8190),
		.dout(new_net_8191)
	);

	bfr new_net_8192_bfr_after (
		.din(new_net_8191),
		.dout(new_net_8192)
	);

	bfr new_net_8193_bfr_after (
		.din(new_net_8192),
		.dout(new_net_8193)
	);

	bfr new_net_8194_bfr_after (
		.din(new_net_8193),
		.dout(new_net_8194)
	);

	bfr new_net_8195_bfr_after (
		.din(new_net_8194),
		.dout(new_net_8195)
	);

	bfr new_net_8196_bfr_after (
		.din(new_net_8195),
		.dout(new_net_8196)
	);

	bfr new_net_8197_bfr_after (
		.din(new_net_8196),
		.dout(new_net_8197)
	);

	bfr new_net_8198_bfr_after (
		.din(new_net_8197),
		.dout(new_net_8198)
	);

	bfr new_net_8199_bfr_after (
		.din(new_net_8198),
		.dout(new_net_8199)
	);

	bfr new_net_8200_bfr_after (
		.din(new_net_8199),
		.dout(new_net_8200)
	);

	bfr new_net_8201_bfr_after (
		.din(new_net_8200),
		.dout(new_net_8201)
	);

	bfr new_net_8202_bfr_after (
		.din(new_net_8201),
		.dout(new_net_8202)
	);

	bfr new_net_8203_bfr_after (
		.din(new_net_8202),
		.dout(new_net_8203)
	);

	bfr new_net_8204_bfr_after (
		.din(new_net_8203),
		.dout(new_net_8204)
	);

	bfr new_net_8205_bfr_after (
		.din(new_net_8204),
		.dout(new_net_8205)
	);

	bfr new_net_2340_bfr_after (
		.din(new_net_8205),
		.dout(new_net_2340)
	);

	bfr new_net_2130_bfr_after (
		.din(_0642_),
		.dout(new_net_2130)
	);

	bfr new_net_2151_bfr_after (
		.din(_0756_),
		.dout(new_net_2151)
	);

	bfr new_net_8206_bfr_after (
		.din(_1241_),
		.dout(new_net_8206)
	);

	bfr new_net_8207_bfr_after (
		.din(new_net_8206),
		.dout(new_net_8207)
	);

	bfr new_net_8208_bfr_after (
		.din(new_net_8207),
		.dout(new_net_8208)
	);

	bfr new_net_8209_bfr_after (
		.din(new_net_8208),
		.dout(new_net_8209)
	);

	bfr new_net_8210_bfr_after (
		.din(new_net_8209),
		.dout(new_net_8210)
	);

	bfr new_net_2220_bfr_after (
		.din(new_net_8210),
		.dout(new_net_2220)
	);

	bfr new_net_2225_bfr_after (
		.din(_0025_),
		.dout(new_net_2225)
	);

	bfr new_net_8211_bfr_after (
		.din(new_net_2359),
		.dout(new_net_8211)
	);

	bfr new_net_8212_bfr_after (
		.din(new_net_8211),
		.dout(new_net_8212)
	);

	bfr new_net_8213_bfr_after (
		.din(new_net_8212),
		.dout(new_net_8213)
	);

	bfr new_net_8214_bfr_after (
		.din(new_net_8213),
		.dout(new_net_8214)
	);

	bfr new_net_8215_bfr_after (
		.din(new_net_8214),
		.dout(new_net_8215)
	);

	bfr new_net_8216_bfr_after (
		.din(new_net_8215),
		.dout(new_net_8216)
	);

	bfr new_net_8217_bfr_after (
		.din(new_net_8216),
		.dout(new_net_8217)
	);

	bfr new_net_8218_bfr_after (
		.din(new_net_8217),
		.dout(new_net_8218)
	);

	bfr new_net_8219_bfr_after (
		.din(new_net_8218),
		.dout(new_net_8219)
	);

	bfr new_net_8220_bfr_after (
		.din(new_net_8219),
		.dout(new_net_8220)
	);

	bfr new_net_8221_bfr_after (
		.din(new_net_8220),
		.dout(new_net_8221)
	);

	bfr new_net_8222_bfr_after (
		.din(new_net_8221),
		.dout(new_net_8222)
	);

	bfr new_net_8223_bfr_after (
		.din(new_net_8222),
		.dout(new_net_8223)
	);

	bfr new_net_8224_bfr_after (
		.din(new_net_8223),
		.dout(new_net_8224)
	);

	bfr new_net_8225_bfr_after (
		.din(new_net_8224),
		.dout(new_net_8225)
	);

	bfr new_net_8226_bfr_after (
		.din(new_net_8225),
		.dout(new_net_8226)
	);

	bfr new_net_8227_bfr_after (
		.din(new_net_8226),
		.dout(new_net_8227)
	);

	bfr new_net_8228_bfr_after (
		.din(new_net_8227),
		.dout(new_net_8228)
	);

	bfr new_net_8229_bfr_after (
		.din(new_net_8228),
		.dout(new_net_8229)
	);

	bfr new_net_8230_bfr_after (
		.din(new_net_8229),
		.dout(new_net_8230)
	);

	bfr new_net_8231_bfr_after (
		.din(new_net_8230),
		.dout(new_net_8231)
	);

	bfr new_net_8232_bfr_after (
		.din(new_net_8231),
		.dout(new_net_8232)
	);

	bfr new_net_8233_bfr_after (
		.din(new_net_8232),
		.dout(new_net_8233)
	);

	bfr new_net_8234_bfr_after (
		.din(new_net_8233),
		.dout(new_net_8234)
	);

	bfr new_net_8235_bfr_after (
		.din(new_net_8234),
		.dout(new_net_8235)
	);

	bfr new_net_8236_bfr_after (
		.din(new_net_8235),
		.dout(new_net_8236)
	);

	bfr new_net_8237_bfr_after (
		.din(new_net_8236),
		.dout(new_net_8237)
	);

	bfr new_net_8238_bfr_after (
		.din(new_net_8237),
		.dout(new_net_8238)
	);

	bfr new_net_8239_bfr_after (
		.din(new_net_8238),
		.dout(new_net_8239)
	);

	bfr new_net_8240_bfr_after (
		.din(new_net_8239),
		.dout(new_net_8240)
	);

	bfr new_net_8241_bfr_after (
		.din(new_net_8240),
		.dout(new_net_8241)
	);

	bfr new_net_8242_bfr_after (
		.din(new_net_8241),
		.dout(new_net_8242)
	);

	bfr new_net_8243_bfr_after (
		.din(new_net_8242),
		.dout(new_net_8243)
	);

	bfr new_net_8244_bfr_after (
		.din(new_net_8243),
		.dout(new_net_8244)
	);

	bfr new_net_8245_bfr_after (
		.din(new_net_8244),
		.dout(new_net_8245)
	);

	bfr new_net_8246_bfr_after (
		.din(new_net_8245),
		.dout(new_net_8246)
	);

	bfr new_net_8247_bfr_after (
		.din(new_net_8246),
		.dout(new_net_8247)
	);

	bfr new_net_8248_bfr_after (
		.din(new_net_8247),
		.dout(new_net_8248)
	);

	bfr new_net_8249_bfr_after (
		.din(new_net_8248),
		.dout(new_net_8249)
	);

	bfr G5197_bfr_after (
		.din(new_net_8249),
		.dout(G5197)
	);

	bfr new_net_8250_bfr_after (
		.din(G7),
		.dout(new_net_8250)
	);

	bfr new_net_2250_bfr_after (
		.din(new_net_8250),
		.dout(new_net_2250)
	);

	bfr new_net_8251_bfr_after (
		.din(_0440_),
		.dout(new_net_8251)
	);

	bfr new_net_8252_bfr_after (
		.din(new_net_8251),
		.dout(new_net_8252)
	);

	bfr new_net_2313_bfr_after (
		.din(new_net_8252),
		.dout(new_net_2313)
	);

	bfr new_net_8253_bfr_after (
		.din(_0425_),
		.dout(new_net_8253)
	);

	bfr new_net_8254_bfr_after (
		.din(new_net_8253),
		.dout(new_net_8254)
	);

	bfr new_net_2308_bfr_after (
		.din(new_net_8254),
		.dout(new_net_2308)
	);

	bfr new_net_8255_bfr_after (
		.din(new_net_2411),
		.dout(new_net_8255)
	);

	bfr new_net_8256_bfr_after (
		.din(new_net_8255),
		.dout(new_net_8256)
	);

	bfr new_net_8257_bfr_after (
		.din(new_net_8256),
		.dout(new_net_8257)
	);

	bfr new_net_8258_bfr_after (
		.din(new_net_8257),
		.dout(new_net_8258)
	);

	bfr new_net_8259_bfr_after (
		.din(new_net_8258),
		.dout(new_net_8259)
	);

	bfr new_net_8260_bfr_after (
		.din(new_net_8259),
		.dout(new_net_8260)
	);

	bfr new_net_8261_bfr_after (
		.din(new_net_8260),
		.dout(new_net_8261)
	);

	bfr new_net_8262_bfr_after (
		.din(new_net_8261),
		.dout(new_net_8262)
	);

	bfr new_net_8263_bfr_after (
		.din(new_net_8262),
		.dout(new_net_8263)
	);

	bfr new_net_8264_bfr_after (
		.din(new_net_8263),
		.dout(new_net_8264)
	);

	bfr new_net_8265_bfr_after (
		.din(new_net_8264),
		.dout(new_net_8265)
	);

	bfr new_net_8266_bfr_after (
		.din(new_net_8265),
		.dout(new_net_8266)
	);

	bfr new_net_8267_bfr_after (
		.din(new_net_8266),
		.dout(new_net_8267)
	);

	bfr new_net_8268_bfr_after (
		.din(new_net_8267),
		.dout(new_net_8268)
	);

	bfr new_net_8269_bfr_after (
		.din(new_net_8268),
		.dout(new_net_8269)
	);

	bfr new_net_8270_bfr_after (
		.din(new_net_8269),
		.dout(new_net_8270)
	);

	bfr new_net_8271_bfr_after (
		.din(new_net_8270),
		.dout(new_net_8271)
	);

	bfr new_net_8272_bfr_after (
		.din(new_net_8271),
		.dout(new_net_8272)
	);

	bfr new_net_8273_bfr_after (
		.din(new_net_8272),
		.dout(new_net_8273)
	);

	bfr new_net_8274_bfr_after (
		.din(new_net_8273),
		.dout(new_net_8274)
	);

	bfr new_net_8275_bfr_after (
		.din(new_net_8274),
		.dout(new_net_8275)
	);

	bfr new_net_8276_bfr_after (
		.din(new_net_8275),
		.dout(new_net_8276)
	);

	bfr new_net_8277_bfr_after (
		.din(new_net_8276),
		.dout(new_net_8277)
	);

	bfr new_net_8278_bfr_after (
		.din(new_net_8277),
		.dout(new_net_8278)
	);

	bfr new_net_8279_bfr_after (
		.din(new_net_8278),
		.dout(new_net_8279)
	);

	bfr G5243_bfr_after (
		.din(new_net_8279),
		.dout(G5243)
	);

	bfr new_net_8280_bfr_after (
		.din(_0958_),
		.dout(new_net_8280)
	);

	bfr new_net_8281_bfr_after (
		.din(new_net_8280),
		.dout(new_net_8281)
	);

	bfr new_net_2189_bfr_after (
		.din(new_net_8281),
		.dout(new_net_2189)
	);

endmodule