module c499(N1, N5, N9, N13, N17, N21, N25, N29, N33, N37, N41, N45, N49, N53, N57, N61, N65, N69, N73, N77, N81, N85, N89, N93, N97, N101, N105, N109, N113, N117, N121, N125, N129, N130, N131, N132, N133, N134, N135, N136, N137, N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755);
	wire new_net_1603;
	wire new_net_1732;
	wire _148_;
	wire _274_;
	wire new_net_562;
	wire new_net_514;
	wire new_net_848;
	wire new_net_226;
	wire new_net_295;
	wire new_net_638;
	wire new_net_935;
	wire new_net_1109;
	wire new_net_987;
	wire new_net_1288;
	wire new_net_5;
	wire new_net_23;
	wire new_net_89;
	wire new_net_329;
	wire new_net_347;
	wire new_net_663;
	wire new_net_1022;
	wire new_net_1034;
	wire new_net_1258;
	wire new_net_1337;
	wire new_net_483;
	wire new_net_546;
	wire _149_;
	wire _275_;
	wire new_net_399;
	wire new_net_838;
	wire new_net_531;
	wire new_net_999;
	wire new_net_1054;
	wire new_net_1066;
	wire new_net_1275;
	wire new_net_1408;
	wire new_net_40;
	wire new_net_106;
	wire new_net_124;
	wire new_net_244;
	wire new_net_466;
	wire new_net_956;
	wire new_net_1097;
	wire new_net_1359;
	wire new_net_1371;
	wire new_net_1658;
	wire new_net_1541;
	wire new_net_278;
	wire _150_;
	wire _276_;
	wire new_net_227;
	wire new_net_365;
	wire new_net_563;
	wire new_net_705;
	wire new_net_633;
	wire new_net_1076;
	wire new_net_1122;
	wire new_net_1430;
	wire new_net_1708;
	wire new_net_1352;
	wire new_net_1606;
	wire new_net_1400;
	wire new_net_24;
	wire new_net_312;
	wire new_net_330;
	wire new_net_348;
	wire new_net_787;
	wire new_net_759;
	wire new_net_866;
	wire new_net_768;
	wire new_net_1304;
	wire new_net_1316;
	wire new_net_1464;
	wire new_net_1457;
	wire new_net_818;
	wire _277_;
	wire _151_;
	wire new_net_400;
	wire new_net_484;
	wire new_net_547;
	wire new_net_433;
	wire new_net_902;
	wire new_net_914;
	wire new_net_1584;
	wire new_net_1217;
	wire new_net_107;
	wire new_net_245;
	wire new_net_296;
	wire new_net_467;
	wire new_net_515;
	wire new_net_604;
	wire new_net_849;
	wire new_net_936;
	wire new_net_1058;
	wire new_net_1098;
	wire new_net_1315;
	wire _278_;
	wire _152_;
	wire new_net_6;
	wire new_net_90;
	wire new_net_279;
	wire new_net_856;
	wire new_net_648;
	wire new_net_661;
	wire new_net_366;
	wire new_net_1023;
	wire new_net_1121;
	wire new_net_1331;
	wire new_net_1506;
	wire new_net_313;
	wire new_net_331;
	wire new_net_532;
	wire new_net_588;
	wire new_net_630;
	wire new_net_670;
	wire new_net_839;
	wire _332_;
	wire new_net_1000;
	wire new_net_1055;
	wire new_net_1266;
	wire new_net_1435;
	wire new_net_434;
	wire _279_;
	wire _153_;
	wire new_net_41;
	wire new_net_125;
	wire new_net_548;
	wire new_net_890;
	wire new_net_957;
	wire new_net_1360;
	wire new_net_1372;
	wire new_net_1532;
	wire new_net_1568;
	wire new_net_228;
	wire new_net_297;
	wire new_net_468;
	wire new_net_516;
	wire new_net_564;
	wire new_net_729;
	wire new_net_1077;
	wire new_net_1214;
	wire new_net_1252;
	wire new_net_1383;
	wire new_net_1469;
	wire new_net_1673;
	wire new_net_1386;
	wire new_net_1727;
	wire new_net_1559;
	wire new_net_1638;
	wire new_net_349;
	wire new_net_788;
	wire _280_;
	wire _154_;
	wire new_net_7;
	wire new_net_25;
	wire new_net_760;
	wire new_net_769;
	wire new_net_873;
	wire new_net_606;
	wire new_net_1317;
	wire new_net_1525;
	wire new_net_1693;
	wire new_net_1279;
	wire new_net_401;
	wire new_net_485;
	wire new_net_533;
	wire new_net_819;
	wire new_net_891;
	wire new_net_903;
	wire new_net_1585;
	wire new_net_1597;
	wire new_net_1659;
	wire new_net_1657;
	wire new_net_1203;
	wire new_net_1420;
	wire new_net_1338;
	wire new_net_22;
	wire new_net_1336;
	wire new_net_1084;
	wire _281_;
	wire _155_;
	wire new_net_42;
	wire new_net_549;
	wire new_net_108;
	wire new_net_246;
	wire new_net_126;
	wire new_net_850;
	wire new_net_937;
	wire new_net_1099;
	wire new_net_1511;
	wire new_net_1442;
	wire new_net_1230;
	wire new_net_1713;
	wire new_net_229;
	wire new_net_280;
	wire new_net_298;
	wire new_net_367;
	wire new_net_565;
	wire new_net_577;
	wire new_net_1024;
	wire new_net_1036;
	wire new_net_1260;
	wire new_net_1327;
	wire new_net_1364;
	wire new_net_1404;
	wire new_net_1580;
	wire new_net_1573;
	wire new_net_1537;
	wire new_net_314;
	wire new_net_332;
	wire new_net_637;
	wire _282_;
	wire _156_;
	wire new_net_8;
	wire new_net_26;
	wire new_net_92;
	wire new_net_350;
	wire new_net_840;
	wire new_net_1257;
	wire new_net_1174;
	wire new_net_1428;
	wire new_net_402;
	wire new_net_435;
	wire new_net_486;
	wire new_net_867;
	wire new_net_958;
	wire new_net_1361;
	wire new_net_1373;
	wire new_net_1391;
	wire new_net_1484;
	wire new_net_1660;
	wire new_net_1681;
	wire new_net_1643;
	wire new_net_1070;
	wire new_net_247;
	wire new_net_623;
	wire new_net_517;
	wire _283_;
	wire _157_;
	wire new_net_109;
	wire new_net_730;
	wire new_net_469;
	wire new_net_658;
	wire new_net_707;
	wire new_net_1664;
	wire new_net_1125;
	wire new_net_1587;
	wire new_net_770;
	wire new_net_874;
	wire new_net_281;
	wire new_net_299;
	wire new_net_368;
	wire new_net_789;
	wire new_net_1306;
	wire new_net_1318;
	wire new_net_1343;
	wire new_net_1407;
	wire new_net_1516;
	wire _350_;
	wire new_net_351;
	wire _158_;
	wire _284_;
	wire new_net_9;
	wire new_net_315;
	wire new_net_333;
	wire new_net_93;
	wire new_net_534;
	wire new_net_892;
	wire new_net_904;
	wire new_net_1447;
	wire new_net_1152;
	wire new_net_1498;
	wire new_net_43;
	wire new_net_127;
	wire new_net_436;
	wire new_net_550;
	wire new_net_851;
	wire new_net_938;
	wire new_net_1100;
	wire new_net_1112;
	wire new_net_1485;
	wire new_net_1508;
	wire new_net_1728;
	wire new_net_1454;
	wire new_net_1476;
	wire new_net_470;
	wire _285_;
	wire _159_;
	wire new_net_230;
	wire new_net_248;
	wire new_net_566;
	wire new_net_518;
	wire new_net_1025;
	wire new_net_1037;
	wire new_net_1261;
	wire new_net_1650;
	wire new_net_1489;
	wire new_net_27;
	wire new_net_282;
	wire new_net_300;
	wire new_net_369;
	wire new_net_841;
	wire new_net_1002;
	wire new_net_1057;
	wire new_net_1069;
	wire new_net_1284;
	wire new_net_1326;
	wire new_net_1621;
	wire new_net_1705;
	wire new_net_1293;
	wire new_net_1669;
	wire new_net_403;
	wire new_net_535;
	wire new_net_352;
	wire _160_;
	wire _286_;
	wire new_net_10;
	wire new_net_487;
	wire new_net_959;
	wire new_net_1362;
	wire new_net_1374;
	wire new_net_1634;
	wire new_net_1350;
	wire new_net_1348;
	wire new_net_1607;
	wire new_net_976;
	wire new_net_44;
	wire new_net_110;
	wire new_net_128;
	wire new_net_551;
	wire new_net_731;
	wire new_net_1079;
	wire new_net_1216;
	wire new_net_1385;
	wire new_net_1242;
	wire new_net_1159;
	wire new_net_1376;
	wire new_net_567;
	wire new_net_771;
	wire new_net_875;
	wire new_net_519;
	wire new_net_471;
	wire _161_;
	wire _287_;
	wire new_net_231;
	wire new_net_249;
	wire new_net_653;
	wire new_net_1551;
	wire new_net_28;
	wire new_net_94;
	wire new_net_283;
	wire new_net_301;
	wire new_net_316;
	wire new_net_334;
	wire new_net_370;
	wire new_net_893;
	wire new_net_905;
	wire new_net_1045;
	wire new_net_1186;
	wire new_net_1655;
	wire new_net_488;
	wire new_net_437;
	wire new_net_852;
	wire _162_;
	wire _288_;
	wire new_net_11;
	wire new_net_404;
	wire new_net_353;
	wire new_net_939;
	wire new_net_1101;
	wire new_net_45;
	wire new_net_111;
	wire new_net_591;
	wire new_net_651;
	wire new_net_761;
	wire new_net_1026;
	wire new_net_1038;
	wire new_net_1262;
	wire new_net_1329;
	wire new_net_1341;
	wire new_net_1599;
	wire new_net_472;
	wire new_net_597;
	wire new_net_842;
	wire new_net_250;
	wire new_net_627;
	wire _289_;
	wire _163_;
	wire new_net_232;
	wire new_net_520;
	wire new_net_820;
	wire new_net_536;
	wire new_net_95;
	wire new_net_284;
	wire new_net_317;
	wire new_net_335;
	wire new_net_371;
	wire new_net_960;
	wire new_net_996;
	wire new_net_1164;
	wire new_net_1363;
	wire new_net_576;
	wire new_net_354;
	wire new_net_552;
	wire new_net_639;
	wire new_net_438;
	wire _164_;
	wire _290_;
	wire new_net_12;
	wire new_net_601;
	wire new_net_709;
	wire new_net_1463;
	wire new_net_1271;
	wire new_net_791;
	wire new_net_869;
	wire new_net_46;
	wire new_net_112;
	wire new_net_762;
	wire new_net_772;
	wire new_net_1308;
	wire new_net_1320;
	wire new_net_1409;
	wire new_net_1421;
	wire new_net_251;
	wire new_net_668;
	wire new_net_521;
	wire new_net_821;
	wire new_net_473;
	wire new_net_587;
	wire new_net_616;
	wire new_net_233;
	wire new_net_302;
	wire _165_;
	wire new_net_1137;
	wire new_net_1396;
	wire new_net_1604;
	wire new_net_568;
	wire new_net_853;
	wire new_net_537;
	wire new_net_655;
	wire new_net_96;
	wire new_net_285;
	wire new_net_318;
	wire new_net_336;
	wire new_net_372;
	wire new_net_405;
	wire new_net_988;
	wire new_net_1289;
	wire new_net_553;
	wire new_net_439;
	wire new_net_580;
	wire new_net_130;
	wire new_net_640;
	wire _166_;
	wire _292_;
	wire new_net_1027;
	wire new_net_1039;
	wire new_net_1213;
	wire new_net_1171;
	wire new_net_1380;
	wire new_net_1094;
	wire new_net_113;
	wire new_net_585;
	wire new_net_603;
	wire new_net_624;
	wire new_net_1004;
	wire new_net_1047;
	wire new_net_1059;
	wire new_net_1286;
	wire new_net_1455;
	wire new_net_1467;
	wire new_net_804;
	wire new_net_474;
	wire new_net_234;
	wire new_net_303;
	wire new_net_650;
	wire new_net_876;
	wire new_net_522;
	wire _167_;
	wire _293_;
	wire new_net_30;
	wire new_net_961;
	wire new_net_129;
	wire new_net_1542;
	wire new_net_209;
	wire new_net_490;
	wire new_net_733;
	wire new_net_13;
	wire new_net_97;
	wire new_net_319;
	wire new_net_337;
	wire new_net_355;
	wire new_net_406;
	wire new_net_1081;
	wire new_net_1218;
	wire new_net_1431;
	wire _352_;
	wire new_net_1564;
	wire new_net_792;
	wire new_net_554;
	wire new_net_440;
	wire new_net_763;
	wire _294_;
	wire _000_;
	wire _168_;
	wire new_net_47;
	wire new_net_1309;
	wire new_net_1321;
	wire new_net_310;
	wire new_net_822;
	wire new_net_114;
	wire new_net_252;
	wire new_net_267;
	wire new_net_578;
	wire new_net_607;
	wire new_net_895;
	wire new_net_907;
	wire new_net_1465;
	wire new_net_1589;
	wire new_net_1458;
	wire new_net_1382;
	wire _001_;
	wire _295_;
	wire _169_;
	wire new_net_523;
	wire new_net_286;
	wire new_net_538;
	wire new_net_235;
	wire new_net_373;
	wire new_net_843;
	wire new_net_917;
	wire new_net_1729;
	wire new_net_1521;
	wire new_net_14;
	wire new_net_98;
	wire new_net_131;
	wire new_net_320;
	wire new_net_338;
	wire new_net_356;
	wire new_net_407;
	wire new_net_857;
	wire new_net_579;
	wire new_net_1028;
	wire new_net_1414;
	wire new_net_1332;
	wire new_net_915;
	wire new_net_1080;
	wire new_net_1507;
	wire new_net_1547;
	wire _002_;
	wire _296_;
	wire _170_;
	wire new_net_48;
	wire new_net_441;
	wire new_net_667;
	wire new_net_555;
	wire new_net_1005;
	wire new_net_1048;
	wire new_net_1060;
	wire new_net_1267;
	wire new_net_1436;
	wire new_net_31;
	wire new_net_115;
	wire new_net_253;
	wire new_net_304;
	wire new_net_475;
	wire new_net_582;
	wire new_net_641;
	wire new_net_962;
	wire new_net_1353;
	wire new_net_1365;
	wire new_net_1576;
	wire new_net_1533;
	wire new_net_1035;
	wire new_net_1033;
	wire _297_;
	wire _003_;
	wire _171_;
	wire new_net_491;
	wire new_net_374;
	wire new_net_711;
	wire new_net_287;
	wire new_net_539;
	wire new_net_1082;
	wire new_net_1219;
	wire new_net_1253;
	wire new_net_925;
	wire new_net_1470;
	wire new_net_1674;
	wire new_net_1387;
	wire new_net_15;
	wire new_net_99;
	wire new_net_132;
	wire new_net_321;
	wire new_net_339;
	wire new_net_408;
	wire new_net_764;
	wire new_net_1223;
	wire new_net_1310;
	wire new_net_1322;
	wire new_net_1560;
	wire new_net_1639;
	wire new_net_823;
	wire _298_;
	wire _004_;
	wire _172_;
	wire new_net_573;
	wire new_net_442;
	wire new_net_581;
	wire new_net_896;
	wire new_net_908;
	wire new_net_1590;
	wire new_net_1001;
	wire new_net_1339;
	wire new_net_32;
	wire new_net_236;
	wire new_net_305;
	wire new_net_476;
	wire new_net_524;
	wire new_net_571;
	wire new_net_586;
	wire new_net_614;
	wire new_net_659;
	wire new_net_918;
	wire new_net_1512;
	wire new_net_1302;
	wire _353_;
	wire new_net_1443;
	wire _299_;
	wire _173_;
	wire _005_;
	wire new_net_288;
	wire new_net_357;
	wire new_net_492;
	wire new_net_654;
	wire new_net_1029;
	wire new_net_1041;
	wire new_net_1265;
	wire new_net_1494;
	wire new_net_1538;
	wire new_net_16;
	wire new_net_49;
	wire new_net_133;
	wire new_net_340;
	wire new_net_409;
	wire new_net_556;
	wire new_net_652;
	wire new_net_1006;
	wire new_net_1040;
	wire new_net_1049;
	wire new_net_254;
	wire new_net_877;
	wire _006_;
	wire _174_;
	wire _300_;
	wire new_net_116;
	wire new_net_844;
	wire new_net_963;
	wire new_net_1354;
	wire new_net_1366;
	wire new_net_1392;
	wire new_net_1644;
	wire new_net_33;
	wire new_net_237;
	wire new_net_375;
	wire new_net_525;
	wire new_net_540;
	wire new_net_592;
	wire new_net_628;
	wire new_net_662;
	wire new_net_1083;
	wire new_net_1220;
	wire new_net_1617;
	wire new_net_1699;
	wire new_net_1665;
	wire new_net_1588;
	wire new_net_1209;
	wire new_net_358;
	wire new_net_765;
	wire _301_;
	wire _007_;
	wire _175_;
	wire new_net_322;
	wire new_net_100;
	wire new_net_289;
	wire new_net_1311;
	wire new_net_1323;
	wire new_net_1426;
	wire new_net_1344;
	wire new_net_1710;
	wire new_net_17;
	wire new_net_50;
	wire new_net_134;
	wire new_net_410;
	wire new_net_443;
	wire new_net_557;
	wire new_net_824;
	wire new_net_897;
	wire new_net_909;
	wire new_net_1591;
	wire new_net_1448;
	wire new_net_1113;
	wire new_net_1153;
	wire new_net_1370;
	wire new_net_477;
	wire _302_;
	wire _008_;
	wire _176_;
	wire new_net_117;
	wire new_net_306;
	wire new_net_255;
	wire new_net_919;
	wire new_net_1105;
	wire new_net_1117;
	wire new_net_888;
	wire new_net_34;
	wire new_net_376;
	wire new_net_493;
	wire new_net_541;
	wire new_net_583;
	wire new_net_664;
	wire new_net_734;
	wire new_net_773;
	wire new_net_1030;
	wire new_net_1042;
	wire new_net_1182;
	wire new_net_1477;
	wire new_net_1651;
	wire new_net_1490;
	wire new_net_341;
	wire new_net_615;
	wire new_net_101;
	wire new_net_290;
	wire _009_;
	wire _177_;
	wire _303_;
	wire new_net_881;
	wire new_net_323;
	wire new_net_1007;
	wire new_net_955;
	wire new_net_916;
	wire new_net_18;
	wire new_net_51;
	wire new_net_444;
	wire new_net_870;
	wire new_net_964;
	wire new_net_1355;
	wire new_net_1367;
	wire new_net_1612;
	wire new_net_1666;
	wire new_net_1735;
	wire _354_;
	wire new_net_713;
	wire new_net_774;
	wire new_net_526;
	wire _010_;
	wire _178_;
	wire _304_;
	wire new_net_478;
	wire new_net_238;
	wire new_net_307;
	wire new_net_1072;
	wire new_net_1608;
	wire new_net_1733;
	wire new_net_735;
	wire new_net_878;
	wire new_net_35;
	wire new_net_359;
	wire new_net_494;
	wire new_net_1312;
	wire new_net_1324;
	wire new_net_1413;
	wire new_net_1425;
	wire new_net_1552;
	wire new_net_1725;
	wire new_net_558;
	wire new_net_825;
	wire new_net_324;
	wire _305_;
	wire _011_;
	wire _179_;
	wire new_net_135;
	wire new_net_342;
	wire new_net_411;
	wire new_net_793;
	wire new_net_426;
	wire new_net_19;
	wire new_net_52;
	wire new_net_118;
	wire new_net_256;
	wire new_net_845;
	wire new_net_920;
	wire new_net_1106;
	wire new_net_1118;
	wire new_net_1491;
	wire new_net_1514;
	wire new_net_1629;
	wire new_net_1627;
	wire new_net_479;
	wire new_net_542;
	wire new_net_669;
	wire new_net_377;
	wire _012_;
	wire _180_;
	wire _306_;
	wire new_net_239;
	wire new_net_642;
	wire new_net_527;
	wire new_net_1299;
	wire new_net_1133;
	wire new_net_1600;
	wire new_net_794;
	wire new_net_36;
	wire new_net_102;
	wire new_net_360;
	wire new_net_596;
	wire new_net_632;
	wire new_net_1008;
	wire new_net_1051;
	wire new_net_1063;
	wire new_net_1290;
	wire new_net_834;
	wire new_net_984;
	wire new_net_1613;
	wire new_net_1285;
	wire new_net_343;
	wire new_net_412;
	wire new_net_559;
	wire _181_;
	wire _013_;
	wire _307_;
	wire new_net_136;
	wire new_net_445;
	wire new_net_325;
	wire new_net_965;
	wire new_net_1167;
	wire new_net_997;
	wire new_net_1165;
	wire new_net_611;
	wire new_net_1090;
	wire new_net_1307;
	wire new_net_775;
	wire new_net_20;
	wire new_net_53;
	wire new_net_119;
	wire new_net_257;
	wire new_net_308;
	wire new_net_1073;
	wire new_net_1085;
	wire new_net_1222;
	wire new_net_1379;
	wire new_net_168;
	wire new_net_1194;
	wire new_net_1405;
	wire new_net_736;
	wire new_net_879;
	wire new_net_480;
	wire new_net_543;
	wire new_net_575;
	wire _182_;
	wire _014_;
	wire _308_;
	wire new_net_378;
	wire new_net_495;
	wire new_net_1074;
	wire new_net_1720;
	wire new_net_666;
	wire new_net_826;
	wire new_net_103;
	wire new_net_292;
	wire new_net_361;
	wire new_net_899;
	wire new_net_911;
	wire new_net_941;
	wire new_net_1593;
	wire new_net_1605;
	wire new_net_1397;
	wire new_net_1711;
	wire new_net_446;
	wire new_net_846;
	wire new_net_137;
	wire new_net_344;
	wire _183_;
	wire _015_;
	wire _309_;
	wire new_net_921;
	wire new_net_1107;
	wire new_net_1119;
	wire new_net_657;
	wire new_net_54;
	wire new_net_120;
	wire new_net_240;
	wire new_net_309;
	wire new_net_528;
	wire new_net_645;
	wire new_net_1032;
	wire new_net_1044;
	wire new_net_1268;
	wire new_net_1381;
	wire new_net_795;
	wire new_net_496;
	wire _184_;
	wire _016_;
	wire _310_;
	wire new_net_37;
	wire new_net_1009;
	wire new_net_1052;
	wire new_net_1064;
	wire new_net_1291;
	wire new_net_1517;
	wire new_net_871;
	wire new_net_293;
	wire new_net_326;
	wire new_net_362;
	wire new_net_413;
	wire new_net_560;
	wire new_net_942;
	wire new_net_966;
	wire new_net_1357;
	wire new_net_1369;
	wire new_net_1410;
	wire new_net_1721;
	wire new_net_1328;
	wire new_net_1543;
	wire new_net_345;
	wire new_net_626;
	wire new_net_649;
	wire new_net_258;
	wire new_net_715;
	wire _185_;
	wire _017_;
	wire _311_;
	wire new_net_21;
	wire new_net_138;
	wire new_net_1263;
	wire new_net_1432;
	wire new_net_1145;
	wire new_net_880;
	wire new_net_121;
	wire new_net_241;
	wire new_net_379;
	wire new_net_481;
	wire new_net_529;
	wire new_net_544;
	wire new_net_737;
	wire new_net_1314;
	wire new_net_1415;
	wire new_net_1565;
	wire new_net_732;
	wire new_net_665;
	wire new_net_827;
	wire new_net_104;
	wire _018_;
	wire _186_;
	wire _312_;
	wire new_net_38;
	wire new_net_900;
	wire new_net_912;
	wire new_net_1594;
	wire new_net_1724;
	wire new_net_1466;
	wire new_net_1459;
	wire new_net_327;
	wire new_net_363;
	wire new_net_414;
	wire new_net_447;
	wire new_net_151;
	wire new_net_561;
	wire new_net_847;
	wire new_net_922;
	wire new_net_1108;
	wire new_net_1120;
	wire new_net_1688;
	wire new_net_55;
	wire new_net_766;
	wire new_net_259;
	wire new_net_574;
	wire new_net_139;
	wire new_net_346;
	wire new_net_717;
	wire _019_;
	wire _187_;
	wire _313_;
	wire new_net_63;
	wire new_net_195;
	wire new_net_1417;
	wire new_net_1333;
	wire new_net_497;
	wire new_net_872;
	wire new_net_545;
	wire new_net_122;
	wire new_net_242;
	wire new_net_380;
	wire new_net_482;
	wire new_net_796;
	wire new_net_1010;
	wire new_net_1053;
	wire new_net_1548;
	wire new_net_218;
	wire new_net_1439;
	wire new_net_1437;
	wire new_net_644;
	wire _020_;
	wire _188_;
	wire _314_;
	wire new_net_105;
	wire new_net_294;
	wire new_net_943;
	wire new_net_940;
	wire new_net_1102;
	wire new_net_1358;
	wire new_net_1731;
	wire new_net_1577;
	wire new_net_1570;
	wire new_net_1534;
	wire new_net_619;
	wire new_net_777;
	wire new_net_328;
	wire new_net_364;
	wire new_net_415;
	wire new_net_448;
	wire new_net_584;
	wire new_net_589;
	wire new_net_647;
	wire new_net_1075;
	wire new_net_1723;
	wire new_net_1471;
	wire new_net_91;
	wire new_net_1675;
	wire new_net_718;
	wire new_net_311;
	wire new_net_767;
	wire new_net_738;
	wire new_net_140;
	wire new_net_530;
	wire _189_;
	wire _021_;
	wire _315_;
	wire new_net_56;
	wire new_net_1388;
	wire new_net_1561;
	wire new_net_1640;
	wire new_net_1067;
	wire new_net_1065;
	wire new_net_868;
	wire new_net_1319;
	wire new_net_828;
	wire new_net_39;
	wire new_net_123;
	wire new_net_243;
	wire new_net_381;
	wire new_net_498;
	wire new_net_901;
	wire new_net_913;
	wire new_net_1595;
	wire new_net_1695;
	wire new_net_1661;
	wire new_net_1205;
	wire new_net_1422;
	wire new_net_1340;
	wire new_net_1453;
	wire new_net_1086;
	wire new_net_968;
	wire new_net_1513;
	wire new_net_1303;
	wire new_net_1444;
	wire _022_;
	wire _064_;
	wire _106_;
	wire _190_;
	wire _232_;
	wire _316_;
	wire _358_;
	wire new_net_157;
	wire new_net_208;
	wire new_net_923;
	wire new_net_1149;
	wire new_net_260;
	wire new_net_416;
	wire new_net_449;
	wire new_net_599;
	wire new_net_643;
	wire new_net_1132;
	wire new_net_1144;
	wire new_net_1270;
	wire new_net_1178;
	wire new_net_1176;
	wire _023_;
	wire _065_;
	wire _107_;
	wire _191_;
	wire _233_;
	wire _317_;
	wire _359_;
	wire new_net_621;
	wire new_net_1011;
	wire new_net_1155;
	wire new_net_1393;
	wire new_net_1486;
	wire new_net_1645;
	wire new_net_1718;
	wire new_net_73;
	wire new_net_175;
	wire new_net_193;
	wire new_net_382;
	wire new_net_944;
	wire new_net_1616;
	wire new_net_1628;
	wire new_net_1670;
	wire new_net_1700;
	wire new_net_1127;
	wire new_net_1427;
	wire _192_;
	wire _234_;
	wire _024_;
	wire _066_;
	wire _108_;
	wire _318_;
	wire _360_;
	wire new_net_158;
	wire new_net_693;
	wire new_net_778;
	wire new_net_1345;
	wire _357_;
	wire new_net_57;
	wire new_net_141;
	wire new_net_261;
	wire new_net_450;
	wire new_net_719;
	wire new_net_979;
	wire new_net_991;
	wire new_net_1449;
	wire new_net_1114;
	wire _291_;
	wire _193_;
	wire _235_;
	wire _025_;
	wire _067_;
	wire _109_;
	wire _319_;
	wire _361_;
	wire new_net_829;
	wire new_net_499;
	wire new_net_1236;
	wire new_net_1500;
	wire new_net_1556;
	wire new_net_74;
	wire new_net_383;
	wire new_net_681;
	wire new_net_924;
	wire new_net_1478;
	wire new_net_1495;
	wire new_net_1518;
	wire new_net_1652;
	wire _194_;
	wire _236_;
	wire _026_;
	wire _068_;
	wire _110_;
	wire _320_;
	wire new_net_210;
	wire new_net_417;
	wire new_net_159;
	wire new_net_967;
	wire new_net_1623;
	wire new_net_1295;
	wire new_net_1596;
	wire new_net_58;
	wire new_net_142;
	wire new_net_262;
	wire new_net_451;
	wire new_net_1012;
	wire new_net_1156;
	wire new_net_1168;
	wire new_net_1224;
	wire new_net_1294;
	wire new_net_1540;
	wire new_net_980;
	wire new_net_1609;
	wire new_net_978;
	wire new_net_176;
	wire new_net_500;
	wire _027_;
	wire _069_;
	wire _111_;
	wire _195_;
	wire _237_;
	wire _321_;
	wire new_net_194;
	wire new_net_945;
	wire new_net_1281;
	wire new_net_1451;
	wire new_net_1161;
	wire new_net_384;
	wire new_net_779;
	wire new_net_1089;
	wire new_net_1179;
	wire new_net_1191;
	wire new_net_1202;
	wire new_net_1395;
	wire new_net_1563;
	wire new_net_1575;
	wire new_net_1706;
	wire new_net_1553;
	wire new_net_418;
	wire new_net_862;
	wire new_net_720;
	wire _196_;
	wire _238_;
	wire _028_;
	wire _070_;
	wire _112_;
	wire _322_;
	wire new_net_211;
	wire new_net_1190;
	wire new_net_1188;
	wire new_net_263;
	wire new_net_452;
	wire new_net_830;
	wire new_net_1225;
	wire new_net_1237;
	wire new_net_1249;
	wire new_net_1692;
	wire new_net_1704;
	wire new_net_625;
	wire _239_;
	wire _029_;
	wire _071_;
	wire _113_;
	wire _197_;
	wire _323_;
	wire new_net_75;
	wire new_net_808;
	wire new_net_177;
	wire new_net_1601;
	wire new_net_739;
	wire new_net_160;
	wire new_net_682;
	wire new_net_797;
	wire new_net_1134;
	wire new_net_1146;
	wire new_net_1272;
	wire new_net_1614;
	wire new_net_143;
	wire _030_;
	wire _072_;
	wire _114_;
	wire _198_;
	wire _240_;
	wire _324_;
	wire new_net_59;
	wire new_net_1013;
	wire new_net_1157;
	wire new_net_264;
	wire new_net_453;
	wire new_net_501;
	wire new_net_672;
	wire new_net_946;
	wire new_net_1618;
	wire new_net_1630;
	wire new_net_1672;
	wire new_net_1273;
	wire new_net_1479;
	wire new_net_1195;
	wire new_net_1406;
	wire new_net_1719;
	wire new_net_695;
	wire new_net_385;
	wire new_net_598;
	wire _031_;
	wire _073_;
	wire _115_;
	wire _199_;
	wire _241_;
	wire _325_;
	wire new_net_76;
	wire new_net_1539;
	wire new_net_1259;
	wire new_net_809;
	wire new_net_161;
	wire new_net_212;
	wire new_net_419;
	wire new_net_612;
	wire new_net_740;
	wire new_net_863;
	wire new_net_883;
	wire new_net_969;
	wire new_net_981;
	wire new_net_1139;
	wire new_net_1398;
	wire _032_;
	wire _074_;
	wire _116_;
	wire _200_;
	wire _242_;
	wire _326_;
	wire new_net_60;
	wire new_net_144;
	wire new_net_1226;
	wire new_net_1238;
	wire new_net_992;
	wire new_net_990;
	wire new_net_1462;
	wire new_net_178;
	wire new_net_196;
	wire new_net_265;
	wire new_net_454;
	wire new_net_502;
	wire new_net_926;
	wire new_net_1497;
	wire new_net_1520;
	wire new_net_1215;
	wire new_net_1056;
	wire new_net_1096;
	wire _075_;
	wire _033_;
	wire _117_;
	wire _201_;
	wire _243_;
	wire _327_;
	wire new_net_386;
	wire new_net_602;
	wire new_net_1123;
	wire new_net_1135;
	wire new_net_1313;
	wire new_net_1716;
	wire new_net_162;
	wire new_net_213;
	wire new_net_420;
	wire new_net_683;
	wire new_net_1014;
	wire new_net_1158;
	wire new_net_1170;
	wire new_net_1199;
	wire new_net_1296;
	wire new_net_1411;
	wire new_net_460;
	wire new_net_646;
	wire new_net_673;
	wire _034_;
	wire _076_;
	wire _118_;
	wire _202_;
	wire _244_;
	wire _328_;
	wire new_net_61;
	wire new_net_947;
	wire new_net_1264;
	wire new_net_1433;
	wire new_net_781;
	wire new_net_77;
	wire new_net_179;
	wire new_net_197;
	wire new_net_751;
	wire new_net_799;
	wire new_net_1091;
	wire new_net_1181;
	wire new_net_1193;
	wire new_net_1204;
	wire new_net_1566;
	wire new_net_387;
	wire new_net_741;
	wire _035_;
	wire _077_;
	wire _119_;
	wire _203_;
	wire _245_;
	wire _329_;
	wire new_net_636;
	wire new_net_884;
	wire new_net_1460;
	wire new_net_1671;
	wire new_net_1384;
	wire new_net_1557;
	wire new_net_1636;
	wire new_net_569;
	wire new_net_145;
	wire new_net_163;
	wire new_net_214;
	wire new_net_421;
	wire new_net_1227;
	wire new_net_1239;
	wire new_net_1682;
	wire new_net_1694;
	wire new_net_1061;
	wire new_net_1475;
	wire new_net_1523;
	wire new_net_1717;
	wire new_net_1691;
	wire new_net_1689;
	wire new_net_1277;
	wire new_net_503;
	wire new_net_266;
	wire new_net_455;
	wire _204_;
	wire _246_;
	wire _036_;
	wire _078_;
	wire _120_;
	wire _330_;
	wire new_net_62;
	wire new_net_1201;
	wire new_net_1418;
	wire new_net_1416;
	wire new_net_1334;
	wire new_net_1509;
	wire new_net_1549;
	wire new_net_78;
	wire new_net_180;
	wire new_net_721;
	wire new_net_1124;
	wire new_net_1136;
	wire new_net_1274;
	wire new_net_750;
	wire new_net_790;
	wire new_net_1440;
	wire new_net_1269;
	wire new_net_1438;
	wire new_net_722;
	wire new_net_388;
	wire new_net_631;
	wire _205_;
	wire _247_;
	wire _037_;
	wire _079_;
	wire _121_;
	wire _331_;
	wire new_net_1015;
	wire new_net_1103;
	wire new_net_1714;
	wire new_net_1578;
	wire new_net_1535;
	wire new_net_1019;
	wire new_net_810;
	wire new_net_684;
	wire new_net_146;
	wire new_net_164;
	wire new_net_215;
	wire new_net_422;
	wire new_net_882;
	wire new_net_948;
	wire new_net_1377;
	wire new_net_1620;
	wire new_net_1255;
	wire new_net_1504;
	wire new_net_927;
	wire new_net_1472;
	wire new_net_613;
	wire new_net_752;
	wire new_net_800;
	wire new_net_504;
	wire new_net_570;
	wire new_net_697;
	wire _038_;
	wire _080_;
	wire _122_;
	wire _206_;
	wire new_net_1389;
	wire new_net_1482;
	wire new_net_1641;
	wire new_net_1068;
	wire new_net_1668;
	wire new_net_181;
	wire new_net_742;
	wire new_net_971;
	wire new_net_983;
	wire new_net_1147;
	wire new_net_1250;
	wire new_net_1662;
	wire new_net_1206;
	wire new_net_1003;
	wire new_net_1423;
	wire new_net_674;
	wire _039_;
	wire _081_;
	wire _123_;
	wire _207_;
	wire _249_;
	wire _333_;
	wire new_net_1228;
	wire new_net_1240;
	wire new_net_1683;
	wire new_net_1087;
	wire new_net_291;
	wire new_net_831;
	wire new_net_165;
	wire new_net_216;
	wire new_net_423;
	wire new_net_928;
	wire new_net_1445;
	wire new_net_1499;
	wire new_net_1522;
	wire new_net_1110;
	wire new_net_507;
	wire new_net_1496;
	wire new_net_199;
	wire new_net_854;
	wire _208_;
	wire _250_;
	wire _040_;
	wire _082_;
	wire _124_;
	wire _334_;
	wire new_net_64;
	wire new_net_79;
	wire new_net_1402;
	wire new_net_1592;
	wire new_net_1726;
	wire new_net_1474;
	wire new_net_182;
	wire new_net_389;
	wire new_net_634;
	wire new_net_811;
	wire new_net_1016;
	wire new_net_1148;
	wire new_net_1160;
	wire new_net_1172;
	wire new_net_1298;
	wire new_net_1544;
	wire new_net_1648;
	wire new_net_489;
	wire new_net_1487;
	wire new_net_1480;
	wire new_net_1646;
	wire _209_;
	wire _251_;
	wire _041_;
	wire _083_;
	wire _125_;
	wire _335_;
	wire new_net_147;
	wire new_net_885;
	wire new_net_949;
	wire new_net_1325;
	wire new_net_1619;
	wire new_net_1703;
	wire new_net_1701;
	wire new_net_1667;
	wire new_net_753;
	wire new_net_801;
	wire new_net_505;
	wire new_net_600;
	wire new_net_457;
	wire new_net_217;
	wire new_net_268;
	wire new_net_424;
	wire new_net_1093;
	wire new_net_1183;
	wire new_net_1211;
	wire new_net_1632;
	wire new_net_1346;
	wire new_net_974;
	wire new_net_80;
	wire new_net_743;
	wire _210_;
	wire _252_;
	wire _042_;
	wire _084_;
	wire _126_;
	wire _336_;
	wire new_net_898;
	wire new_net_972;
	wire new_net_1450;
	wire new_net_1115;
	wire new_net_832;
	wire new_net_629;
	wire new_net_183;
	wire new_net_390;
	wire new_net_620;
	wire new_net_1229;
	wire new_net_1241;
	wire new_net_1276;
	wire new_net_1684;
	wire new_net_1696;
	wire _043_;
	wire _085_;
	wire _127_;
	wire _211_;
	wire _253_;
	wire _337_;
	wire new_net_148;
	wire new_net_166;
	wire new_net_929;
	wire new_net_1184;
	wire new_net_1653;
	wire new_net_1492;
	wire new_net_65;
	wire new_net_200;
	wire new_net_269;
	wire new_net_506;
	wire new_net_458;
	wire new_net_605;
	wire new_net_675;
	wire new_net_728;
	wire new_net_1126;
	wire new_net_1138;
	wire _212_;
	wire _254_;
	wire _044_;
	wire _086_;
	wire _128_;
	wire _338_;
	wire new_net_572;
	wire new_net_782;
	wire new_net_617;
	wire new_net_1017;
	wire new_net_595;
	wire new_net_687;
	wire new_net_950;
	wire new_net_1622;
	wire new_net_1676;
	wire new_net_1712;
	wire new_net_1610;
	wire new_net_1530;
	wire new_net_1282;
	wire new_net_1452;
	wire new_net_425;
	wire _213_;
	wire _255_;
	wire _045_;
	wire _087_;
	wire _129_;
	wire _339_;
	wire new_net_149;
	wire new_net_167;
	wire new_net_723;
	wire new_net_1554;
	wire new_net_66;
	wire new_net_81;
	wire new_net_201;
	wire new_net_973;
	wire new_net_985;
	wire new_net_993;
	wire _214_;
	wire _256_;
	wire _046_;
	wire _088_;
	wire _130_;
	wire _340_;
	wire new_net_184;
	wire new_net_660;
	wire new_net_391;
	wire new_net_812;
	wire new_net_930;
	wire new_net_1501;
	wire new_net_1524;
	wire new_net_1394;
	wire new_net_1602;
	wire new_net_270;
	wire new_net_459;
	wire _047_;
	wire _089_;
	wire _131_;
	wire _215_;
	wire _257_;
	wire _341_;
	wire new_net_150;
	wire new_net_219;
	wire new_net_986;
	wire new_net_1615;
	wire new_net_910;
	wire new_net_1287;
	wire new_net_82;
	wire new_net_676;
	wire new_net_833;
	wire new_net_994;
	wire new_net_1018;
	wire new_net_1150;
	wire new_net_1162;
	wire new_net_1300;
	wire new_net_1546;
	wire new_net_1709;
	wire new_net_1169;
	wire new_net_1378;
	wire new_net_1092;
	wire new_net_1050;
	wire new_net_185;
	wire new_net_392;
	wire _048_;
	wire _090_;
	wire _132_;
	wire _216_;
	wire _258_;
	wire _342_;
	wire new_net_886;
	wire new_net_951;
	wire new_net_802;
	wire new_net_1196;
	wire new_net_803;
	wire new_net_724;
	wire new_net_1095;
	wire new_net_1185;
	wire new_net_1197;
	wire new_net_1208;
	wire new_net_1401;
	wire new_net_1569;
	wire new_net_1631;
	wire new_net_169;
	wire _049_;
	wire _091_;
	wire _133_;
	wire _217_;
	wire _259_;
	wire _343_;
	wire new_net_67;
	wire new_net_508;
	wire new_net_202;
	wire new_net_1429;
	wire new_net_1562;
	wire new_net_1399;
	wire new_net_83;
	wire new_net_685;
	wire new_net_813;
	wire new_net_1231;
	wire new_net_1243;
	wire new_net_1686;
	wire new_net_1698;
	wire _050_;
	wire _092_;
	wire _134_;
	wire _218_;
	wire _260_;
	wire _344_;
	wire new_net_186;
	wire new_net_931;
	wire new_net_1173;
	wire new_net_1292;
	wire new_net_1456;
	wire new_net_744;
	wire new_net_855;
	wire new_net_754;
	wire new_net_0;
	wire new_net_220;
	wire new_net_427;
	wire new_net_671;
	wire new_net_1128;
	wire new_net_1140;
	wire new_net_1254;
	wire new_net_1519;
	wire new_net_1685;
	wire new_net_203;
	wire new_net_749;
	wire new_net_152;
	wire _051_;
	wire _093_;
	wire _135_;
	wire _219_;
	wire _261_;
	wire _345_;
	wire new_net_68;
	wire new_net_699;
	wire new_net_1412;
	wire new_net_1330;
	wire new_net_1078;
	wire new_net_1505;
	wire new_net_1545;
	wire new_net_84;
	wire new_net_393;
	wire new_net_677;
	wire new_net_689;
	wire new_net_858;
	wire new_net_952;
	wire new_net_1624;
	wire new_net_1678;
	wire new_net_1434;
	wire new_net_701;
	wire _220_;
	wire _262_;
	wire _052_;
	wire _094_;
	wire _136_;
	wire _346_;
	wire new_net_187;
	wire new_net_593;
	wire new_net_725;
	wire new_net_1356;
	wire new_net_1574;
	wire new_net_1567;
	wire new_net_1531;
	wire new_net_1734;
	wire new_net_1031;
	wire new_net_1581;
	wire new_net_509;
	wire new_net_1;
	wire new_net_170;
	wire new_net_221;
	wire new_net_272;
	wire new_net_428;
	wire new_net_461;
	wire new_net_745;
	wire new_net_755;
	wire new_net_887;
	wire new_net_1251;
	wire new_net_780;
	wire new_net_1468;
	wire new_net_1461;
	wire new_net_1221;
	wire new_net_1558;
	wire new_net_1637;
	wire new_net_814;
	wire _221_;
	wire _263_;
	wire _053_;
	wire _095_;
	wire _137_;
	wire _347_;
	wire new_net_1232;
	wire new_net_1244;
	wire new_net_1687;
	wire new_net_1062;
	wire new_net_1690;
	wire new_net_85;
	wire new_net_394;
	wire new_net_932;
	wire new_net_1503;
	wire new_net_1278;
	wire new_net_1526;
	wire new_net_1633;
	wire new_net_1730;
	wire new_net_1419;
	wire new_net_1335;
	wire _054_;
	wire _096_;
	wire _138_;
	wire _222_;
	wire _264_;
	wire _348_;
	wire new_net_608;
	wire new_net_783;
	wire new_net_1129;
	wire new_net_1141;
	wire new_net_1510;
	wire new_net_1550;
	wire new_net_29;
	wire new_net_1441;
	wire new_net_861;
	wire new_net_835;
	wire new_net_69;
	wire new_net_153;
	wire new_net_171;
	wire new_net_204;
	wire new_net_222;
	wire new_net_273;
	wire new_net_510;
	wire new_net_462;
	wire new_net_1104;
	wire new_net_1403;
	wire new_net_1579;
	wire new_net_1572;
	wire new_net_1536;
	wire _055_;
	wire _097_;
	wire _139_;
	wire _223_;
	wire _265_;
	wire _349_;
	wire new_net_953;
	wire new_net_1625;
	wire new_net_1679;
	wire new_net_271;
	wire new_net_1473;
	wire new_net_188;
	wire new_net_618;
	wire new_net_678;
	wire new_net_726;
	wire new_net_805;
	wire new_net_1175;
	wire new_net_1187;
	wire new_net_1210;
	wire new_net_1571;
	wire new_net_1677;
	wire new_net_1390;
	wire new_net_1297;
	wire new_net_1483;
	wire new_net_1642;
	wire _248_;
	wire new_net_746;
	wire new_net_784;
	wire new_net_859;
	wire new_net_429;
	wire new_net_756;
	wire _224_;
	wire _266_;
	wire _056_;
	wire _098_;
	wire _140_;
	wire new_net_1071;
	wire new_net_1697;
	wire new_net_1663;
	wire new_net_1586;
	wire new_net_1207;
	wire new_net_815;
	wire new_net_70;
	wire new_net_154;
	wire new_net_205;
	wire new_net_223;
	wire new_net_274;
	wire new_net_511;
	wire new_net_1233;
	wire new_net_1245;
	wire new_net_1342;
	wire new_net_1424;
	wire new_net_970;
	wire new_net_1515;
	wire new_net_894;
	wire new_net_395;
	wire _225_;
	wire _267_;
	wire _057_;
	wire _099_;
	wire _141_;
	wire _351_;
	wire new_net_86;
	wire new_net_933;
	wire new_net_1527;
	wire new_net_1722;
	wire new_net_1446;
	wire new_net_1234;
	wire new_net_1111;
	wire new_net_1151;
	wire new_net_1368;
	wire new_net_2;
	wire new_net_189;
	wire new_net_1020;
	wire new_net_1130;
	wire new_net_1142;
	wire new_net_1198;
	wire new_net_1256;
	wire new_net_1301;
	wire new_net_1715;
	wire new_net_1043;
	wire new_net_1180;
	wire new_net_430;
	wire new_net_172;
	wire new_net_836;
	wire new_net_656;
	wire new_net_463;
	wire _226_;
	wire _268_;
	wire _142_;
	wire _058_;
	wire _100_;
	wire new_net_1649;
	wire new_net_1488;
	wire new_net_1481;
	wire new_net_1647;
	wire new_net_610;
	wire new_net_864;
	wire new_net_224;
	wire new_net_275;
	wire new_net_512;
	wire new_net_954;
	wire new_net_1626;
	wire new_net_1680;
	wire new_net_1702;
	wire new_net_87;
	wire new_net_691;
	wire new_net_727;
	wire new_net_703;
	wire new_net_806;
	wire _059_;
	wire _101_;
	wire _227_;
	wire _269_;
	wire _143_;
	wire new_net_1349;
	wire new_net_1347;
	wire new_net_1351;
	wire new_net_975;
	wire new_net_747;
	wire new_net_785;
	wire new_net_679;
	wire new_net_860;
	wire new_net_757;
	wire new_net_190;
	wire new_net_590;
	wire new_net_889;
	wire new_net_977;
	wire new_net_989;
	wire new_net_1116;
	wire new_net_71;
	wire new_net_206;
	wire new_net_464;
	wire new_net_816;
	wire new_net_155;
	wire new_net_173;
	wire _228_;
	wire _270_;
	wire _060_;
	wire _102_;
	wire new_net_1375;
	wire new_net_396;
	wire new_net_1502;
	wire new_net_3;
	wire new_net_225;
	wire new_net_276;
	wire new_net_934;
	wire new_net_1528;
	wire new_net_1635;
	wire new_net_397;
	wire _229_;
	wire _271_;
	wire _061_;
	wire _103_;
	wire _145_;
	wire _355_;
	wire new_net_1021;
	wire new_net_1131;
	wire new_net_1143;
	wire new_net_1493;
	wire new_net_1654;
	wire new_net_837;
	wire new_net_594;
	wire new_net_622;
	wire new_net_191;
	wire new_net_431;
	wire new_net_776;
	wire new_net_998;
	wire new_net_1154;
	wire new_net_1166;
	wire new_net_1280;
	wire new_net_1707;
	wire new_net_1598;
	wire new_net_513;
	wire new_net_207;
	wire new_net_156;
	wire _230_;
	wire _272_;
	wire _146_;
	wire _062_;
	wire _104_;
	wire _356_;
	wire new_net_72;
	wire new_net_982;
	wire new_net_1529;
	wire new_net_1611;
	wire new_net_906;
	wire new_net_1283;
	wire new_net_1248;
	wire new_net_807;
	wire new_net_4;
	wire new_net_88;
	wire new_net_277;
	wire new_net_1177;
	wire _144_;
	wire new_net_1189;
	wire new_net_1200;
	wire new_net_1212;
	wire new_net_1246;
	wire new_net_995;
	wire new_net_1163;
	wire new_net_1582;
	wire new_net_609;
	wire new_net_1088;
	wire new_net_1046;
	wire new_net_1555;
	wire new_net_1305;
	wire new_net_748;
	wire new_net_786;
	wire new_net_758;
	wire new_net_865;
	wire new_net_398;
	wire _231_;
	wire _273_;
	wire _147_;
	wire _063_;
	wire _105_;
	wire new_net_798;
	wire new_net_1192;
	wire new_net_635;
	wire new_net_817;
	wire new_net_680;
	wire new_net_174;
	wire new_net_192;
	wire new_net_432;
	wire new_net_465;
	wire new_net_1235;
	wire new_net_1247;
	wire new_net_1583;
	wire new_net_1656;
	wire new_net_198;
	wire new_net_456;
	input N1;
	input N101;
	input N105;
	input N109;
	input N113;
	input N117;
	input N121;
	input N125;
	input N129;
	input N13;
	input N130;
	input N131;
	input N132;
	input N133;
	input N134;
	input N135;
	input N136;
	input N137;
	input N17;
	input N21;
	input N25;
	input N29;
	input N33;
	input N37;
	input N41;
	input N45;
	input N49;
	input N5;
	input N53;
	input N57;
	input N61;
	input N65;
	input N69;
	input N73;
	input N77;
	input N81;
	input N85;
	input N89;
	input N9;
	input N93;
	input N97;
	output N724;
	output N725;
	output N726;
	output N727;
	output N728;
	output N729;
	output N730;
	output N731;
	output N732;
	output N733;
	output N734;
	output N735;
	output N736;
	output N737;
	output N738;
	output N739;
	output N740;
	output N741;
	output N742;
	output N743;
	output N744;
	output N745;
	output N746;
	output N747;
	output N748;
	output N749;
	output N750;
	output N751;
	output N752;
	output N753;
	output N754;
	output N755;

	or_ii _362_ (
		.a(new_net_671),
		.b(new_net_447),
		.c(_336_)
	);

	or_bi _363_ (
		.a(new_net_344),
		.b(new_net_215),
		.c(_337_)
	);

	and_bi _364_ (
		.a(new_net_342),
		.b(new_net_212),
		.c(_338_)
	);

	or_bi _365_ (
		.a(_338_),
		.b(_337_),
		.c(_339_)
	);

	or_bi _366_ (
		.a(new_net_94),
		.b(new_net_359),
		.c(_340_)
	);

	and_bi _367_ (
		.a(new_net_98),
		.b(new_net_362),
		.c(_341_)
	);

	or_bi _368_ (
		.a(_341_),
		.b(_340_),
		.c(_342_)
	);

	or_bi _369_ (
		.a(new_net_532),
		.b(new_net_143),
		.c(_343_)
	);

	and_bi _370_ (
		.a(new_net_533),
		.b(new_net_144),
		.c(_344_)
	);

	or_bi _371_ (
		.a(_344_),
		.b(_343_),
		.c(_345_)
	);

	or_bi _372_ (
		.a(new_net_562),
		.b(new_net_252),
		.c(_346_)
	);

	and_bi _373_ (
		.a(new_net_563),
		.b(new_net_253),
		.c(_347_)
	);

	and_bi _374_ (
		.a(_346_),
		.b(_347_),
		.c(_348_)
	);

	or_bb _375_ (
		.a(new_net_209),
		.b(new_net_52),
		.c(_349_)
	);

	and_bb _376_ (
		.a(new_net_207),
		.b(new_net_49),
		.c(_350_)
	);

	and_bi _377_ (
		.a(_349_),
		.b(_350_),
		.c(_351_)
	);

	or_bi _378_ (
		.a(new_net_469),
		.b(new_net_437),
		.c(_352_)
	);

	and_bi _379_ (
		.a(new_net_474),
		.b(new_net_442),
		.c(_353_)
	);

	or_bi _380_ (
		.a(_353_),
		.b(_352_),
		.c(_354_)
	);

	or_bi _381_ (
		.a(new_net_443),
		.b(new_net_505),
		.c(_355_)
	);

	and_bi _382_ (
		.a(new_net_444),
		.b(new_net_506),
		.c(_356_)
	);

	and_bi _383_ (
		.a(_355_),
		.b(_356_),
		.c(_357_)
	);

	or_bb _384_ (
		.a(new_net_230),
		.b(new_net_188),
		.c(_358_)
	);

	and_bb _385_ (
		.a(new_net_234),
		.b(new_net_193),
		.c(_359_)
	);

	and_bi _386_ (
		.a(_358_),
		.b(_359_),
		.c(_360_)
	);

	or_bi _387_ (
		.a(new_net_163),
		.b(new_net_398),
		.c(_361_)
	);

	and_bi _388_ (
		.a(new_net_161),
		.b(new_net_395),
		.c(_000_)
	);

	or_bi _389_ (
		.a(_000_),
		.b(_361_),
		.c(_001_)
	);

	or_bi _390_ (
		.a(new_net_86),
		.b(new_net_0),
		.c(_002_)
	);

	and_bi _391_ (
		.a(new_net_87),
		.b(new_net_1),
		.c(_003_)
	);

	and_bi _392_ (
		.a(_002_),
		.b(_003_),
		.c(_004_)
	);

	or_bb _393_ (
		.a(new_net_90),
		.b(new_net_552),
		.c(_005_)
	);

	and_bb _394_ (
		.a(new_net_93),
		.b(new_net_555),
		.c(_006_)
	);

	and_bi _395_ (
		.a(_005_),
		.b(_006_),
		.c(_007_)
	);

	or_bi _396_ (
		.a(new_net_23),
		.b(new_net_174),
		.c(_008_)
	);

	and_bi _397_ (
		.a(new_net_24),
		.b(new_net_175),
		.c(_009_)
	);

	and_bi _398_ (
		.a(new_net_218),
		.b(new_net_256),
		.c(_010_)
	);

	or_ii _399_ (
		.a(new_net_672),
		.b(new_net_453),
		.c(_011_)
	);

	or_bi _400_ (
		.a(new_net_326),
		.b(new_net_189),
		.c(_012_)
	);

	and_bi _401_ (
		.a(new_net_330),
		.b(new_net_191),
		.c(_013_)
	);

	or_bi _402_ (
		.a(_013_),
		.b(_012_),
		.c(_014_)
	);

	or_bi _403_ (
		.a(new_net_223),
		.b(new_net_54),
		.c(_015_)
	);

	and_bi _404_ (
		.a(new_net_222),
		.b(new_net_50),
		.c(_016_)
	);

	or_bi _405_ (
		.a(_016_),
		.b(_015_),
		.c(_017_)
	);

	or_bi _406_ (
		.a(new_net_417),
		.b(new_net_489),
		.c(_018_)
	);

	and_bi _407_ (
		.a(new_net_418),
		.b(new_net_490),
		.c(_019_)
	);

	or_bi _408_ (
		.a(_019_),
		.b(_018_),
		.c(_020_)
	);

	or_bi _409_ (
		.a(new_net_306),
		.b(new_net_534),
		.c(_021_)
	);

	and_bi _410_ (
		.a(new_net_307),
		.b(new_net_535),
		.c(_022_)
	);

	and_bi _411_ (
		.a(_021_),
		.b(_022_),
		.c(_023_)
	);

	or_bb _412_ (
		.a(new_net_419),
		.b(new_net_360),
		.c(_024_)
	);

	and_bb _413_ (
		.a(new_net_422),
		.b(new_net_363),
		.c(_025_)
	);

	and_bi _414_ (
		.a(_024_),
		.b(_025_),
		.c(_026_)
	);

	or_bi _415_ (
		.a(new_net_319),
		.b(new_net_138),
		.c(_027_)
	);

	and_bi _416_ (
		.a(new_net_316),
		.b(new_net_136),
		.c(_028_)
	);

	or_bi _417_ (
		.a(_028_),
		.b(_027_),
		.c(_029_)
	);

	or_bi _418_ (
		.a(new_net_129),
		.b(new_net_236),
		.c(_030_)
	);

	and_bi _419_ (
		.a(new_net_130),
		.b(new_net_237),
		.c(_031_)
	);

	and_bi _420_ (
		.a(_030_),
		.b(_031_),
		.c(_032_)
	);

	or_bb _421_ (
		.a(new_net_249),
		.b(new_net_216),
		.c(_033_)
	);

	and_bb _422_ (
		.a(new_net_248),
		.b(new_net_213),
		.c(_034_)
	);

	and_bi _423_ (
		.a(_033_),
		.b(_034_),
		.c(_035_)
	);

	or_bi _424_ (
		.a(new_net_178),
		.b(new_net_147),
		.c(_036_)
	);

	and_bi _425_ (
		.a(new_net_181),
		.b(new_net_150),
		.c(_037_)
	);

	or_bi _426_ (
		.a(_037_),
		.b(_036_),
		.c(_038_)
	);

	or_bi _427_ (
		.a(new_net_427),
		.b(new_net_491),
		.c(_039_)
	);

	and_bi _428_ (
		.a(new_net_428),
		.b(new_net_492),
		.c(_040_)
	);

	and_bi _429_ (
		.a(_039_),
		.b(_040_),
		.c(_041_)
	);

	or_bb _430_ (
		.a(new_net_546),
		.b(new_net_322),
		.c(_042_)
	);

	and_bb _431_ (
		.a(new_net_549),
		.b(new_net_323),
		.c(_043_)
	);

	and_bi _432_ (
		.a(_042_),
		.b(_043_),
		.c(_044_)
	);

	and_bi _433_ (
		.a(new_net_39),
		.b(new_net_55),
		.c(_045_)
	);

	and_bi _434_ (
		.a(new_net_56),
		.b(new_net_40),
		.c(_046_)
	);

	or_bb _435_ (
		.a(_046_),
		.b(_045_),
		.c(_047_)
	);

	or_ii _436_ (
		.a(new_net_673),
		.b(new_net_448),
		.c(_048_)
	);

	or_bi _437_ (
		.a(new_net_370),
		.b(new_net_233),
		.c(_049_)
	);

	and_bi _438_ (
		.a(new_net_367),
		.b(new_net_231),
		.c(_050_)
	);

	or_bi _439_ (
		.a(_050_),
		.b(_049_),
		.c(_051_)
	);

	or_bi _440_ (
		.a(new_net_379),
		.b(new_net_206),
		.c(_052_)
	);

	and_bi _441_ (
		.a(new_net_382),
		.b(new_net_211),
		.c(_053_)
	);

	or_bi _442_ (
		.a(_053_),
		.b(_052_),
		.c(_054_)
	);

	or_bi _443_ (
		.a(new_net_254),
		.b(new_net_357),
		.c(_055_)
	);

	and_bi _444_ (
		.a(new_net_255),
		.b(new_net_358),
		.c(_056_)
	);

	or_bi _445_ (
		.a(_056_),
		.b(_055_),
		.c(_057_)
	);

	or_bi _446_ (
		.a(new_net_153),
		.b(new_net_445),
		.c(_058_)
	);

	and_bi _447_ (
		.a(new_net_154),
		.b(new_net_446),
		.c(_059_)
	);

	and_bi _448_ (
		.a(_058_),
		.b(_059_),
		.c(_060_)
	);

	or_bb _449_ (
		.a(new_net_113),
		.b(new_net_97),
		.c(_061_)
	);

	and_bb _450_ (
		.a(new_net_110),
		.b(new_net_96),
		.c(_062_)
	);

	and_bi _451_ (
		.a(_061_),
		.b(_062_),
		.c(_063_)
	);

	or_bi _452_ (
		.a(new_net_59),
		.b(new_net_31),
		.c(_064_)
	);

	and_bi _453_ (
		.a(new_net_63),
		.b(new_net_35),
		.c(_065_)
	);

	or_bi _454_ (
		.a(_065_),
		.b(_064_),
		.c(_066_)
	);

	or_bi _455_ (
		.a(new_net_558),
		.b(new_net_75),
		.c(_067_)
	);

	and_bi _456_ (
		.a(new_net_559),
		.b(new_net_76),
		.c(_068_)
	);

	and_bi _457_ (
		.a(_067_),
		.b(_068_),
		.c(_069_)
	);

	or_bb _458_ (
		.a(new_net_405),
		.b(new_net_341),
		.c(_070_)
	);

	and_bb _459_ (
		.a(new_net_408),
		.b(new_net_345),
		.c(_071_)
	);

	and_bi _460_ (
		.a(_070_),
		.b(_071_),
		.c(_072_)
	);

	or_bi _461_ (
		.a(new_net_352),
		.b(new_net_275),
		.c(_073_)
	);

	and_bi _462_ (
		.a(new_net_350),
		.b(new_net_274),
		.c(_074_)
	);

	or_bi _463_ (
		.a(_074_),
		.b(_073_),
		.c(_075_)
	);

	or_bi _464_ (
		.a(new_net_266),
		.b(new_net_377),
		.c(_076_)
	);

	and_bi _465_ (
		.a(new_net_267),
		.b(new_net_378),
		.c(_077_)
	);

	and_bi _466_ (
		.a(new_net_391),
		.b(new_net_431),
		.c(_078_)
	);

	or_bb _467_ (
		.a(new_net_461),
		.b(new_net_166),
		.c(_079_)
	);

	or_bi _468_ (
		.a(new_net_432),
		.b(new_net_392),
		.c(_080_)
	);

	and_bi _469_ (
		.a(new_net_167),
		.b(new_net_495),
		.c(_081_)
	);

	and_bi _470_ (
		.a(_079_),
		.b(_081_),
		.c(_082_)
	);

	and_bi _471_ (
		.a(new_net_528),
		.b(new_net_501),
		.c(_083_)
	);

	and_bi _472_ (
		.a(new_net_502),
		.b(new_net_529),
		.c(_084_)
	);

	or_bb _473_ (
		.a(_084_),
		.b(_083_),
		.c(_085_)
	);

	and_bi _474_ (
		.a(new_net_118),
		.b(new_net_6),
		.c(_086_)
	);

	inv _475_ (
		.din(new_net_37),
		.dout(_087_)
	);

	or_bi _476_ (
		.a(new_net_257),
		.b(new_net_219),
		.c(_088_)
	);

	and_bi _477_ (
		.a(new_net_151),
		.b(new_net_276),
		.c(_089_)
	);

	and_bi _478_ (
		.a(new_net_273),
		.b(new_net_149),
		.c(_090_)
	);

	or_bb _479_ (
		.a(_090_),
		.b(_089_),
		.c(_091_)
	);

	or_ii _480_ (
		.a(new_net_449),
		.b(new_net_674),
		.c(_092_)
	);

	or_bi _481_ (
		.a(new_net_34),
		.b(new_net_139),
		.c(_093_)
	);

	and_bi _482_ (
		.a(new_net_32),
		.b(new_net_137),
		.c(_094_)
	);

	and_bi _483_ (
		.a(_093_),
		.b(_094_),
		.c(_095_)
	);

	and_bi _484_ (
		.a(new_net_314),
		.b(new_net_196),
		.c(_096_)
	);

	and_bi _485_ (
		.a(new_net_197),
		.b(new_net_315),
		.c(_097_)
	);

	or_bb _486_ (
		.a(_097_),
		.b(_096_),
		.c(_098_)
	);

	or_bb _487_ (
		.a(new_net_411),
		.b(new_net_176),
		.c(_099_)
	);

	and_bb _488_ (
		.a(new_net_412),
		.b(new_net_177),
		.c(_100_)
	);

	and_bi _489_ (
		.a(_099_),
		.b(_100_),
		.c(_101_)
	);

	or_bb _490_ (
		.a(new_net_380),
		.b(new_net_221),
		.c(_102_)
	);

	and_bb _491_ (
		.a(new_net_383),
		.b(new_net_224),
		.c(_103_)
	);

	and_bi _492_ (
		.a(_102_),
		.b(_103_),
		.c(_104_)
	);

	or_bi _493_ (
		.a(new_net_283),
		.b(new_net_243),
		.c(_105_)
	);

	and_bi _494_ (
		.a(new_net_281),
		.b(new_net_242),
		.c(_106_)
	);

	or_bi _495_ (
		.a(_106_),
		.b(_105_),
		.c(_107_)
	);

	or_bi _496_ (
		.a(new_net_536),
		.b(new_net_47),
		.c(_108_)
	);

	and_bi _497_ (
		.a(new_net_537),
		.b(new_net_48),
		.c(_109_)
	);

	and_bi _498_ (
		.a(_108_),
		.b(_109_),
		.c(_110_)
	);

	or_bb _499_ (
		.a(new_net_131),
		.b(new_net_554),
		.c(_111_)
	);

	and_bb _500_ (
		.a(new_net_134),
		.b(new_net_553),
		.c(_112_)
	);

	and_bi _501_ (
		.a(_111_),
		.b(_112_),
		.c(_113_)
	);

	and_bi _502_ (
		.a(new_net_228),
		.b(new_net_487),
		.c(_114_)
	);

	and_bi _503_ (
		.a(new_net_488),
		.b(new_net_229),
		.c(_115_)
	);

	or_bb _504_ (
		.a(_115_),
		.b(_114_),
		.c(_116_)
	);

	and_bi _505_ (
		.a(new_net_182),
		.b(new_net_353),
		.c(_117_)
	);

	and_bi _506_ (
		.a(new_net_351),
		.b(new_net_180),
		.c(_118_)
	);

	or_bb _507_ (
		.a(_118_),
		.b(_117_),
		.c(_119_)
	);

	or_ii _508_ (
		.a(new_net_675),
		.b(new_net_452),
		.c(_120_)
	);

	or_bi _509_ (
		.a(new_net_61),
		.b(new_net_317),
		.c(_121_)
	);

	and_bi _510_ (
		.a(new_net_62),
		.b(new_net_321),
		.c(_122_)
	);

	and_bi _511_ (
		.a(_121_),
		.b(_122_),
		.c(_123_)
	);

	and_bi _512_ (
		.a(new_net_507),
		.b(new_net_455),
		.c(_124_)
	);

	and_bi _513_ (
		.a(new_net_456),
		.b(new_net_508),
		.c(_125_)
	);

	or_bb _514_ (
		.a(_125_),
		.b(_124_),
		.c(_126_)
	);

	or_bb _515_ (
		.a(new_net_564),
		.b(new_net_425),
		.c(_127_)
	);

	and_bb _516_ (
		.a(new_net_565),
		.b(new_net_426),
		.c(_128_)
	);

	and_bi _517_ (
		.a(_127_),
		.b(_128_),
		.c(_129_)
	);

	or_bb _518_ (
		.a(new_net_371),
		.b(new_net_329),
		.c(_130_)
	);

	and_bb _519_ (
		.a(new_net_368),
		.b(new_net_328),
		.c(_131_)
	);

	and_bi _520_ (
		.a(_130_),
		.b(_131_),
		.c(_132_)
	);

	or_bi _521_ (
		.a(new_net_296),
		.b(new_net_260),
		.c(_133_)
	);

	and_bi _522_ (
		.a(new_net_299),
		.b(new_net_264),
		.c(_134_)
	);

	or_bi _523_ (
		.a(_134_),
		.b(_133_),
		.c(_135_)
	);

	or_bi _524_ (
		.a(new_net_145),
		.b(new_net_238),
		.c(_136_)
	);

	and_bi _525_ (
		.a(new_net_146),
		.b(new_net_239),
		.c(_137_)
	);

	and_bi _526_ (
		.a(new_net_278),
		.b(new_net_310),
		.c(_138_)
	);

	or_bb _527_ (
		.a(new_net_347),
		.b(new_net_91),
		.c(_139_)
	);

	or_bi _528_ (
		.a(new_net_311),
		.b(new_net_279),
		.c(_140_)
	);

	and_bi _529_ (
		.a(new_net_92),
		.b(new_net_566),
		.c(_141_)
	);

	and_bi _530_ (
		.a(_139_),
		.b(_141_),
		.c(_142_)
	);

	and_bi _531_ (
		.a(new_net_463),
		.b(new_net_71),
		.c(_143_)
	);

	and_bi _532_ (
		.a(new_net_72),
		.b(new_net_464),
		.c(_144_)
	);

	or_bb _533_ (
		.a(_144_),
		.b(_143_),
		.c(_145_)
	);

	or_bi _534_ (
		.a(new_net_335),
		.b(new_net_518),
		.c(_146_)
	);

	or_bb _535_ (
		.a(new_net_542),
		.b(new_net_100),
		.c(_147_)
	);

	or_bi _536_ (
		.a(new_net_521),
		.b(new_net_336),
		.c(_148_)
	);

	or_bb _537_ (
		.a(new_net_25),
		.b(new_net_101),
		.c(_149_)
	);

	and_bb _538_ (
		.a(new_net_41),
		.b(new_net_550),
		.c(_150_)
	);

	or_ii _539_ (
		.a(new_net_676),
		.b(new_net_450),
		.c(_151_)
	);

	or_bi _540_ (
		.a(new_net_410),
		.b(new_net_250),
		.c(_152_)
	);

	and_bi _541_ (
		.a(new_net_406),
		.b(new_net_247),
		.c(_153_)
	);

	or_bi _542_ (
		.a(_153_),
		.b(_152_),
		.c(_154_)
	);

	or_bi _543_ (
		.a(new_net_111),
		.b(new_net_420),
		.c(_155_)
	);

	and_bi _544_ (
		.a(new_net_114),
		.b(new_net_424),
		.c(_156_)
	);

	or_bi _545_ (
		.a(_156_),
		.b(_155_),
		.c(_157_)
	);

	or_bi _546_ (
		.a(new_net_194),
		.b(new_net_294),
		.c(_158_)
	);

	and_bi _547_ (
		.a(new_net_195),
		.b(new_net_295),
		.c(_159_)
	);

	or_bi _548_ (
		.a(_159_),
		.b(_158_),
		.c(_160_)
	);

	or_bi _549_ (
		.a(new_net_102),
		.b(new_net_389),
		.c(_161_)
	);

	and_bi _550_ (
		.a(new_net_103),
		.b(new_net_390),
		.c(_162_)
	);

	and_bi _551_ (
		.a(_161_),
		.b(_162_),
		.c(_163_)
	);

	or_bb _552_ (
		.a(new_net_348),
		.b(new_net_132),
		.c(_164_)
	);

	and_bi _553_ (
		.a(new_net_133),
		.b(new_net_567),
		.c(_165_)
	);

	and_bi _554_ (
		.a(_164_),
		.b(_165_),
		.c(_166_)
	);

	and_bi _555_ (
		.a(new_net_530),
		.b(new_net_475),
		.c(_167_)
	);

	and_bi _556_ (
		.a(new_net_476),
		.b(new_net_531),
		.c(_168_)
	);

	or_bb _557_ (
		.a(_168_),
		.b(_167_),
		.c(_169_)
	);

	or_bb _558_ (
		.a(new_net_17),
		.b(_150_),
		.c(_170_)
	);

	or_bb _559_ (
		.a(new_net_13),
		.b(new_net_286),
		.c(_171_)
	);

	or_ii _560_ (
		.a(new_net_18),
		.b(new_net_288),
		.c(_172_)
	);

	or_ii _561_ (
		.a(new_net_677),
		.b(new_net_69),
		.c(_173_)
	);

	or_bb _562_ (
		.a(new_net_520),
		.b(new_net_338),
		.c(_174_)
	);

	and_bi _563_ (
		.a(_173_),
		.b(new_net_678),
		.c(_175_)
	);

	and_bi _564_ (
		.a(_170_),
		.b(new_net_679),
		.c(_176_)
	);

	and_bi _565_ (
		.a(new_net_396),
		.b(new_net_261),
		.c(_177_)
	);

	and_bi _566_ (
		.a(new_net_265),
		.b(new_net_399),
		.c(_178_)
	);

	or_bb _567_ (
		.a(_178_),
		.b(_177_),
		.c(_179_)
	);

	or_ii _568_ (
		.a(new_net_680),
		.b(new_net_454),
		.c(_180_)
	);

	or_bi _569_ (
		.a(new_net_241),
		.b(new_net_438),
		.c(_181_)
	);

	and_bi _570_ (
		.a(new_net_244),
		.b(new_net_440),
		.c(_182_)
	);

	and_bi _571_ (
		.a(_181_),
		.b(_182_),
		.c(_183_)
	);

	and_bi _572_ (
		.a(new_net_433),
		.b(new_net_355),
		.c(_184_)
	);

	and_bi _573_ (
		.a(new_net_356),
		.b(new_net_434),
		.c(_185_)
	);

	or_bb _574_ (
		.a(_185_),
		.b(_184_),
		.c(_186_)
	);

	or_bb _575_ (
		.a(new_net_499),
		.b(new_net_302),
		.c(_187_)
	);

	and_bb _576_ (
		.a(new_net_500),
		.b(new_net_303),
		.c(_188_)
	);

	and_bi _577_ (
		.a(_187_),
		.b(_188_),
		.c(_189_)
	);

	or_bb _578_ (
		.a(new_net_168),
		.b(new_net_325),
		.c(_190_)
	);

	and_bb _579_ (
		.a(new_net_169),
		.b(new_net_324),
		.c(_191_)
	);

	and_bi _580_ (
		.a(_190_),
		.b(_191_),
		.c(_192_)
	);

	or_bi _581_ (
		.a(new_net_560),
		.b(new_net_73),
		.c(_193_)
	);

	and_bi _582_ (
		.a(new_net_561),
		.b(new_net_74),
		.c(_194_)
	);

	and_bi _583_ (
		.a(new_net_104),
		.b(new_net_127),
		.c(_195_)
	);

	and_bi _584_ (
		.a(new_net_165),
		.b(new_net_300),
		.c(_196_)
	);

	and_bi _585_ (
		.a(new_net_297),
		.b(new_net_160),
		.c(_197_)
	);

	or_bb _586_ (
		.a(_197_),
		.b(_196_),
		.c(_198_)
	);

	or_ii _587_ (
		.a(new_net_681),
		.b(new_net_451),
		.c(_199_)
	);

	or_bi _588_ (
		.a(new_net_284),
		.b(new_net_472),
		.c(_200_)
	);

	and_bi _589_ (
		.a(new_net_282),
		.b(new_net_470),
		.c(_201_)
	);

	and_bi _590_ (
		.a(_200_),
		.b(_201_),
		.c(_202_)
	);

	and_bi _591_ (
		.a(new_net_393),
		.b(new_net_292),
		.c(_203_)
	);

	and_bi _592_ (
		.a(new_net_293),
		.b(new_net_394),
		.c(_204_)
	);

	or_bb _593_ (
		.a(_204_),
		.b(_203_),
		.c(_205_)
	);

	or_bb _594_ (
		.a(new_net_481),
		.b(new_net_270),
		.c(_206_)
	);

	and_bb _595_ (
		.a(new_net_482),
		.b(new_net_271),
		.c(_207_)
	);

	and_bi _596_ (
		.a(_206_),
		.b(_207_),
		.c(_208_)
	);

	or_bb _597_ (
		.a(new_net_462),
		.b(new_net_548),
		.c(_209_)
	);

	and_bi _598_ (
		.a(new_net_547),
		.b(new_net_496),
		.c(_210_)
	);

	and_bi _599_ (
		.a(_209_),
		.b(_210_),
		.c(_211_)
	);

	or_bi _600_ (
		.a(new_net_526),
		.b(new_net_21),
		.c(_212_)
	);

	and_bi _601_ (
		.a(new_net_527),
		.b(new_net_22),
		.c(_213_)
	);

	or_bi _602_ (
		.a(new_net_67),
		.b(new_net_27),
		.c(_214_)
	);

	or_bb _603_ (
		.a(new_net_88),
		.b(new_net_155),
		.c(_215_)
	);

	or_bb _604_ (
		.a(new_net_125),
		.b(new_net_204),
		.c(_216_)
	);

	or_bb _605_ (
		.a(new_net_141),
		.b(new_net_65),
		.c(_217_)
	);

	or_bb _606_ (
		.a(new_net_184),
		.b(new_net_289),
		.c(_218_)
	);

	and_bi _607_ (
		.a(new_net_361),
		.b(new_net_198),
		.c(_219_)
	);

	and_bi _608_ (
		.a(new_net_199),
		.b(new_net_364),
		.c(_220_)
	);

	and_ii _609_ (
		.a(_220_),
		.b(_219_),
		.c(N726)
	);

	or_bi _610_ (
		.a(new_net_185),
		.b(new_net_337),
		.c(_221_)
	);

	and_bi _611_ (
		.a(new_net_312),
		.b(new_net_135),
		.c(_222_)
	);

	and_bi _612_ (
		.a(new_net_140),
		.b(new_net_313),
		.c(_223_)
	);

	and_ii _613_ (
		.a(_223_),
		.b(_222_),
		.c(N724)
	);

	and_bi _614_ (
		.a(new_net_10),
		.b(new_net_124),
		.c(_224_)
	);

	inv _615_ (
		.din(new_net_403),
		.dout(_225_)
	);

	or_bb _616_ (
		.a(new_net_515),
		.b(new_net_142),
		.c(_226_)
	);

	or_bi _617_ (
		.a(new_net_465),
		.b(new_net_334),
		.c(_227_)
	);

	and_bi _618_ (
		.a(new_net_485),
		.b(new_net_36),
		.c(_228_)
	);

	and_bi _619_ (
		.a(new_net_33),
		.b(new_net_486),
		.c(_229_)
	);

	and_ii _620_ (
		.a(_229_),
		.b(_228_),
		.c(N728)
	);

	or_bi _621_ (
		.a(new_net_186),
		.b(new_net_517),
		.c(_230_)
	);

	and_bi _622_ (
		.a(new_net_538),
		.b(new_net_320),
		.c(_231_)
	);

	and_bi _623_ (
		.a(new_net_318),
		.b(new_net_539),
		.c(_232_)
	);

	and_ii _624_ (
		.a(_232_),
		.b(_231_),
		.c(N725)
	);

	or_bi _625_ (
		.a(new_net_128),
		.b(new_net_105),
		.c(_233_)
	);

	and_bi _626_ (
		.a(new_net_28),
		.b(new_net_68),
		.c(_234_)
	);

	or_bb _627_ (
		.a(new_net_81),
		.b(new_net_57),
		.c(_235_)
	);

	and_bb _628_ (
		.a(new_net_106),
		.b(new_net_126),
		.c(_236_)
	);

	or_bb _629_ (
		.a(new_net_8),
		.b(new_net_119),
		.c(_237_)
	);

	or_bb _630_ (
		.a(new_net_682),
		.b(_236_),
		.c(_238_)
	);

	or_bb _631_ (
		.a(new_net_404),
		.b(new_net_38),
		.c(_239_)
	);

	or_bb _632_ (
		.a(new_net_89),
		.b(new_net_58),
		.c(_240_)
	);

	and_bi _633_ (
		.a(_239_),
		.b(new_net_683),
		.c(_241_)
	);

	and_bi _634_ (
		.a(_238_),
		.b(new_net_684),
		.c(_242_)
	);

	or_bb _635_ (
		.a(new_net_332),
		.b(new_net_70),
		.c(_243_)
	);

	or_bb _636_ (
		.a(new_net_373),
		.b(new_net_26),
		.c(_244_)
	);

	or_bi _637_ (
		.a(new_net_385),
		.b(new_net_7),
		.c(_245_)
	);

	and_bi _638_ (
		.a(new_net_210),
		.b(new_net_429),
		.c(_246_)
	);

	and_bi _639_ (
		.a(new_net_430),
		.b(new_net_208),
		.c(_247_)
	);

	and_ii _640_ (
		.a(_247_),
		.b(_246_),
		.c(new_net_709)
	);

	or_bi _641_ (
		.a(new_net_333),
		.b(new_net_15),
		.c(_248_)
	);

	or_bb _642_ (
		.a(new_net_493),
		.b(new_net_551),
		.c(_249_)
	);

	or_bb _643_ (
		.a(new_net_509),
		.b(new_net_157),
		.c(_250_)
	);

	or_bi _644_ (
		.a(new_net_263),
		.b(new_net_524),
		.c(_251_)
	);

	and_bi _645_ (
		.a(new_net_262),
		.b(new_net_525),
		.c(_252_)
	);

	and_bi _646_ (
		.a(_251_),
		.b(_252_),
		.c(new_net_707)
	);

	or_bb _647_ (
		.a(new_net_494),
		.b(new_net_42),
		.c(_253_)
	);

	or_bb _648_ (
		.a(new_net_2),
		.b(new_net_159),
		.c(_254_)
	);

	and_bi _649_ (
		.a(new_net_29),
		.b(new_net_240),
		.c(_255_)
	);

	and_bi _650_ (
		.a(new_net_245),
		.b(new_net_30),
		.c(_256_)
	);

	and_ii _651_ (
		.a(_256_),
		.b(_255_),
		.c(new_net_715)
	);

	or_bb _652_ (
		.a(new_net_512),
		.b(new_net_84),
		.c(_257_)
	);

	and_bi _653_ (
		.a(new_net_116),
		.b(new_net_298),
		.c(_258_)
	);

	and_bi _654_ (
		.a(new_net_301),
		.b(new_net_117),
		.c(_259_)
	);

	and_ii _655_ (
		.a(_259_),
		.b(_258_),
		.c(new_net_691)
	);

	or_bb _656_ (
		.a(new_net_3),
		.b(new_net_85),
		.c(_260_)
	);

	and_bi _657_ (
		.a(new_net_202),
		.b(new_net_280),
		.c(_261_)
	);

	and_bi _658_ (
		.a(new_net_285),
		.b(new_net_203),
		.c(_262_)
	);

	and_ii _659_ (
		.a(_262_),
		.b(_261_),
		.c(new_net_693)
	);

	or_bi _660_ (
		.a(new_net_511),
		.b(new_net_123),
		.c(_263_)
	);

	and_bi _661_ (
		.a(new_net_327),
		.b(new_net_304),
		.c(_264_)
	);

	and_bi _662_ (
		.a(new_net_305),
		.b(new_net_331),
		.c(_265_)
	);

	and_ii _663_ (
		.a(_265_),
		.b(_264_),
		.c(new_net_687)
	);

	or_bi _664_ (
		.a(new_net_5),
		.b(new_net_122),
		.c(_266_)
	);

	and_bi _665_ (
		.a(new_net_220),
		.b(new_net_401),
		.c(_267_)
	);

	and_bi _666_ (
		.a(new_net_402),
		.b(new_net_225),
		.c(_268_)
	);

	and_ii _667_ (
		.a(_268_),
		.b(_267_),
		.c(new_net_701)
	);

	or_bi _668_ (
		.a(new_net_510),
		.b(new_net_11),
		.c(_269_)
	);

	or_bi _669_ (
		.a(new_net_369),
		.b(new_net_483),
		.c(_270_)
	);

	and_bi _670_ (
		.a(new_net_372),
		.b(new_net_484),
		.c(_271_)
	);

	and_bi _671_ (
		.a(_270_),
		.b(_271_),
		.c(new_net_713)
	);

	or_bi _672_ (
		.a(new_net_4),
		.b(new_net_12),
		.c(_272_)
	);

	or_bi _673_ (
		.a(new_net_381),
		.b(new_net_540),
		.c(_273_)
	);

	and_bi _674_ (
		.a(new_net_384),
		.b(new_net_541),
		.c(_274_)
	);

	and_bi _675_ (
		.a(_273_),
		.b(_274_),
		.c(new_net_711)
	);

	or_bb _676_ (
		.a(new_net_374),
		.b(new_net_543),
		.c(_275_)
	);

	or_bb _677_ (
		.a(new_net_43),
		.b(new_net_158),
		.c(_276_)
	);

	and_bi _678_ (
		.a(new_net_79),
		.b(new_net_400),
		.c(_277_)
	);

	and_bi _679_ (
		.a(new_net_397),
		.b(new_net_80),
		.c(_278_)
	);

	and_ii _680_ (
		.a(_278_),
		.b(_277_),
		.c(new_net_695)
	);

	or_bb _681_ (
		.a(new_net_46),
		.b(new_net_82),
		.c(_279_)
	);

	and_bi _682_ (
		.a(new_net_170),
		.b(new_net_164),
		.c(_280_)
	);

	and_bi _683_ (
		.a(new_net_162),
		.b(new_net_171),
		.c(_281_)
	);

	and_ii _684_ (
		.a(_281_),
		.b(_280_),
		.c(new_net_705)
	);

	and_bi _685_ (
		.a(new_net_120),
		.b(new_net_44),
		.c(_282_)
	);

	and_bi _686_ (
		.a(new_net_258),
		.b(new_net_192),
		.c(_283_)
	);

	and_bi _687_ (
		.a(new_net_190),
		.b(new_net_259),
		.c(_284_)
	);

	or_bb _688_ (
		.a(_284_),
		.b(_283_),
		.c(new_net_697)
	);

	and_bi _689_ (
		.a(new_net_14),
		.b(new_net_187),
		.c(_285_)
	);

	and_bi _690_ (
		.a(new_net_365),
		.b(new_net_423),
		.c(_286_)
	);

	and_bi _691_ (
		.a(new_net_421),
		.b(new_net_366),
		.c(_287_)
	);

	or_bb _692_ (
		.a(_287_),
		.b(_286_),
		.c(N727)
	);

	or_bb _693_ (
		.a(new_net_107),
		.b(new_net_205),
		.c(_288_)
	);

	or_bb _694_ (
		.a(new_net_459),
		.b(new_net_516),
		.c(_289_)
	);

	or_bb _695_ (
		.a(new_net_477),
		.b(new_net_287),
		.c(_290_)
	);

	and_bi _696_ (
		.a(new_net_346),
		.b(new_net_497),
		.c(_291_)
	);

	and_bi _697_ (
		.a(new_net_498),
		.b(new_net_343),
		.c(_292_)
	);

	and_ii _698_ (
		.a(_292_),
		.b(_291_),
		.c(N738)
	);

	or_bi _699_ (
		.a(new_net_45),
		.b(new_net_9),
		.c(_293_)
	);

	and_bi _700_ (
		.a(new_net_235),
		.b(new_net_544),
		.c(_294_)
	);

	and_bi _701_ (
		.a(new_net_545),
		.b(new_net_232),
		.c(_295_)
	);

	and_ii _702_ (
		.a(_295_),
		.b(_294_),
		.c(new_net_699)
	);

	or_bi _703_ (
		.a(new_net_478),
		.b(new_net_16),
		.c(_296_)
	);

	and_bi _704_ (
		.a(new_net_409),
		.b(new_net_226),
		.c(_297_)
	);

	and_bi _705_ (
		.a(new_net_227),
		.b(new_net_407),
		.c(_298_)
	);

	and_ii _706_ (
		.a(_298_),
		.b(_297_),
		.c(N739)
	);

	and_bi _707_ (
		.a(new_net_121),
		.b(new_net_388),
		.c(_299_)
	);

	and_bi _708_ (
		.a(new_net_108),
		.b(new_net_53),
		.c(_300_)
	);

	and_bi _709_ (
		.a(new_net_51),
		.b(new_net_109),
		.c(_301_)
	);

	or_bb _710_ (
		.a(_301_),
		.b(_300_),
		.c(new_net_685)
	);

	or_bb _711_ (
		.a(new_net_387),
		.b(new_net_156),
		.c(_302_)
	);

	and_bi _712_ (
		.a(new_net_200),
		.b(new_net_441),
		.c(_303_)
	);

	and_bi _713_ (
		.a(new_net_439),
		.b(new_net_201),
		.c(_304_)
	);

	and_ii _714_ (
		.a(_304_),
		.b(_303_),
		.c(new_net_689)
	);

	or_bb _715_ (
		.a(new_net_386),
		.b(new_net_83),
		.c(_305_)
	);

	and_bi _716_ (
		.a(new_net_308),
		.b(new_net_473),
		.c(_306_)
	);

	and_bi _717_ (
		.a(new_net_471),
		.b(new_net_309),
		.c(_307_)
	);

	and_ii _718_ (
		.a(_307_),
		.b(_306_),
		.c(new_net_703)
	);

	or_bb _719_ (
		.a(new_net_460),
		.b(new_net_66),
		.c(_308_)
	);

	or_bi _720_ (
		.a(new_net_413),
		.b(new_net_519),
		.c(_309_)
	);

	and_bi _721_ (
		.a(new_net_435),
		.b(new_net_179),
		.c(_310_)
	);

	and_bi _722_ (
		.a(new_net_183),
		.b(new_net_436),
		.c(_311_)
	);

	and_ii _723_ (
		.a(_311_),
		.b(_310_),
		.c(N733)
	);

	or_bi _724_ (
		.a(new_net_468),
		.b(new_net_522),
		.c(_312_)
	);

	and_bi _725_ (
		.a(new_net_503),
		.b(new_net_60),
		.c(_313_)
	);

	and_bi _726_ (
		.a(new_net_64),
		.b(new_net_504),
		.c(_314_)
	);

	and_ii _727_ (
		.a(_314_),
		.b(_313_),
		.c(N729)
	);

	or_bb _728_ (
		.a(new_net_414),
		.b(new_net_290),
		.c(_315_)
	);

	and_bi _729_ (
		.a(new_net_214),
		.b(new_net_556),
		.c(_316_)
	);

	and_bi _730_ (
		.a(new_net_557),
		.b(new_net_217),
		.c(_317_)
	);

	and_ii _731_ (
		.a(_317_),
		.b(_316_),
		.c(N734)
	);

	or_bb _732_ (
		.a(new_net_467),
		.b(new_net_291),
		.c(_318_)
	);

	and_bi _733_ (
		.a(new_net_95),
		.b(new_net_77),
		.c(_319_)
	);

	and_bi _734_ (
		.a(new_net_78),
		.b(new_net_99),
		.c(_320_)
	);

	and_ii _735_ (
		.a(_320_),
		.b(_319_),
		.c(N730)
	);

	or_bi _736_ (
		.a(new_net_416),
		.b(new_net_19),
		.c(_321_)
	);

	and_bi _737_ (
		.a(new_net_172),
		.b(new_net_246),
		.c(_322_)
	);

	and_bi _738_ (
		.a(new_net_251),
		.b(new_net_173),
		.c(_323_)
	);

	and_ii _739_ (
		.a(_323_),
		.b(_322_),
		.c(N735)
	);

	or_bi _740_ (
		.a(new_net_479),
		.b(new_net_339),
		.c(_324_)
	);

	and_bi _741_ (
		.a(new_net_268),
		.b(new_net_272),
		.c(_325_)
	);

	and_bi _742_ (
		.a(new_net_277),
		.b(new_net_269),
		.c(_326_)
	);

	and_ii _743_ (
		.a(_326_),
		.b(_325_),
		.c(N736)
	);

	or_bi _744_ (
		.a(new_net_480),
		.b(new_net_523),
		.c(_327_)
	);

	and_bi _745_ (
		.a(new_net_375),
		.b(new_net_349),
		.c(_328_)
	);

	and_bi _746_ (
		.a(new_net_354),
		.b(new_net_376),
		.c(_329_)
	);

	and_ii _747_ (
		.a(_329_),
		.b(_328_),
		.c(N737)
	);

	and_bi _748_ (
		.a(new_net_20),
		.b(new_net_466),
		.c(_330_)
	);

	and_bi _749_ (
		.a(new_net_457),
		.b(new_net_112),
		.c(_331_)
	);

	and_bi _750_ (
		.a(new_net_115),
		.b(new_net_458),
		.c(_332_)
	);

	or_bb _751_ (
		.a(_332_),
		.b(_331_),
		.c(N731)
	);

	or_bi _752_ (
		.a(new_net_415),
		.b(new_net_340),
		.c(_333_)
	);

	and_bi _753_ (
		.a(new_net_513),
		.b(new_net_148),
		.c(_334_)
	);

	and_bi _754_ (
		.a(new_net_152),
		.b(new_net_514),
		.c(_335_)
	);

	and_ii _755_ (
		.a(_335_),
		.b(_334_),
		.c(N732)
	);

	spl2 new_net_599_v_fanout (
		.a(new_net_599),
		.b(new_net_251),
		.c(new_net_246)
	);

	spl2 _330__v_fanout (
		.a(_330_),
		.b(new_net_458),
		.c(new_net_457)
	);

	spl2 _227__v_fanout (
		.a(_227_),
		.b(new_net_486),
		.c(new_net_485)
	);

	spl2 _321__v_fanout (
		.a(_321_),
		.b(new_net_173),
		.c(new_net_172)
	);

	spl2 _296__v_fanout (
		.a(_296_),
		.b(new_net_227),
		.c(new_net_226)
	);

	spl2 new_net_640_v_fanout (
		.a(new_net_640),
		.b(new_net_140),
		.c(new_net_135)
	);

	spl2 _285__v_fanout (
		.a(_285_),
		.b(new_net_366),
		.c(new_net_365)
	);

	spl2 new_net_628_v_fanout (
		.a(new_net_628),
		.b(new_net_421),
		.c(new_net_423)
	);

	spl2 _290__v_fanout (
		.a(_290_),
		.b(new_net_498),
		.c(new_net_497)
	);

	spl2 _333__v_fanout (
		.a(_333_),
		.b(new_net_514),
		.c(new_net_513)
	);

	spl2 _312__v_fanout (
		.a(_312_),
		.b(new_net_504),
		.c(new_net_503)
	);

	spl2 _324__v_fanout (
		.a(_324_),
		.b(new_net_269),
		.c(new_net_268)
	);

	spl2 new_net_634_v_fanout (
		.a(new_net_634),
		.b(new_net_364),
		.c(new_net_361)
	);

	spl2 new_net_629_v_fanout (
		.a(new_net_629),
		.b(new_net_277),
		.c(new_net_272)
	);

	spl2 new_net_613_v_fanout (
		.a(new_net_613),
		.b(new_net_99),
		.c(new_net_95)
	);

	spl2 _230__v_fanout (
		.a(_230_),
		.b(new_net_539),
		.c(new_net_538)
	);

	spl2 new_net_614_v_fanout (
		.a(new_net_614),
		.b(new_net_217),
		.c(new_net_214)
	);

	spl2 new_net_651_v_fanout (
		.a(new_net_651),
		.b(new_net_354),
		.c(new_net_349)
	);

	spl2 _309__v_fanout (
		.a(_309_),
		.b(new_net_436),
		.c(new_net_435)
	);

	spl2 _218__v_fanout (
		.a(_218_),
		.b(new_net_199),
		.c(new_net_198)
	);

	spl2 new_net_596_v_fanout (
		.a(new_net_596),
		.b(new_net_64),
		.c(new_net_60)
	);

	spl2 new_net_605_v_fanout (
		.a(new_net_605),
		.b(new_net_407),
		.c(new_net_409)
	);

	spl2 _327__v_fanout (
		.a(_327_),
		.b(new_net_376),
		.c(new_net_375)
	);

	spl2 _315__v_fanout (
		.a(_315_),
		.b(new_net_557),
		.c(new_net_556)
	);

	spl2 _221__v_fanout (
		.a(_221_),
		.b(new_net_313),
		.c(new_net_312)
	);

	spl2 _318__v_fanout (
		.a(_318_),
		.b(new_net_78),
		.c(new_net_77)
	);

	spl2 _263__v_fanout (
		.a(_263_),
		.b(new_net_305),
		.c(new_net_304)
	);

	spl2 new_net_618_v_fanout (
		.a(new_net_618),
		.b(new_net_384),
		.c(new_net_381)
	);

	spl2 _254__v_fanout (
		.a(_254_),
		.b(new_net_30),
		.c(new_net_29)
	);

	spl2 new_net_568_v_fanout (
		.a(new_net_568),
		.b(new_net_183),
		.c(new_net_179)
	);

	spl2 new_net_637_v_fanout (
		.a(new_net_637),
		.b(new_net_235),
		.c(new_net_232)
	);

	spl2 new_net_648_v_fanout (
		.a(new_net_648),
		.b(new_net_439),
		.c(new_net_441)
	);

	spl2 _279__v_fanout (
		.a(_279_),
		.b(new_net_171),
		.c(new_net_170)
	);

	spl2 _257__v_fanout (
		.a(_257_),
		.b(new_net_117),
		.c(new_net_116)
	);

	spl2 _260__v_fanout (
		.a(_260_),
		.b(new_net_203),
		.c(new_net_202)
	);

	spl2 new_net_645_v_fanout (
		.a(new_net_645),
		.b(new_net_51),
		.c(new_net_53)
	);

	spl2 _299__v_fanout (
		.a(_299_),
		.b(new_net_109),
		.c(new_net_108)
	);

	spl2 new_net_571_v_fanout (
		.a(new_net_571),
		.b(new_net_36),
		.c(new_net_33)
	);

	spl2 new_net_592_v_fanout (
		.a(new_net_592),
		.b(new_net_152),
		.c(new_net_148)
	);

	spl2 new_net_588_v_fanout (
		.a(new_net_588),
		.b(new_net_225),
		.c(new_net_220)
	);

	spl2 new_net_623_v_fanout (
		.a(new_net_623),
		.b(new_net_369),
		.c(new_net_372)
	);

	spl2 _293__v_fanout (
		.a(_293_),
		.b(new_net_545),
		.c(new_net_544)
	);

	spl2 _269__v_fanout (
		.a(_269_),
		.b(new_net_484),
		.c(new_net_483)
	);

	spl2 _272__v_fanout (
		.a(_272_),
		.b(new_net_541),
		.c(new_net_540)
	);

	spl2 _266__v_fanout (
		.a(_266_),
		.b(new_net_402),
		.c(new_net_401)
	);

	spl2 new_net_602_v_fanout (
		.a(new_net_602),
		.b(new_net_331),
		.c(new_net_327)
	);

	spl2 _282__v_fanout (
		.a(_282_),
		.b(new_net_259),
		.c(new_net_258)
	);

	spl2 new_net_611_v_fanout (
		.a(new_net_611),
		.b(new_net_263),
		.c(new_net_262)
	);

	spl2 new_net_633_v_fanout (
		.a(new_net_633),
		.b(new_net_162),
		.c(new_net_164)
	);

	spl2 new_net_654_v_fanout (
		.a(new_net_654),
		.b(new_net_400),
		.c(new_net_397)
	);

	spl2 _245__v_fanout (
		.a(_245_),
		.b(new_net_430),
		.c(new_net_429)
	);

	spl2 _302__v_fanout (
		.a(_302_),
		.b(new_net_201),
		.c(new_net_200)
	);

	spl2 new_net_619_v_fanout (
		.a(new_net_619),
		.b(new_net_208),
		.c(new_net_210)
	);

	spl2 new_net_593_v_fanout (
		.a(new_net_593),
		.b(new_net_301),
		.c(new_net_298)
	);

	spl2 new_net_624_v_fanout (
		.a(new_net_624),
		.b(new_net_245),
		.c(new_net_240)
	);

	spl2 _305__v_fanout (
		.a(_305_),
		.b(new_net_309),
		.c(new_net_308)
	);

	spl2 new_net_609_v_fanout (
		.a(new_net_609),
		.b(new_net_190),
		.c(new_net_192)
	);

	spl2 new_net_585_v_fanout (
		.a(new_net_585),
		.b(new_net_346),
		.c(new_net_343)
	);

	spl2 new_net_577_v_fanout (
		.a(new_net_577),
		.b(new_net_115),
		.c(new_net_112)
	);

	spl2 new_net_580_v_fanout (
		.a(new_net_580),
		.b(new_net_320),
		.c(new_net_318)
	);

	spl2 _250__v_fanout (
		.a(_250_),
		.b(new_net_525),
		.c(new_net_524)
	);

	spl2 _276__v_fanout (
		.a(_276_),
		.b(new_net_80),
		.c(new_net_79)
	);

	spl2 new_net_574_v_fanout (
		.a(new_net_574),
		.b(new_net_471),
		.c(new_net_473)
	);

	spl4L _226__v_fanout (
		.a(_226_),
		.b(new_net_467),
		.c(new_net_465),
		.d(new_net_468),
		.e(new_net_466)
	);

	spl4L new_net_665_v_fanout (
		.a(new_net_665),
		.b(new_net_20),
		.c(new_net_16),
		.d(new_net_19),
		.e(new_net_14)
	);

	spl4L _217__v_fanout (
		.a(_217_),
		.b(new_net_186),
		.c(new_net_184),
		.d(new_net_187),
		.e(new_net_185)
	);

	spl2 new_net_584_v_fanout (
		.a(new_net_584),
		.b(new_net_285),
		.c(new_net_280)
	);

	spl4L new_net_666_v_fanout (
		.a(new_net_666),
		.b(new_net_519),
		.c(new_net_517),
		.d(new_net_523),
		.e(new_net_522)
	);

	spl4L _308__v_fanout (
		.a(_308_),
		.b(new_net_414),
		.c(new_net_413),
		.d(new_net_415),
		.e(new_net_416)
	);

	spl4L new_net_668_v_fanout (
		.a(new_net_668),
		.b(new_net_291),
		.c(new_net_287),
		.d(new_net_290),
		.e(new_net_289)
	);

	spl4L _289__v_fanout (
		.a(_289_),
		.b(new_net_478),
		.c(new_net_477),
		.d(new_net_479),
		.e(new_net_480)
	);

	spl4L new_net_661_v_fanout (
		.a(new_net_661),
		.b(new_net_339),
		.c(new_net_334),
		.d(new_net_337),
		.e(new_net_340)
	);

	spl4L _244__v_fanout (
		.a(_244_),
		.b(new_net_388),
		.c(new_net_385),
		.d(new_net_386),
		.e(new_net_387)
	);

	spl4L new_net_667_v_fanout (
		.a(new_net_667),
		.b(new_net_11),
		.c(new_net_7),
		.d(new_net_9),
		.e(new_net_12)
	);

	spl4L new_net_669_v_fanout (
		.a(new_net_669),
		.b(new_net_157),
		.c(new_net_159),
		.d(new_net_158),
		.e(new_net_156)
	);

	spl4L _253__v_fanout (
		.a(_253_),
		.b(new_net_3),
		.c(new_net_2),
		.d(new_net_4),
		.e(new_net_5)
	);

	spl4L _275__v_fanout (
		.a(_275_),
		.b(new_net_45),
		.c(new_net_43),
		.d(new_net_46),
		.e(new_net_44)
	);

	spl4L _249__v_fanout (
		.a(_249_),
		.b(new_net_512),
		.c(new_net_509),
		.d(new_net_510),
		.e(new_net_511)
	);

	spl4L new_net_670_v_fanout (
		.a(new_net_670),
		.b(new_net_85),
		.c(new_net_82),
		.d(new_net_83),
		.e(new_net_84)
	);

	spl4L new_net_662_v_fanout (
		.a(new_net_662),
		.b(new_net_122),
		.c(new_net_120),
		.d(new_net_121),
		.e(new_net_123)
	);

	spl2 _216__v_fanout (
		.a(_216_),
		.b(new_net_142),
		.c(new_net_141)
	);

	spl2 _288__v_fanout (
		.a(_288_),
		.b(new_net_460),
		.c(new_net_459)
	);

	spl2 _243__v_fanout (
		.a(_243_),
		.b(new_net_374),
		.c(new_net_373)
	);

	spl2 _248__v_fanout (
		.a(_248_),
		.b(new_net_494),
		.c(new_net_493)
	);

	spl2 _176__v_fanout (
		.a(_176_),
		.b(new_net_205),
		.c(new_net_204)
	);

	spl2 _242__v_fanout (
		.a(_242_),
		.b(new_net_333),
		.c(new_net_332)
	);

	bfr new_net_717_bfr_before (
		.din(new_net_717),
		.dout(new_net_665)
	);

	bfr new_net_718_bfr_before (
		.din(new_net_718),
		.dout(new_net_717)
	);

	bfr new_net_719_bfr_before (
		.din(new_net_719),
		.dout(new_net_718)
	);

	bfr new_net_720_bfr_before (
		.din(new_net_720),
		.dout(new_net_719)
	);

	spl2 new_net_664_v_fanout (
		.a(new_net_664),
		.b(new_net_720),
		.c(new_net_15)
	);

	bfr new_net_721_bfr_before (
		.din(new_net_721),
		.dout(new_net_664)
	);

	spl2 new_net_663_v_fanout (
		.a(new_net_663),
		.b(new_net_721),
		.c(new_net_17)
	);

	bfr new_net_722_bfr_after (
		.din(_225_),
		.dout(new_net_722)
	);

	bfr new_net_723_bfr_after (
		.din(new_net_722),
		.dout(new_net_723)
	);

	bfr new_net_724_bfr_after (
		.din(new_net_723),
		.dout(new_net_724)
	);

	bfr new_net_725_bfr_after (
		.din(new_net_724),
		.dout(new_net_725)
	);

	bfr new_net_726_bfr_after (
		.din(new_net_725),
		.dout(new_net_726)
	);

	bfr new_net_727_bfr_after (
		.din(new_net_726),
		.dout(new_net_727)
	);

	spl2 _225__v_fanout (
		.a(new_net_727),
		.b(new_net_516),
		.c(new_net_515)
	);

	bfr new_net_728_bfr_after (
		.din(_087_),
		.dout(new_net_728)
	);

	bfr new_net_729_bfr_after (
		.din(new_net_728),
		.dout(new_net_729)
	);

	bfr new_net_730_bfr_after (
		.din(new_net_729),
		.dout(new_net_730)
	);

	bfr new_net_731_bfr_after (
		.din(new_net_730),
		.dout(new_net_731)
	);

	bfr new_net_732_bfr_after (
		.din(new_net_731),
		.dout(new_net_732)
	);

	bfr new_net_733_bfr_after (
		.din(new_net_732),
		.dout(new_net_733)
	);

	spl2 _087__v_fanout (
		.a(new_net_733),
		.b(new_net_66),
		.c(new_net_65)
	);

	bfr new_net_734_bfr_before (
		.din(new_net_734),
		.dout(new_net_42)
	);

	bfr new_net_735_bfr_before (
		.din(new_net_735),
		.dout(new_net_734)
	);

	bfr new_net_736_bfr_before (
		.din(new_net_736),
		.dout(new_net_735)
	);

	bfr new_net_737_bfr_before (
		.din(new_net_737),
		.dout(new_net_736)
	);

	bfr new_net_738_bfr_before (
		.din(new_net_738),
		.dout(new_net_737)
	);

	spl2 _149__v_fanout (
		.a(_149_),
		.b(new_net_738),
		.c(new_net_41)
	);

	bfr new_net_739_bfr_before (
		.din(new_net_739),
		.dout(new_net_551)
	);

	bfr new_net_740_bfr_before (
		.din(new_net_740),
		.dout(new_net_739)
	);

	bfr new_net_741_bfr_before (
		.din(new_net_741),
		.dout(new_net_740)
	);

	bfr new_net_742_bfr_before (
		.din(new_net_742),
		.dout(new_net_741)
	);

	bfr new_net_743_bfr_before (
		.din(new_net_743),
		.dout(new_net_742)
	);

	spl2 _147__v_fanout (
		.a(_147_),
		.b(new_net_743),
		.c(new_net_550)
	);

	bfr new_net_744_bfr_before (
		.din(new_net_744),
		.dout(new_net_107)
	);

	bfr new_net_745_bfr_before (
		.din(new_net_745),
		.dout(new_net_744)
	);

	bfr new_net_746_bfr_before (
		.din(new_net_746),
		.dout(new_net_745)
	);

	bfr new_net_747_bfr_before (
		.din(new_net_747),
		.dout(new_net_746)
	);

	bfr new_net_748_bfr_before (
		.din(new_net_748),
		.dout(new_net_747)
	);

	spl2 _235__v_fanout (
		.a(_235_),
		.b(new_net_748),
		.c(new_net_106)
	);

	bfr new_net_749_bfr_before (
		.din(new_net_749),
		.dout(new_net_125)
	);

	bfr new_net_750_bfr_before (
		.din(new_net_750),
		.dout(new_net_749)
	);

	bfr new_net_751_bfr_before (
		.din(new_net_751),
		.dout(new_net_750)
	);

	bfr new_net_752_bfr_before (
		.din(new_net_752),
		.dout(new_net_751)
	);

	bfr new_net_753_bfr_before (
		.din(new_net_753),
		.dout(new_net_752)
	);

	spl2 _215__v_fanout (
		.a(_215_),
		.b(new_net_126),
		.c(new_net_753)
	);

	bfr new_net_754_bfr_before (
		.din(new_net_754),
		.dout(new_net_26)
	);

	bfr new_net_755_bfr_before (
		.din(new_net_755),
		.dout(new_net_754)
	);

	bfr new_net_756_bfr_before (
		.din(new_net_756),
		.dout(new_net_755)
	);

	bfr new_net_757_bfr_before (
		.din(new_net_757),
		.dout(new_net_756)
	);

	bfr new_net_758_bfr_before (
		.din(new_net_758),
		.dout(new_net_757)
	);

	bfr new_net_759_bfr_before (
		.din(new_net_759),
		.dout(new_net_758)
	);

	bfr new_net_760_bfr_before (
		.din(new_net_760),
		.dout(new_net_759)
	);

	spl2 _148__v_fanout (
		.a(_148_),
		.b(new_net_760),
		.c(new_net_25)
	);

	bfr new_net_761_bfr_before (
		.din(new_net_761),
		.dout(new_net_70)
	);

	bfr new_net_762_bfr_before (
		.din(new_net_762),
		.dout(new_net_761)
	);

	bfr new_net_763_bfr_before (
		.din(new_net_763),
		.dout(new_net_762)
	);

	bfr new_net_764_bfr_before (
		.din(new_net_764),
		.dout(new_net_763)
	);

	bfr new_net_765_bfr_before (
		.din(new_net_765),
		.dout(new_net_764)
	);

	spl2 _171__v_fanout (
		.a(_171_),
		.b(new_net_765),
		.c(new_net_69)
	);

	spl2 _086__v_fanout (
		.a(_086_),
		.b(new_net_38),
		.c(new_net_37)
	);

	bfr new_net_766_bfr_before (
		.din(new_net_766),
		.dout(new_net_543)
	);

	bfr new_net_767_bfr_before (
		.din(new_net_767),
		.dout(new_net_766)
	);

	bfr new_net_768_bfr_before (
		.din(new_net_768),
		.dout(new_net_767)
	);

	bfr new_net_769_bfr_before (
		.din(new_net_769),
		.dout(new_net_768)
	);

	bfr new_net_770_bfr_before (
		.din(new_net_770),
		.dout(new_net_769)
	);

	bfr new_net_771_bfr_before (
		.din(new_net_771),
		.dout(new_net_770)
	);

	bfr new_net_772_bfr_before (
		.din(new_net_772),
		.dout(new_net_771)
	);

	spl2 _146__v_fanout (
		.a(_146_),
		.b(new_net_772),
		.c(new_net_542)
	);

	spl2 _224__v_fanout (
		.a(_224_),
		.b(new_net_404),
		.c(new_net_403)
	);

	bfr new_net_773_bfr_before (
		.din(new_net_773),
		.dout(new_net_670)
	);

	bfr new_net_774_bfr_before (
		.din(new_net_774),
		.dout(new_net_773)
	);

	bfr new_net_775_bfr_before (
		.din(new_net_775),
		.dout(new_net_774)
	);

	bfr new_net_776_bfr_before (
		.din(new_net_776),
		.dout(new_net_775)
	);

	bfr new_net_777_bfr_before (
		.din(new_net_777),
		.dout(new_net_776)
	);

	bfr new_net_778_bfr_before (
		.din(new_net_778),
		.dout(new_net_777)
	);

	bfr new_net_779_bfr_before (
		.din(new_net_779),
		.dout(new_net_778)
	);

	bfr new_net_780_bfr_before (
		.din(new_net_780),
		.dout(new_net_779)
	);

	bfr new_net_781_bfr_before (
		.din(new_net_781),
		.dout(new_net_780)
	);

	spl2 _234__v_fanout (
		.a(_234_),
		.b(new_net_81),
		.c(new_net_781)
	);

	spl2 _214__v_fanout (
		.a(_214_),
		.b(new_net_89),
		.c(new_net_88)
	);

	bfr new_net_782_bfr_after (
		.din(_233_),
		.dout(new_net_782)
	);

	spl2 _233__v_fanout (
		.a(new_net_782),
		.b(new_net_58),
		.c(new_net_57)
	);

	bfr new_net_783_bfr_before (
		.din(new_net_783),
		.dout(new_net_667)
	);

	bfr new_net_784_bfr_before (
		.din(new_net_784),
		.dout(new_net_783)
	);

	bfr new_net_785_bfr_before (
		.din(new_net_785),
		.dout(new_net_784)
	);

	bfr new_net_786_bfr_before (
		.din(new_net_786),
		.dout(new_net_785)
	);

	bfr new_net_787_bfr_before (
		.din(new_net_787),
		.dout(new_net_786)
	);

	bfr new_net_788_bfr_before (
		.din(new_net_788),
		.dout(new_net_787)
	);

	bfr new_net_789_bfr_before (
		.din(new_net_789),
		.dout(new_net_788)
	);

	bfr new_net_790_bfr_before (
		.din(new_net_790),
		.dout(new_net_789)
	);

	bfr new_net_791_bfr_before (
		.din(new_net_791),
		.dout(new_net_790)
	);

	bfr new_net_792_bfr_before (
		.din(new_net_792),
		.dout(new_net_791)
	);

	spl4L _085__v_fanout (
		.a(_085_),
		.b(new_net_10),
		.c(new_net_6),
		.d(new_net_792),
		.e(new_net_8)
	);

	bfr new_net_793_bfr_before (
		.din(new_net_793),
		.dout(new_net_663)
	);

	bfr new_net_794_bfr_before (
		.din(new_net_794),
		.dout(new_net_793)
	);

	bfr new_net_795_bfr_before (
		.din(new_net_795),
		.dout(new_net_794)
	);

	bfr new_net_796_bfr_before (
		.din(new_net_796),
		.dout(new_net_795)
	);

	spl3L _169__v_fanout (
		.a(_169_),
		.b(new_net_18),
		.c(new_net_13),
		.d(new_net_796)
	);

	bfr new_net_797_bfr_before (
		.din(new_net_797),
		.dout(new_net_668)
	);

	bfr new_net_798_bfr_before (
		.din(new_net_798),
		.dout(new_net_797)
	);

	bfr new_net_799_bfr_before (
		.din(new_net_799),
		.dout(new_net_798)
	);

	bfr new_net_800_bfr_before (
		.din(new_net_800),
		.dout(new_net_799)
	);

	bfr new_net_801_bfr_before (
		.din(new_net_801),
		.dout(new_net_800)
	);

	bfr new_net_802_bfr_before (
		.din(new_net_802),
		.dout(new_net_801)
	);

	bfr new_net_803_bfr_before (
		.din(new_net_803),
		.dout(new_net_802)
	);

	bfr new_net_804_bfr_before (
		.din(new_net_804),
		.dout(new_net_803)
	);

	bfr new_net_805_bfr_before (
		.din(new_net_805),
		.dout(new_net_804)
	);

	bfr new_net_806_bfr_before (
		.din(new_net_806),
		.dout(new_net_805)
	);

	bfr new_net_807_bfr_before (
		.din(new_net_807),
		.dout(new_net_806)
	);

	spl3L _010__v_fanout (
		.a(_010_),
		.b(new_net_288),
		.c(new_net_286),
		.d(new_net_807)
	);

	bfr new_net_808_bfr_after (
		.din(_088_),
		.dout(new_net_808)
	);

	bfr new_net_809_bfr_after (
		.din(new_net_808),
		.dout(new_net_809)
	);

	spl2 _088__v_fanout (
		.a(new_net_809),
		.b(new_net_101),
		.c(new_net_100)
	);

	bfr new_net_810_bfr_after (
		.din(_195_),
		.dout(new_net_810)
	);

	bfr new_net_811_bfr_before (
		.din(new_net_811),
		.dout(new_net_669)
	);

	bfr new_net_812_bfr_before (
		.din(new_net_812),
		.dout(new_net_811)
	);

	bfr new_net_813_bfr_before (
		.din(new_net_813),
		.dout(new_net_812)
	);

	bfr new_net_814_bfr_before (
		.din(new_net_814),
		.dout(new_net_813)
	);

	bfr new_net_815_bfr_before (
		.din(new_net_815),
		.dout(new_net_814)
	);

	bfr new_net_816_bfr_before (
		.din(new_net_816),
		.dout(new_net_815)
	);

	bfr new_net_817_bfr_before (
		.din(new_net_817),
		.dout(new_net_816)
	);

	bfr new_net_818_bfr_before (
		.din(new_net_818),
		.dout(new_net_817)
	);

	bfr new_net_819_bfr_before (
		.din(new_net_819),
		.dout(new_net_818)
	);

	spl2 _195__v_fanout (
		.a(new_net_810),
		.b(new_net_819),
		.c(new_net_155)
	);

	bfr new_net_820_bfr_before (
		.din(new_net_820),
		.dout(new_net_666)
	);

	bfr new_net_821_bfr_before (
		.din(new_net_821),
		.dout(new_net_820)
	);

	bfr new_net_822_bfr_before (
		.din(new_net_822),
		.dout(new_net_821)
	);

	bfr new_net_823_bfr_before (
		.din(new_net_823),
		.dout(new_net_822)
	);

	bfr new_net_824_bfr_before (
		.din(new_net_824),
		.dout(new_net_823)
	);

	bfr new_net_825_bfr_before (
		.din(new_net_825),
		.dout(new_net_824)
	);

	bfr new_net_826_bfr_before (
		.din(new_net_826),
		.dout(new_net_825)
	);

	bfr new_net_827_bfr_before (
		.din(new_net_827),
		.dout(new_net_826)
	);

	bfr new_net_828_bfr_before (
		.din(new_net_828),
		.dout(new_net_827)
	);

	bfr new_net_829_bfr_before (
		.din(new_net_829),
		.dout(new_net_828)
	);

	bfr new_net_830_bfr_before (
		.din(new_net_830),
		.dout(new_net_829)
	);

	spl4L _145__v_fanout (
		.a(_145_),
		.b(new_net_520),
		.c(new_net_521),
		.d(new_net_830),
		.e(new_net_518)
	);

	spl2 _212__v_fanout (
		.a(_212_),
		.b(new_net_28),
		.c(new_net_27)
	);

	bfr new_net_831_bfr_after (
		.din(_116_),
		.dout(new_net_831)
	);

	bfr new_net_832_bfr_before (
		.din(new_net_832),
		.dout(new_net_661)
	);

	bfr new_net_833_bfr_before (
		.din(new_net_833),
		.dout(new_net_832)
	);

	bfr new_net_834_bfr_before (
		.din(new_net_834),
		.dout(new_net_833)
	);

	bfr new_net_835_bfr_before (
		.din(new_net_835),
		.dout(new_net_834)
	);

	bfr new_net_836_bfr_before (
		.din(new_net_836),
		.dout(new_net_835)
	);

	bfr new_net_837_bfr_before (
		.din(new_net_837),
		.dout(new_net_836)
	);

	bfr new_net_838_bfr_before (
		.din(new_net_838),
		.dout(new_net_837)
	);

	bfr new_net_839_bfr_before (
		.din(new_net_839),
		.dout(new_net_838)
	);

	bfr new_net_840_bfr_before (
		.din(new_net_840),
		.dout(new_net_839)
	);

	bfr new_net_841_bfr_before (
		.din(new_net_841),
		.dout(new_net_840)
	);

	bfr new_net_842_bfr_before (
		.din(new_net_842),
		.dout(new_net_841)
	);

	spl4L _116__v_fanout (
		.a(new_net_831),
		.b(new_net_336),
		.c(new_net_842),
		.d(new_net_338),
		.e(new_net_335)
	);

	bfr new_net_843_bfr_after (
		.din(_047_),
		.dout(new_net_843)
	);

	bfr new_net_844_bfr_before (
		.din(new_net_844),
		.dout(new_net_662)
	);

	bfr new_net_845_bfr_before (
		.din(new_net_845),
		.dout(new_net_844)
	);

	bfr new_net_846_bfr_before (
		.din(new_net_846),
		.dout(new_net_845)
	);

	bfr new_net_847_bfr_before (
		.din(new_net_847),
		.dout(new_net_846)
	);

	bfr new_net_848_bfr_before (
		.din(new_net_848),
		.dout(new_net_847)
	);

	bfr new_net_849_bfr_before (
		.din(new_net_849),
		.dout(new_net_848)
	);

	bfr new_net_850_bfr_before (
		.din(new_net_850),
		.dout(new_net_849)
	);

	bfr new_net_851_bfr_before (
		.din(new_net_851),
		.dout(new_net_850)
	);

	bfr new_net_852_bfr_before (
		.din(new_net_852),
		.dout(new_net_851)
	);

	bfr new_net_853_bfr_before (
		.din(new_net_853),
		.dout(new_net_852)
	);

	spl4L _047__v_fanout (
		.a(new_net_843),
		.b(new_net_119),
		.c(new_net_118),
		.d(new_net_853),
		.e(new_net_124)
	);

	spl2 _213__v_fanout (
		.a(_213_),
		.b(new_net_68),
		.c(new_net_67)
	);

	spl2 _009__v_fanout (
		.a(_009_),
		.b(new_net_257),
		.c(new_net_256)
	);

	spl2 _193__v_fanout (
		.a(_193_),
		.b(new_net_105),
		.c(new_net_104)
	);

	spl2 _194__v_fanout (
		.a(_194_),
		.b(new_net_128),
		.c(new_net_127)
	);

	spl2 _008__v_fanout (
		.a(_008_),
		.b(new_net_219),
		.c(new_net_218)
	);

	spl2 _082__v_fanout (
		.a(_082_),
		.b(new_net_529),
		.c(new_net_528)
	);

	spl2 _142__v_fanout (
		.a(_142_),
		.b(new_net_464),
		.c(new_net_463)
	);

	spl2 _211__v_fanout (
		.a(_211_),
		.b(new_net_22),
		.c(new_net_21)
	);

	spl2 _166__v_fanout (
		.a(_166_),
		.b(new_net_531),
		.c(new_net_530)
	);

	spl2 _007__v_fanout (
		.a(_007_),
		.b(new_net_175),
		.c(new_net_174)
	);

	bfr new_net_854_bfr_after (
		.din(_129_),
		.dout(new_net_854)
	);

	spl2 _129__v_fanout (
		.a(new_net_854),
		.b(new_net_72),
		.c(new_net_71)
	);

	spl2 _113__v_fanout (
		.a(_113_),
		.b(new_net_229),
		.c(new_net_228)
	);

	bfr new_net_855_bfr_after (
		.din(_208_),
		.dout(new_net_855)
	);

	spl2 _208__v_fanout (
		.a(new_net_855),
		.b(new_net_527),
		.c(new_net_526)
	);

	spl2 _348__v_fanout (
		.a(_348_),
		.b(new_net_24),
		.c(new_net_23)
	);

	spl2 _101__v_fanout (
		.a(_101_),
		.b(new_net_488),
		.c(new_net_487)
	);

	spl2 _023__v_fanout (
		.a(_023_),
		.b(new_net_56),
		.c(new_net_55)
	);

	bfr new_net_856_bfr_after (
		.din(_163_),
		.dout(new_net_856)
	);

	spl2 _163__v_fanout (
		.a(new_net_856),
		.b(new_net_476),
		.c(new_net_475)
	);

	spl2 _192__v_fanout (
		.a(_192_),
		.b(new_net_74),
		.c(new_net_73)
	);

	spl2 _189__v_fanout (
		.a(_189_),
		.b(new_net_561),
		.c(new_net_560)
	);

	spl2 _044__v_fanout (
		.a(_044_),
		.b(new_net_40),
		.c(new_net_39)
	);

	bfr new_net_857_bfr_after (
		.din(_060_),
		.dout(new_net_857)
	);

	spl2 _060__v_fanout (
		.a(new_net_857),
		.b(new_net_502),
		.c(new_net_501)
	);

	spl2 new_net_658_v_fanout (
		.a(new_net_658),
		.b(new_net_132),
		.c(new_net_133)
	);

	spl2 _078__v_fanout (
		.a(_078_),
		.b(new_net_462),
		.c(new_net_461)
	);

	spl2 _080__v_fanout (
		.a(_080_),
		.b(new_net_496),
		.c(new_net_495)
	);

	spl2 _138__v_fanout (
		.a(_138_),
		.b(new_net_348),
		.c(new_net_347)
	);

	spl2 new_net_659_v_fanout (
		.a(new_net_659),
		.b(new_net_167),
		.c(new_net_166)
	);

	spl2 _140__v_fanout (
		.a(_140_),
		.b(new_net_567),
		.c(new_net_566)
	);

	spl2 new_net_660_v_fanout (
		.a(new_net_660),
		.b(new_net_547),
		.c(new_net_548)
	);

	spl2 new_net_657_v_fanout (
		.a(new_net_657),
		.b(new_net_92),
		.c(new_net_91)
	);

	spl3L _041__v_fanout (
		.a(_041_),
		.b(new_net_549),
		.c(new_net_546),
		.d(new_net_660)
	);

	spl2 _205__v_fanout (
		.a(_205_),
		.b(new_net_482),
		.c(new_net_481)
	);

	spl3L _110__v_fanout (
		.a(_110_),
		.b(new_net_131),
		.c(new_net_658),
		.d(new_net_134)
	);

	spl3L _004__v_fanout (
		.a(_004_),
		.b(new_net_657),
		.c(new_net_90),
		.d(new_net_93)
	);

	spl4L _357__v_fanout (
		.a(_357_),
		.b(new_net_554),
		.c(new_net_552),
		.d(new_net_553),
		.e(new_net_555)
	);

	spl2 _098__v_fanout (
		.a(_098_),
		.b(new_net_412),
		.c(new_net_411)
	);

	spl2 _020__v_fanout (
		.a(_020_),
		.b(new_net_535),
		.c(new_net_534)
	);

	spl3L _069__v_fanout (
		.a(_069_),
		.b(new_net_169),
		.c(new_net_168),
		.d(new_net_659)
	);

	spl2 _057__v_fanout (
		.a(_057_),
		.b(new_net_446),
		.c(new_net_445)
	);

	spl2 _186__v_fanout (
		.a(_186_),
		.b(new_net_500),
		.c(new_net_499)
	);

	spl2 _126__v_fanout (
		.a(_126_),
		.b(new_net_565),
		.c(new_net_564)
	);

	spl4L _032__v_fanout (
		.a(_032_),
		.b(new_net_325),
		.c(new_net_322),
		.d(new_net_323),
		.e(new_net_324)
	);

	spl2 _160__v_fanout (
		.a(_160_),
		.b(new_net_390),
		.c(new_net_389)
	);

	spl2 _345__v_fanout (
		.a(_345_),
		.b(new_net_253),
		.c(new_net_252)
	);

	spl2 _076__v_fanout (
		.a(_076_),
		.b(new_net_392),
		.c(new_net_391)
	);

	spl2 _137__v_fanout (
		.a(_137_),
		.b(new_net_311),
		.c(new_net_310)
	);

	spl2 _077__v_fanout (
		.a(_077_),
		.b(new_net_432),
		.c(new_net_431)
	);

	spl2 _136__v_fanout (
		.a(_136_),
		.b(new_net_279),
		.c(new_net_278)
	);

	spl2 _001__v_fanout (
		.a(_001_),
		.b(new_net_1),
		.c(new_net_0)
	);

	spl2 _063__v_fanout (
		.a(_063_),
		.b(new_net_559),
		.c(new_net_558)
	);

	spl2 _354__v_fanout (
		.a(_354_),
		.b(new_net_506),
		.c(new_net_505)
	);

	spl2 _072__v_fanout (
		.a(_072_),
		.b(new_net_267),
		.c(new_net_266)
	);

	spl2 _202__v_fanout (
		.a(_202_),
		.b(new_net_394),
		.c(new_net_393)
	);

	spl2 _054__v_fanout (
		.a(_054_),
		.b(new_net_358),
		.c(new_net_357)
	);

	spl2 _038__v_fanout (
		.a(_038_),
		.b(new_net_492),
		.c(new_net_491)
	);

	spl2 _183__v_fanout (
		.a(_183_),
		.b(new_net_434),
		.c(new_net_433)
	);

	spl2 _157__v_fanout (
		.a(_157_),
		.b(new_net_295),
		.c(new_net_294)
	);

	spl2 _014__v_fanout (
		.a(_014_),
		.b(new_net_418),
		.c(new_net_417)
	);

	spl2 _066__v_fanout (
		.a(_066_),
		.b(new_net_76),
		.c(new_net_75)
	);

	spl2 _342__v_fanout (
		.a(_342_),
		.b(new_net_144),
		.c(new_net_143)
	);

	spl2 _351__v_fanout (
		.a(_351_),
		.b(new_net_444),
		.c(new_net_443)
	);

	spl2 _135__v_fanout (
		.a(_135_),
		.b(new_net_239),
		.c(new_net_238)
	);

	spl2 _029__v_fanout (
		.a(_029_),
		.b(new_net_237),
		.c(new_net_236)
	);

	spl2 _339__v_fanout (
		.a(_339_),
		.b(new_net_533),
		.c(new_net_532)
	);

	spl2 _107__v_fanout (
		.a(_107_),
		.b(new_net_48),
		.c(new_net_47)
	);

	spl2 _051__v_fanout (
		.a(_051_),
		.b(new_net_255),
		.c(new_net_254)
	);

	spl2 _132__v_fanout (
		.a(_132_),
		.b(new_net_146),
		.c(new_net_145)
	);

	spl2 _026__v_fanout (
		.a(_026_),
		.b(new_net_130),
		.c(new_net_129)
	);

	bfr new_net_858_bfr_after (
		.din(_119_),
		.dout(new_net_858)
	);

	bfr new_net_859_bfr_after (
		.din(new_net_858),
		.dout(new_net_859)
	);

	bfr new_net_860_bfr_after (
		.din(new_net_859),
		.dout(new_net_860)
	);

	spl2 _119__v_fanout (
		.a(new_net_860),
		.b(new_net_426),
		.c(new_net_425)
	);

	bfr new_net_861_bfr_after (
		.din(_179_),
		.dout(new_net_861)
	);

	bfr new_net_862_bfr_after (
		.din(new_net_861),
		.dout(new_net_862)
	);

	bfr new_net_863_bfr_after (
		.din(new_net_862),
		.dout(new_net_863)
	);

	spl2 _179__v_fanout (
		.a(new_net_863),
		.b(new_net_303),
		.c(new_net_302)
	);

	spl2 _104__v_fanout (
		.a(_104_),
		.b(new_net_537),
		.c(new_net_536)
	);

	spl2 _095__v_fanout (
		.a(_095_),
		.b(new_net_315),
		.c(new_net_314)
	);

	spl2 _017__v_fanout (
		.a(_017_),
		.b(new_net_490),
		.c(new_net_489)
	);

	spl2 _154__v_fanout (
		.a(_154_),
		.b(new_net_195),
		.c(new_net_194)
	);

	spl2 _123__v_fanout (
		.a(_123_),
		.b(new_net_508),
		.c(new_net_507)
	);

	spl2 _035__v_fanout (
		.a(_035_),
		.b(new_net_428),
		.c(new_net_427)
	);

	bfr new_net_864_bfr_after (
		.din(_091_),
		.dout(new_net_864)
	);

	bfr new_net_865_bfr_after (
		.din(new_net_864),
		.dout(new_net_865)
	);

	bfr new_net_866_bfr_after (
		.din(new_net_865),
		.dout(new_net_866)
	);

	spl2 _091__v_fanout (
		.a(new_net_866),
		.b(new_net_177),
		.c(new_net_176)
	);

	bfr new_net_867_bfr_after (
		.din(_198_),
		.dout(new_net_867)
	);

	bfr new_net_868_bfr_after (
		.din(new_net_867),
		.dout(new_net_868)
	);

	bfr new_net_869_bfr_after (
		.din(new_net_868),
		.dout(new_net_869)
	);

	spl2 _198__v_fanout (
		.a(new_net_869),
		.b(new_net_271),
		.c(new_net_270)
	);

	spl2 _360__v_fanout (
		.a(_360_),
		.b(new_net_87),
		.c(new_net_86)
	);

	spl2 _075__v_fanout (
		.a(_075_),
		.b(new_net_378),
		.c(new_net_377)
	);

	bfr new_net_870_bfr_after (
		.din(_199_),
		.dout(new_net_870)
	);

	spl2 _199__v_fanout (
		.a(new_net_870),
		.b(new_net_293),
		.c(new_net_292)
	);

	bfr new_net_871_bfr_after (
		.din(_180_),
		.dout(new_net_871)
	);

	spl2 _180__v_fanout (
		.a(new_net_871),
		.b(new_net_356),
		.c(new_net_355)
	);

	bfr new_net_872_bfr_after (
		.din(_151_),
		.dout(new_net_872)
	);

	bfr new_net_873_bfr_after (
		.din(new_net_872),
		.dout(new_net_873)
	);

	bfr new_net_874_bfr_after (
		.din(new_net_873),
		.dout(new_net_874)
	);

	bfr new_net_875_bfr_after (
		.din(new_net_874),
		.dout(new_net_875)
	);

	spl2 _151__v_fanout (
		.a(new_net_875),
		.b(new_net_103),
		.c(new_net_102)
	);

	bfr new_net_876_bfr_after (
		.din(_120_),
		.dout(new_net_876)
	);

	spl2 _120__v_fanout (
		.a(new_net_876),
		.b(new_net_456),
		.c(new_net_455)
	);

	bfr new_net_877_bfr_after (
		.din(_048_),
		.dout(new_net_877)
	);

	bfr new_net_878_bfr_after (
		.din(new_net_877),
		.dout(new_net_878)
	);

	bfr new_net_879_bfr_after (
		.din(new_net_878),
		.dout(new_net_879)
	);

	bfr new_net_880_bfr_after (
		.din(new_net_879),
		.dout(new_net_880)
	);

	spl2 _048__v_fanout (
		.a(new_net_880),
		.b(new_net_154),
		.c(new_net_153)
	);

	bfr new_net_881_bfr_after (
		.din(_011_),
		.dout(new_net_881)
	);

	bfr new_net_882_bfr_after (
		.din(new_net_881),
		.dout(new_net_882)
	);

	bfr new_net_883_bfr_after (
		.din(new_net_882),
		.dout(new_net_883)
	);

	bfr new_net_884_bfr_after (
		.din(new_net_883),
		.dout(new_net_884)
	);

	spl2 _011__v_fanout (
		.a(new_net_884),
		.b(new_net_307),
		.c(new_net_306)
	);

	bfr new_net_885_bfr_after (
		.din(_092_),
		.dout(new_net_885)
	);

	spl2 _092__v_fanout (
		.a(new_net_885),
		.b(new_net_197),
		.c(new_net_196)
	);

	bfr new_net_886_bfr_after (
		.din(_336_),
		.dout(new_net_886)
	);

	bfr new_net_887_bfr_after (
		.din(new_net_886),
		.dout(new_net_887)
	);

	bfr new_net_888_bfr_after (
		.din(new_net_887),
		.dout(new_net_888)
	);

	bfr new_net_889_bfr_after (
		.din(new_net_888),
		.dout(new_net_889)
	);

	spl2 _336__v_fanout (
		.a(new_net_889),
		.b(new_net_563),
		.c(new_net_562)
	);

	bfr new_net_890_bfr_before (
		.din(new_net_890),
		.dout(new_net_633)
	);

	bfr new_net_891_bfr_before (
		.din(new_net_891),
		.dout(new_net_890)
	);

	bfr new_net_892_bfr_before (
		.din(new_net_892),
		.dout(new_net_891)
	);

	bfr new_net_893_bfr_before (
		.din(new_net_893),
		.dout(new_net_892)
	);

	bfr new_net_894_bfr_before (
		.din(new_net_894),
		.dout(new_net_893)
	);

	bfr new_net_895_bfr_before (
		.din(new_net_895),
		.dout(new_net_894)
	);

	bfr new_net_896_bfr_before (
		.din(new_net_896),
		.dout(new_net_895)
	);

	bfr new_net_897_bfr_before (
		.din(new_net_897),
		.dout(new_net_896)
	);

	bfr new_net_898_bfr_before (
		.din(new_net_898),
		.dout(new_net_897)
	);

	bfr new_net_899_bfr_before (
		.din(new_net_899),
		.dout(new_net_898)
	);

	bfr new_net_900_bfr_before (
		.din(new_net_900),
		.dout(new_net_899)
	);

	bfr new_net_901_bfr_before (
		.din(new_net_901),
		.dout(new_net_900)
	);

	bfr new_net_902_bfr_before (
		.din(new_net_902),
		.dout(new_net_901)
	);

	bfr new_net_903_bfr_before (
		.din(new_net_903),
		.dout(new_net_902)
	);

	bfr new_net_904_bfr_before (
		.din(new_net_904),
		.dout(new_net_903)
	);

	bfr new_net_905_bfr_before (
		.din(new_net_905),
		.dout(new_net_904)
	);

	bfr new_net_906_bfr_before (
		.din(new_net_906),
		.dout(new_net_905)
	);

	bfr new_net_907_bfr_before (
		.din(new_net_907),
		.dout(new_net_906)
	);

	bfr new_net_908_bfr_before (
		.din(new_net_908),
		.dout(new_net_907)
	);

	bfr new_net_909_bfr_before (
		.din(new_net_909),
		.dout(new_net_908)
	);

	bfr new_net_910_bfr_before (
		.din(new_net_910),
		.dout(new_net_909)
	);

	bfr new_net_911_bfr_before (
		.din(new_net_911),
		.dout(new_net_910)
	);

	bfr new_net_912_bfr_before (
		.din(new_net_912),
		.dout(new_net_911)
	);

	bfr new_net_913_bfr_before (
		.din(new_net_913),
		.dout(new_net_912)
	);

	bfr new_net_914_bfr_before (
		.din(new_net_914),
		.dout(new_net_913)
	);

	spl3L new_net_632_v_fanout (
		.a(new_net_632),
		.b(new_net_165),
		.c(new_net_160),
		.d(new_net_914)
	);

	spl2 new_net_572_v_fanout (
		.a(new_net_572),
		.b(new_net_31),
		.c(new_net_35)
	);

	bfr new_net_915_bfr_before (
		.din(new_net_915),
		.dout(new_net_596)
	);

	bfr new_net_916_bfr_before (
		.din(new_net_916),
		.dout(new_net_915)
	);

	bfr new_net_917_bfr_before (
		.din(new_net_917),
		.dout(new_net_916)
	);

	bfr new_net_918_bfr_before (
		.din(new_net_918),
		.dout(new_net_917)
	);

	bfr new_net_919_bfr_before (
		.din(new_net_919),
		.dout(new_net_918)
	);

	bfr new_net_920_bfr_before (
		.din(new_net_920),
		.dout(new_net_919)
	);

	bfr new_net_921_bfr_before (
		.din(new_net_921),
		.dout(new_net_920)
	);

	bfr new_net_922_bfr_before (
		.din(new_net_922),
		.dout(new_net_921)
	);

	bfr new_net_923_bfr_before (
		.din(new_net_923),
		.dout(new_net_922)
	);

	bfr new_net_924_bfr_before (
		.din(new_net_924),
		.dout(new_net_923)
	);

	bfr new_net_925_bfr_before (
		.din(new_net_925),
		.dout(new_net_924)
	);

	bfr new_net_926_bfr_before (
		.din(new_net_926),
		.dout(new_net_925)
	);

	bfr new_net_927_bfr_before (
		.din(new_net_927),
		.dout(new_net_926)
	);

	bfr new_net_928_bfr_before (
		.din(new_net_928),
		.dout(new_net_927)
	);

	bfr new_net_929_bfr_before (
		.din(new_net_929),
		.dout(new_net_928)
	);

	bfr new_net_930_bfr_before (
		.din(new_net_930),
		.dout(new_net_929)
	);

	bfr new_net_931_bfr_before (
		.din(new_net_931),
		.dout(new_net_930)
	);

	bfr new_net_932_bfr_before (
		.din(new_net_932),
		.dout(new_net_931)
	);

	bfr new_net_933_bfr_before (
		.din(new_net_933),
		.dout(new_net_932)
	);

	bfr new_net_934_bfr_before (
		.din(new_net_934),
		.dout(new_net_933)
	);

	bfr new_net_935_bfr_before (
		.din(new_net_935),
		.dout(new_net_934)
	);

	bfr new_net_936_bfr_before (
		.din(new_net_936),
		.dout(new_net_935)
	);

	bfr new_net_937_bfr_before (
		.din(new_net_937),
		.dout(new_net_936)
	);

	bfr new_net_938_bfr_before (
		.din(new_net_938),
		.dout(new_net_937)
	);

	bfr new_net_939_bfr_before (
		.din(new_net_939),
		.dout(new_net_938)
	);

	bfr new_net_940_bfr_before (
		.din(new_net_940),
		.dout(new_net_939)
	);

	spl2 new_net_597_v_fanout (
		.a(new_net_597),
		.b(new_net_61),
		.c(new_net_940)
	);

	spl3L new_net_626_v_fanout (
		.a(new_net_626),
		.b(new_net_243),
		.c(new_net_244),
		.d(new_net_242)
	);

	spl2 new_net_655_v_fanout (
		.a(new_net_655),
		.b(new_net_399),
		.c(new_net_395)
	);

	bfr new_net_941_bfr_before (
		.din(new_net_941),
		.dout(new_net_651)
	);

	bfr new_net_942_bfr_before (
		.din(new_net_942),
		.dout(new_net_941)
	);

	bfr new_net_943_bfr_before (
		.din(new_net_943),
		.dout(new_net_942)
	);

	bfr new_net_944_bfr_before (
		.din(new_net_944),
		.dout(new_net_943)
	);

	bfr new_net_945_bfr_before (
		.din(new_net_945),
		.dout(new_net_944)
	);

	bfr new_net_946_bfr_before (
		.din(new_net_946),
		.dout(new_net_945)
	);

	bfr new_net_947_bfr_before (
		.din(new_net_947),
		.dout(new_net_946)
	);

	bfr new_net_948_bfr_before (
		.din(new_net_948),
		.dout(new_net_947)
	);

	bfr new_net_949_bfr_before (
		.din(new_net_949),
		.dout(new_net_948)
	);

	bfr new_net_950_bfr_before (
		.din(new_net_950),
		.dout(new_net_949)
	);

	bfr new_net_951_bfr_before (
		.din(new_net_951),
		.dout(new_net_950)
	);

	bfr new_net_952_bfr_before (
		.din(new_net_952),
		.dout(new_net_951)
	);

	bfr new_net_953_bfr_before (
		.din(new_net_953),
		.dout(new_net_952)
	);

	bfr new_net_954_bfr_before (
		.din(new_net_954),
		.dout(new_net_953)
	);

	bfr new_net_955_bfr_before (
		.din(new_net_955),
		.dout(new_net_954)
	);

	bfr new_net_956_bfr_before (
		.din(new_net_956),
		.dout(new_net_955)
	);

	bfr new_net_957_bfr_before (
		.din(new_net_957),
		.dout(new_net_956)
	);

	bfr new_net_958_bfr_before (
		.din(new_net_958),
		.dout(new_net_957)
	);

	bfr new_net_959_bfr_before (
		.din(new_net_959),
		.dout(new_net_958)
	);

	bfr new_net_960_bfr_before (
		.din(new_net_960),
		.dout(new_net_959)
	);

	bfr new_net_961_bfr_before (
		.din(new_net_961),
		.dout(new_net_960)
	);

	bfr new_net_962_bfr_before (
		.din(new_net_962),
		.dout(new_net_961)
	);

	bfr new_net_963_bfr_before (
		.din(new_net_963),
		.dout(new_net_962)
	);

	bfr new_net_964_bfr_before (
		.din(new_net_964),
		.dout(new_net_963)
	);

	bfr new_net_965_bfr_before (
		.din(new_net_965),
		.dout(new_net_964)
	);

	bfr new_net_966_bfr_before (
		.din(new_net_966),
		.dout(new_net_965)
	);

	spl3L new_net_653_v_fanout (
		.a(new_net_653),
		.b(new_net_966),
		.c(new_net_352),
		.d(new_net_353)
	);

	bfr new_net_967_bfr_before (
		.din(new_net_967),
		.dout(new_net_568)
	);

	bfr new_net_968_bfr_before (
		.din(new_net_968),
		.dout(new_net_967)
	);

	bfr new_net_969_bfr_before (
		.din(new_net_969),
		.dout(new_net_968)
	);

	bfr new_net_970_bfr_before (
		.din(new_net_970),
		.dout(new_net_969)
	);

	bfr new_net_971_bfr_before (
		.din(new_net_971),
		.dout(new_net_970)
	);

	bfr new_net_972_bfr_before (
		.din(new_net_972),
		.dout(new_net_971)
	);

	bfr new_net_973_bfr_before (
		.din(new_net_973),
		.dout(new_net_972)
	);

	bfr new_net_974_bfr_before (
		.din(new_net_974),
		.dout(new_net_973)
	);

	bfr new_net_975_bfr_before (
		.din(new_net_975),
		.dout(new_net_974)
	);

	bfr new_net_976_bfr_before (
		.din(new_net_976),
		.dout(new_net_975)
	);

	bfr new_net_977_bfr_before (
		.din(new_net_977),
		.dout(new_net_976)
	);

	bfr new_net_978_bfr_before (
		.din(new_net_978),
		.dout(new_net_977)
	);

	bfr new_net_979_bfr_before (
		.din(new_net_979),
		.dout(new_net_978)
	);

	bfr new_net_980_bfr_before (
		.din(new_net_980),
		.dout(new_net_979)
	);

	bfr new_net_981_bfr_before (
		.din(new_net_981),
		.dout(new_net_980)
	);

	bfr new_net_982_bfr_before (
		.din(new_net_982),
		.dout(new_net_981)
	);

	bfr new_net_983_bfr_before (
		.din(new_net_983),
		.dout(new_net_982)
	);

	bfr new_net_984_bfr_before (
		.din(new_net_984),
		.dout(new_net_983)
	);

	bfr new_net_985_bfr_before (
		.din(new_net_985),
		.dout(new_net_984)
	);

	bfr new_net_986_bfr_before (
		.din(new_net_986),
		.dout(new_net_985)
	);

	bfr new_net_987_bfr_before (
		.din(new_net_987),
		.dout(new_net_986)
	);

	bfr new_net_988_bfr_before (
		.din(new_net_988),
		.dout(new_net_987)
	);

	bfr new_net_989_bfr_before (
		.din(new_net_989),
		.dout(new_net_988)
	);

	bfr new_net_990_bfr_before (
		.din(new_net_990),
		.dout(new_net_989)
	);

	bfr new_net_991_bfr_before (
		.din(new_net_991),
		.dout(new_net_990)
	);

	bfr new_net_992_bfr_before (
		.din(new_net_992),
		.dout(new_net_991)
	);

	spl2 new_net_569_v_fanout (
		.a(new_net_569),
		.b(new_net_992),
		.c(new_net_180)
	);

	spl2 new_net_641_v_fanout (
		.a(new_net_641),
		.b(new_net_139),
		.c(new_net_138)
	);

	spl4L new_net_644_v_fanout (
		.a(new_net_644),
		.b(new_net_451),
		.c(new_net_447),
		.d(new_net_448),
		.e(new_net_453)
	);

	bfr new_net_993_bfr_before (
		.din(new_net_993),
		.dout(new_net_599)
	);

	bfr new_net_994_bfr_before (
		.din(new_net_994),
		.dout(new_net_993)
	);

	bfr new_net_995_bfr_before (
		.din(new_net_995),
		.dout(new_net_994)
	);

	bfr new_net_996_bfr_before (
		.din(new_net_996),
		.dout(new_net_995)
	);

	bfr new_net_997_bfr_before (
		.din(new_net_997),
		.dout(new_net_996)
	);

	bfr new_net_998_bfr_before (
		.din(new_net_998),
		.dout(new_net_997)
	);

	bfr new_net_999_bfr_before (
		.din(new_net_999),
		.dout(new_net_998)
	);

	bfr new_net_1000_bfr_before (
		.din(new_net_1000),
		.dout(new_net_999)
	);

	bfr new_net_1001_bfr_before (
		.din(new_net_1001),
		.dout(new_net_1000)
	);

	bfr new_net_1002_bfr_before (
		.din(new_net_1002),
		.dout(new_net_1001)
	);

	bfr new_net_1003_bfr_before (
		.din(new_net_1003),
		.dout(new_net_1002)
	);

	bfr new_net_1004_bfr_before (
		.din(new_net_1004),
		.dout(new_net_1003)
	);

	bfr new_net_1005_bfr_before (
		.din(new_net_1005),
		.dout(new_net_1004)
	);

	bfr new_net_1006_bfr_before (
		.din(new_net_1006),
		.dout(new_net_1005)
	);

	bfr new_net_1007_bfr_before (
		.din(new_net_1007),
		.dout(new_net_1006)
	);

	bfr new_net_1008_bfr_before (
		.din(new_net_1008),
		.dout(new_net_1007)
	);

	bfr new_net_1009_bfr_before (
		.din(new_net_1009),
		.dout(new_net_1008)
	);

	bfr new_net_1010_bfr_before (
		.din(new_net_1010),
		.dout(new_net_1009)
	);

	bfr new_net_1011_bfr_before (
		.din(new_net_1011),
		.dout(new_net_1010)
	);

	bfr new_net_1012_bfr_before (
		.din(new_net_1012),
		.dout(new_net_1011)
	);

	bfr new_net_1013_bfr_before (
		.din(new_net_1013),
		.dout(new_net_1012)
	);

	bfr new_net_1014_bfr_before (
		.din(new_net_1014),
		.dout(new_net_1013)
	);

	bfr new_net_1015_bfr_before (
		.din(new_net_1015),
		.dout(new_net_1014)
	);

	bfr new_net_1016_bfr_before (
		.din(new_net_1016),
		.dout(new_net_1015)
	);

	bfr new_net_1017_bfr_before (
		.din(new_net_1017),
		.dout(new_net_1016)
	);

	bfr new_net_1018_bfr_before (
		.din(new_net_1018),
		.dout(new_net_1017)
	);

	spl2 new_net_600_v_fanout (
		.a(new_net_600),
		.b(new_net_1018),
		.c(new_net_250)
	);

	bfr new_net_1019_bfr_before (
		.din(new_net_1019),
		.dout(new_net_580)
	);

	bfr new_net_1020_bfr_before (
		.din(new_net_1020),
		.dout(new_net_1019)
	);

	bfr new_net_1021_bfr_before (
		.din(new_net_1021),
		.dout(new_net_1020)
	);

	bfr new_net_1022_bfr_before (
		.din(new_net_1022),
		.dout(new_net_1021)
	);

	bfr new_net_1023_bfr_before (
		.din(new_net_1023),
		.dout(new_net_1022)
	);

	bfr new_net_1024_bfr_before (
		.din(new_net_1024),
		.dout(new_net_1023)
	);

	bfr new_net_1025_bfr_before (
		.din(new_net_1025),
		.dout(new_net_1024)
	);

	bfr new_net_1026_bfr_before (
		.din(new_net_1026),
		.dout(new_net_1025)
	);

	bfr new_net_1027_bfr_before (
		.din(new_net_1027),
		.dout(new_net_1026)
	);

	bfr new_net_1028_bfr_before (
		.din(new_net_1028),
		.dout(new_net_1027)
	);

	bfr new_net_1029_bfr_before (
		.din(new_net_1029),
		.dout(new_net_1028)
	);

	bfr new_net_1030_bfr_before (
		.din(new_net_1030),
		.dout(new_net_1029)
	);

	bfr new_net_1031_bfr_before (
		.din(new_net_1031),
		.dout(new_net_1030)
	);

	bfr new_net_1032_bfr_before (
		.din(new_net_1032),
		.dout(new_net_1031)
	);

	bfr new_net_1033_bfr_before (
		.din(new_net_1033),
		.dout(new_net_1032)
	);

	bfr new_net_1034_bfr_before (
		.din(new_net_1034),
		.dout(new_net_1033)
	);

	bfr new_net_1035_bfr_before (
		.din(new_net_1035),
		.dout(new_net_1034)
	);

	bfr new_net_1036_bfr_before (
		.din(new_net_1036),
		.dout(new_net_1035)
	);

	bfr new_net_1037_bfr_before (
		.din(new_net_1037),
		.dout(new_net_1036)
	);

	bfr new_net_1038_bfr_before (
		.din(new_net_1038),
		.dout(new_net_1037)
	);

	bfr new_net_1039_bfr_before (
		.din(new_net_1039),
		.dout(new_net_1038)
	);

	bfr new_net_1040_bfr_before (
		.din(new_net_1040),
		.dout(new_net_1039)
	);

	bfr new_net_1041_bfr_before (
		.din(new_net_1041),
		.dout(new_net_1040)
	);

	bfr new_net_1042_bfr_before (
		.din(new_net_1042),
		.dout(new_net_1041)
	);

	bfr new_net_1043_bfr_before (
		.din(new_net_1043),
		.dout(new_net_1042)
	);

	bfr new_net_1044_bfr_before (
		.din(new_net_1044),
		.dout(new_net_1043)
	);

	spl3L new_net_582_v_fanout (
		.a(new_net_582),
		.b(new_net_321),
		.c(new_net_1044),
		.d(new_net_316)
	);

	spl4L new_net_643_v_fanout (
		.a(new_net_643),
		.b(new_net_450),
		.c(new_net_449),
		.d(new_net_454),
		.e(new_net_452)
	);

	spl3L new_net_598_v_fanout (
		.a(new_net_598),
		.b(new_net_63),
		.c(new_net_59),
		.d(new_net_62)
	);

	bfr new_net_1045_bfr_before (
		.din(new_net_1045),
		.dout(new_net_577)
	);

	bfr new_net_1046_bfr_before (
		.din(new_net_1046),
		.dout(new_net_1045)
	);

	bfr new_net_1047_bfr_before (
		.din(new_net_1047),
		.dout(new_net_1046)
	);

	bfr new_net_1048_bfr_before (
		.din(new_net_1048),
		.dout(new_net_1047)
	);

	bfr new_net_1049_bfr_before (
		.din(new_net_1049),
		.dout(new_net_1048)
	);

	bfr new_net_1050_bfr_before (
		.din(new_net_1050),
		.dout(new_net_1049)
	);

	bfr new_net_1051_bfr_before (
		.din(new_net_1051),
		.dout(new_net_1050)
	);

	bfr new_net_1052_bfr_before (
		.din(new_net_1052),
		.dout(new_net_1051)
	);

	bfr new_net_1053_bfr_before (
		.din(new_net_1053),
		.dout(new_net_1052)
	);

	bfr new_net_1054_bfr_before (
		.din(new_net_1054),
		.dout(new_net_1053)
	);

	bfr new_net_1055_bfr_before (
		.din(new_net_1055),
		.dout(new_net_1054)
	);

	bfr new_net_1056_bfr_before (
		.din(new_net_1056),
		.dout(new_net_1055)
	);

	bfr new_net_1057_bfr_before (
		.din(new_net_1057),
		.dout(new_net_1056)
	);

	bfr new_net_1058_bfr_before (
		.din(new_net_1058),
		.dout(new_net_1057)
	);

	bfr new_net_1059_bfr_before (
		.din(new_net_1059),
		.dout(new_net_1058)
	);

	bfr new_net_1060_bfr_before (
		.din(new_net_1060),
		.dout(new_net_1059)
	);

	bfr new_net_1061_bfr_before (
		.din(new_net_1061),
		.dout(new_net_1060)
	);

	bfr new_net_1062_bfr_before (
		.din(new_net_1062),
		.dout(new_net_1061)
	);

	bfr new_net_1063_bfr_before (
		.din(new_net_1063),
		.dout(new_net_1062)
	);

	bfr new_net_1064_bfr_before (
		.din(new_net_1064),
		.dout(new_net_1063)
	);

	bfr new_net_1065_bfr_before (
		.din(new_net_1065),
		.dout(new_net_1064)
	);

	bfr new_net_1066_bfr_before (
		.din(new_net_1066),
		.dout(new_net_1065)
	);

	bfr new_net_1067_bfr_before (
		.din(new_net_1067),
		.dout(new_net_1066)
	);

	bfr new_net_1068_bfr_before (
		.din(new_net_1068),
		.dout(new_net_1067)
	);

	bfr new_net_1069_bfr_before (
		.din(new_net_1069),
		.dout(new_net_1068)
	);

	bfr new_net_1070_bfr_before (
		.din(new_net_1070),
		.dout(new_net_1069)
	);

	spl3L new_net_579_v_fanout (
		.a(new_net_579),
		.b(new_net_110),
		.c(new_net_1070),
		.d(new_net_111)
	);

	spl2 new_net_603_v_fanout (
		.a(new_net_603),
		.b(new_net_329),
		.c(new_net_328)
	);

	bfr new_net_1071_bfr_before (
		.din(new_net_1071),
		.dout(new_net_634)
	);

	bfr new_net_1072_bfr_before (
		.din(new_net_1072),
		.dout(new_net_1071)
	);

	bfr new_net_1073_bfr_before (
		.din(new_net_1073),
		.dout(new_net_1072)
	);

	bfr new_net_1074_bfr_before (
		.din(new_net_1074),
		.dout(new_net_1073)
	);

	bfr new_net_1075_bfr_before (
		.din(new_net_1075),
		.dout(new_net_1074)
	);

	bfr new_net_1076_bfr_before (
		.din(new_net_1076),
		.dout(new_net_1075)
	);

	bfr new_net_1077_bfr_before (
		.din(new_net_1077),
		.dout(new_net_1076)
	);

	bfr new_net_1078_bfr_before (
		.din(new_net_1078),
		.dout(new_net_1077)
	);

	bfr new_net_1079_bfr_before (
		.din(new_net_1079),
		.dout(new_net_1078)
	);

	bfr new_net_1080_bfr_before (
		.din(new_net_1080),
		.dout(new_net_1079)
	);

	bfr new_net_1081_bfr_before (
		.din(new_net_1081),
		.dout(new_net_1080)
	);

	bfr new_net_1082_bfr_before (
		.din(new_net_1082),
		.dout(new_net_1081)
	);

	bfr new_net_1083_bfr_before (
		.din(new_net_1083),
		.dout(new_net_1082)
	);

	bfr new_net_1084_bfr_before (
		.din(new_net_1084),
		.dout(new_net_1083)
	);

	bfr new_net_1085_bfr_before (
		.din(new_net_1085),
		.dout(new_net_1084)
	);

	bfr new_net_1086_bfr_before (
		.din(new_net_1086),
		.dout(new_net_1085)
	);

	bfr new_net_1087_bfr_before (
		.din(new_net_1087),
		.dout(new_net_1086)
	);

	bfr new_net_1088_bfr_before (
		.din(new_net_1088),
		.dout(new_net_1087)
	);

	bfr new_net_1089_bfr_before (
		.din(new_net_1089),
		.dout(new_net_1088)
	);

	bfr new_net_1090_bfr_before (
		.din(new_net_1090),
		.dout(new_net_1089)
	);

	bfr new_net_1091_bfr_before (
		.din(new_net_1091),
		.dout(new_net_1090)
	);

	bfr new_net_1092_bfr_before (
		.din(new_net_1092),
		.dout(new_net_1091)
	);

	bfr new_net_1093_bfr_before (
		.din(new_net_1093),
		.dout(new_net_1092)
	);

	bfr new_net_1094_bfr_before (
		.din(new_net_1094),
		.dout(new_net_1093)
	);

	bfr new_net_1095_bfr_before (
		.din(new_net_1095),
		.dout(new_net_1094)
	);

	bfr new_net_1096_bfr_before (
		.din(new_net_1096),
		.dout(new_net_1095)
	);

	spl2 new_net_635_v_fanout (
		.a(new_net_635),
		.b(new_net_363),
		.c(new_net_1096)
	);

	spl3L new_net_636_v_fanout (
		.a(new_net_636),
		.b(new_net_362),
		.c(new_net_359),
		.d(new_net_360)
	);

	bfr new_net_1097_bfr_before (
		.din(new_net_1097),
		.dout(new_net_637)
	);

	bfr new_net_1098_bfr_before (
		.din(new_net_1098),
		.dout(new_net_1097)
	);

	bfr new_net_1099_bfr_before (
		.din(new_net_1099),
		.dout(new_net_1098)
	);

	bfr new_net_1100_bfr_before (
		.din(new_net_1100),
		.dout(new_net_1099)
	);

	bfr new_net_1101_bfr_before (
		.din(new_net_1101),
		.dout(new_net_1100)
	);

	bfr new_net_1102_bfr_before (
		.din(new_net_1102),
		.dout(new_net_1101)
	);

	bfr new_net_1103_bfr_before (
		.din(new_net_1103),
		.dout(new_net_1102)
	);

	bfr new_net_1104_bfr_before (
		.din(new_net_1104),
		.dout(new_net_1103)
	);

	bfr new_net_1105_bfr_before (
		.din(new_net_1105),
		.dout(new_net_1104)
	);

	bfr new_net_1106_bfr_before (
		.din(new_net_1106),
		.dout(new_net_1105)
	);

	bfr new_net_1107_bfr_before (
		.din(new_net_1107),
		.dout(new_net_1106)
	);

	bfr new_net_1108_bfr_before (
		.din(new_net_1108),
		.dout(new_net_1107)
	);

	bfr new_net_1109_bfr_before (
		.din(new_net_1109),
		.dout(new_net_1108)
	);

	bfr new_net_1110_bfr_before (
		.din(new_net_1110),
		.dout(new_net_1109)
	);

	bfr new_net_1111_bfr_before (
		.din(new_net_1111),
		.dout(new_net_1110)
	);

	bfr new_net_1112_bfr_before (
		.din(new_net_1112),
		.dout(new_net_1111)
	);

	bfr new_net_1113_bfr_before (
		.din(new_net_1113),
		.dout(new_net_1112)
	);

	bfr new_net_1114_bfr_before (
		.din(new_net_1114),
		.dout(new_net_1113)
	);

	bfr new_net_1115_bfr_before (
		.din(new_net_1115),
		.dout(new_net_1114)
	);

	bfr new_net_1116_bfr_before (
		.din(new_net_1116),
		.dout(new_net_1115)
	);

	bfr new_net_1117_bfr_before (
		.din(new_net_1117),
		.dout(new_net_1116)
	);

	bfr new_net_1118_bfr_before (
		.din(new_net_1118),
		.dout(new_net_1117)
	);

	bfr new_net_1119_bfr_before (
		.din(new_net_1119),
		.dout(new_net_1118)
	);

	bfr new_net_1120_bfr_before (
		.din(new_net_1120),
		.dout(new_net_1119)
	);

	bfr new_net_1121_bfr_before (
		.din(new_net_1121),
		.dout(new_net_1120)
	);

	spl3L new_net_639_v_fanout (
		.a(new_net_639),
		.b(new_net_1121),
		.c(new_net_230),
		.d(new_net_231)
	);

	bfr new_net_1122_bfr_before (
		.din(new_net_1122),
		.dout(new_net_624)
	);

	bfr new_net_1123_bfr_before (
		.din(new_net_1123),
		.dout(new_net_1122)
	);

	bfr new_net_1124_bfr_before (
		.din(new_net_1124),
		.dout(new_net_1123)
	);

	bfr new_net_1125_bfr_before (
		.din(new_net_1125),
		.dout(new_net_1124)
	);

	bfr new_net_1126_bfr_before (
		.din(new_net_1126),
		.dout(new_net_1125)
	);

	bfr new_net_1127_bfr_before (
		.din(new_net_1127),
		.dout(new_net_1126)
	);

	bfr new_net_1128_bfr_before (
		.din(new_net_1128),
		.dout(new_net_1127)
	);

	bfr new_net_1129_bfr_before (
		.din(new_net_1129),
		.dout(new_net_1128)
	);

	bfr new_net_1130_bfr_before (
		.din(new_net_1130),
		.dout(new_net_1129)
	);

	bfr new_net_1131_bfr_before (
		.din(new_net_1131),
		.dout(new_net_1130)
	);

	bfr new_net_1132_bfr_before (
		.din(new_net_1132),
		.dout(new_net_1131)
	);

	bfr new_net_1133_bfr_before (
		.din(new_net_1133),
		.dout(new_net_1132)
	);

	bfr new_net_1134_bfr_before (
		.din(new_net_1134),
		.dout(new_net_1133)
	);

	bfr new_net_1135_bfr_before (
		.din(new_net_1135),
		.dout(new_net_1134)
	);

	bfr new_net_1136_bfr_before (
		.din(new_net_1136),
		.dout(new_net_1135)
	);

	bfr new_net_1137_bfr_before (
		.din(new_net_1137),
		.dout(new_net_1136)
	);

	bfr new_net_1138_bfr_before (
		.din(new_net_1138),
		.dout(new_net_1137)
	);

	bfr new_net_1139_bfr_before (
		.din(new_net_1139),
		.dout(new_net_1138)
	);

	bfr new_net_1140_bfr_before (
		.din(new_net_1140),
		.dout(new_net_1139)
	);

	bfr new_net_1141_bfr_before (
		.din(new_net_1141),
		.dout(new_net_1140)
	);

	bfr new_net_1142_bfr_before (
		.din(new_net_1142),
		.dout(new_net_1141)
	);

	bfr new_net_1143_bfr_before (
		.din(new_net_1143),
		.dout(new_net_1142)
	);

	bfr new_net_1144_bfr_before (
		.din(new_net_1144),
		.dout(new_net_1143)
	);

	bfr new_net_1145_bfr_before (
		.din(new_net_1145),
		.dout(new_net_1144)
	);

	bfr new_net_1146_bfr_before (
		.din(new_net_1146),
		.dout(new_net_1145)
	);

	spl2 new_net_625_v_fanout (
		.a(new_net_625),
		.b(new_net_241),
		.c(new_net_1146)
	);

	bfr new_net_1147_bfr_before (
		.din(new_net_1147),
		.dout(new_net_640)
	);

	bfr new_net_1148_bfr_before (
		.din(new_net_1148),
		.dout(new_net_1147)
	);

	bfr new_net_1149_bfr_before (
		.din(new_net_1149),
		.dout(new_net_1148)
	);

	bfr new_net_1150_bfr_before (
		.din(new_net_1150),
		.dout(new_net_1149)
	);

	bfr new_net_1151_bfr_before (
		.din(new_net_1151),
		.dout(new_net_1150)
	);

	bfr new_net_1152_bfr_before (
		.din(new_net_1152),
		.dout(new_net_1151)
	);

	bfr new_net_1153_bfr_before (
		.din(new_net_1153),
		.dout(new_net_1152)
	);

	bfr new_net_1154_bfr_before (
		.din(new_net_1154),
		.dout(new_net_1153)
	);

	bfr new_net_1155_bfr_before (
		.din(new_net_1155),
		.dout(new_net_1154)
	);

	bfr new_net_1156_bfr_before (
		.din(new_net_1156),
		.dout(new_net_1155)
	);

	bfr new_net_1157_bfr_before (
		.din(new_net_1157),
		.dout(new_net_1156)
	);

	bfr new_net_1158_bfr_before (
		.din(new_net_1158),
		.dout(new_net_1157)
	);

	bfr new_net_1159_bfr_before (
		.din(new_net_1159),
		.dout(new_net_1158)
	);

	bfr new_net_1160_bfr_before (
		.din(new_net_1160),
		.dout(new_net_1159)
	);

	bfr new_net_1161_bfr_before (
		.din(new_net_1161),
		.dout(new_net_1160)
	);

	bfr new_net_1162_bfr_before (
		.din(new_net_1162),
		.dout(new_net_1161)
	);

	bfr new_net_1163_bfr_before (
		.din(new_net_1163),
		.dout(new_net_1162)
	);

	bfr new_net_1164_bfr_before (
		.din(new_net_1164),
		.dout(new_net_1163)
	);

	bfr new_net_1165_bfr_before (
		.din(new_net_1165),
		.dout(new_net_1164)
	);

	bfr new_net_1166_bfr_before (
		.din(new_net_1166),
		.dout(new_net_1165)
	);

	bfr new_net_1167_bfr_before (
		.din(new_net_1167),
		.dout(new_net_1166)
	);

	bfr new_net_1168_bfr_before (
		.din(new_net_1168),
		.dout(new_net_1167)
	);

	bfr new_net_1169_bfr_before (
		.din(new_net_1169),
		.dout(new_net_1168)
	);

	bfr new_net_1170_bfr_before (
		.din(new_net_1170),
		.dout(new_net_1169)
	);

	bfr new_net_1171_bfr_before (
		.din(new_net_1171),
		.dout(new_net_1170)
	);

	bfr new_net_1172_bfr_before (
		.din(new_net_1172),
		.dout(new_net_1171)
	);

	spl3L new_net_642_v_fanout (
		.a(new_net_642),
		.b(new_net_1172),
		.c(new_net_136),
		.d(new_net_137)
	);

	bfr new_net_1173_bfr_before (
		.din(new_net_1173),
		.dout(new_net_588)
	);

	bfr new_net_1174_bfr_before (
		.din(new_net_1174),
		.dout(new_net_1173)
	);

	bfr new_net_1175_bfr_before (
		.din(new_net_1175),
		.dout(new_net_1174)
	);

	bfr new_net_1176_bfr_before (
		.din(new_net_1176),
		.dout(new_net_1175)
	);

	bfr new_net_1177_bfr_before (
		.din(new_net_1177),
		.dout(new_net_1176)
	);

	bfr new_net_1178_bfr_before (
		.din(new_net_1178),
		.dout(new_net_1177)
	);

	bfr new_net_1179_bfr_before (
		.din(new_net_1179),
		.dout(new_net_1178)
	);

	bfr new_net_1180_bfr_before (
		.din(new_net_1180),
		.dout(new_net_1179)
	);

	bfr new_net_1181_bfr_before (
		.din(new_net_1181),
		.dout(new_net_1180)
	);

	bfr new_net_1182_bfr_before (
		.din(new_net_1182),
		.dout(new_net_1181)
	);

	bfr new_net_1183_bfr_before (
		.din(new_net_1183),
		.dout(new_net_1182)
	);

	bfr new_net_1184_bfr_before (
		.din(new_net_1184),
		.dout(new_net_1183)
	);

	bfr new_net_1185_bfr_before (
		.din(new_net_1185),
		.dout(new_net_1184)
	);

	bfr new_net_1186_bfr_before (
		.din(new_net_1186),
		.dout(new_net_1185)
	);

	bfr new_net_1187_bfr_before (
		.din(new_net_1187),
		.dout(new_net_1186)
	);

	bfr new_net_1188_bfr_before (
		.din(new_net_1188),
		.dout(new_net_1187)
	);

	bfr new_net_1189_bfr_before (
		.din(new_net_1189),
		.dout(new_net_1188)
	);

	bfr new_net_1190_bfr_before (
		.din(new_net_1190),
		.dout(new_net_1189)
	);

	bfr new_net_1191_bfr_before (
		.din(new_net_1191),
		.dout(new_net_1190)
	);

	bfr new_net_1192_bfr_before (
		.din(new_net_1192),
		.dout(new_net_1191)
	);

	bfr new_net_1193_bfr_before (
		.din(new_net_1193),
		.dout(new_net_1192)
	);

	bfr new_net_1194_bfr_before (
		.din(new_net_1194),
		.dout(new_net_1193)
	);

	bfr new_net_1195_bfr_before (
		.din(new_net_1195),
		.dout(new_net_1194)
	);

	bfr new_net_1196_bfr_before (
		.din(new_net_1196),
		.dout(new_net_1195)
	);

	bfr new_net_1197_bfr_before (
		.din(new_net_1197),
		.dout(new_net_1196)
	);

	spl2 new_net_589_v_fanout (
		.a(new_net_589),
		.b(new_net_1197),
		.c(new_net_224)
	);

	bfr new_net_1198_bfr_before (
		.din(new_net_1198),
		.dout(new_net_605)
	);

	bfr new_net_1199_bfr_before (
		.din(new_net_1199),
		.dout(new_net_1198)
	);

	bfr new_net_1200_bfr_before (
		.din(new_net_1200),
		.dout(new_net_1199)
	);

	bfr new_net_1201_bfr_before (
		.din(new_net_1201),
		.dout(new_net_1200)
	);

	bfr new_net_1202_bfr_before (
		.din(new_net_1202),
		.dout(new_net_1201)
	);

	bfr new_net_1203_bfr_before (
		.din(new_net_1203),
		.dout(new_net_1202)
	);

	bfr new_net_1204_bfr_before (
		.din(new_net_1204),
		.dout(new_net_1203)
	);

	bfr new_net_1205_bfr_before (
		.din(new_net_1205),
		.dout(new_net_1204)
	);

	bfr new_net_1206_bfr_before (
		.din(new_net_1206),
		.dout(new_net_1205)
	);

	bfr new_net_1207_bfr_before (
		.din(new_net_1207),
		.dout(new_net_1206)
	);

	bfr new_net_1208_bfr_before (
		.din(new_net_1208),
		.dout(new_net_1207)
	);

	bfr new_net_1209_bfr_before (
		.din(new_net_1209),
		.dout(new_net_1208)
	);

	bfr new_net_1210_bfr_before (
		.din(new_net_1210),
		.dout(new_net_1209)
	);

	bfr new_net_1211_bfr_before (
		.din(new_net_1211),
		.dout(new_net_1210)
	);

	bfr new_net_1212_bfr_before (
		.din(new_net_1212),
		.dout(new_net_1211)
	);

	bfr new_net_1213_bfr_before (
		.din(new_net_1213),
		.dout(new_net_1212)
	);

	bfr new_net_1214_bfr_before (
		.din(new_net_1214),
		.dout(new_net_1213)
	);

	bfr new_net_1215_bfr_before (
		.din(new_net_1215),
		.dout(new_net_1214)
	);

	bfr new_net_1216_bfr_before (
		.din(new_net_1216),
		.dout(new_net_1215)
	);

	bfr new_net_1217_bfr_before (
		.din(new_net_1217),
		.dout(new_net_1216)
	);

	bfr new_net_1218_bfr_before (
		.din(new_net_1218),
		.dout(new_net_1217)
	);

	bfr new_net_1219_bfr_before (
		.din(new_net_1219),
		.dout(new_net_1218)
	);

	bfr new_net_1220_bfr_before (
		.din(new_net_1220),
		.dout(new_net_1219)
	);

	bfr new_net_1221_bfr_before (
		.din(new_net_1221),
		.dout(new_net_1220)
	);

	bfr new_net_1222_bfr_before (
		.din(new_net_1222),
		.dout(new_net_1221)
	);

	bfr new_net_1223_bfr_before (
		.din(new_net_1223),
		.dout(new_net_1222)
	);

	spl3L new_net_607_v_fanout (
		.a(new_net_607),
		.b(new_net_405),
		.c(new_net_410),
		.d(new_net_1223)
	);

	bfr new_net_1224_bfr_before (
		.din(new_net_1224),
		.dout(new_net_629)
	);

	bfr new_net_1225_bfr_before (
		.din(new_net_1225),
		.dout(new_net_1224)
	);

	bfr new_net_1226_bfr_before (
		.din(new_net_1226),
		.dout(new_net_1225)
	);

	bfr new_net_1227_bfr_before (
		.din(new_net_1227),
		.dout(new_net_1226)
	);

	bfr new_net_1228_bfr_before (
		.din(new_net_1228),
		.dout(new_net_1227)
	);

	bfr new_net_1229_bfr_before (
		.din(new_net_1229),
		.dout(new_net_1228)
	);

	bfr new_net_1230_bfr_before (
		.din(new_net_1230),
		.dout(new_net_1229)
	);

	bfr new_net_1231_bfr_before (
		.din(new_net_1231),
		.dout(new_net_1230)
	);

	bfr new_net_1232_bfr_before (
		.din(new_net_1232),
		.dout(new_net_1231)
	);

	bfr new_net_1233_bfr_before (
		.din(new_net_1233),
		.dout(new_net_1232)
	);

	bfr new_net_1234_bfr_before (
		.din(new_net_1234),
		.dout(new_net_1233)
	);

	bfr new_net_1235_bfr_before (
		.din(new_net_1235),
		.dout(new_net_1234)
	);

	bfr new_net_1236_bfr_before (
		.din(new_net_1236),
		.dout(new_net_1235)
	);

	bfr new_net_1237_bfr_before (
		.din(new_net_1237),
		.dout(new_net_1236)
	);

	bfr new_net_1238_bfr_before (
		.din(new_net_1238),
		.dout(new_net_1237)
	);

	bfr new_net_1239_bfr_before (
		.din(new_net_1239),
		.dout(new_net_1238)
	);

	bfr new_net_1240_bfr_before (
		.din(new_net_1240),
		.dout(new_net_1239)
	);

	bfr new_net_1241_bfr_before (
		.din(new_net_1241),
		.dout(new_net_1240)
	);

	bfr new_net_1242_bfr_before (
		.din(new_net_1242),
		.dout(new_net_1241)
	);

	bfr new_net_1243_bfr_before (
		.din(new_net_1243),
		.dout(new_net_1242)
	);

	bfr new_net_1244_bfr_before (
		.din(new_net_1244),
		.dout(new_net_1243)
	);

	bfr new_net_1245_bfr_before (
		.din(new_net_1245),
		.dout(new_net_1244)
	);

	bfr new_net_1246_bfr_before (
		.din(new_net_1246),
		.dout(new_net_1245)
	);

	bfr new_net_1247_bfr_before (
		.din(new_net_1247),
		.dout(new_net_1246)
	);

	bfr new_net_1248_bfr_before (
		.din(new_net_1248),
		.dout(new_net_1247)
	);

	bfr new_net_1249_bfr_before (
		.din(new_net_1249),
		.dout(new_net_1248)
	);

	spl3L new_net_631_v_fanout (
		.a(new_net_631),
		.b(new_net_1249),
		.c(new_net_276),
		.d(new_net_273)
	);

	bfr new_net_1250_bfr_before (
		.din(new_net_1250),
		.dout(new_net_628)
	);

	bfr new_net_1251_bfr_before (
		.din(new_net_1251),
		.dout(new_net_1250)
	);

	bfr new_net_1252_bfr_before (
		.din(new_net_1252),
		.dout(new_net_1251)
	);

	bfr new_net_1253_bfr_before (
		.din(new_net_1253),
		.dout(new_net_1252)
	);

	bfr new_net_1254_bfr_before (
		.din(new_net_1254),
		.dout(new_net_1253)
	);

	bfr new_net_1255_bfr_before (
		.din(new_net_1255),
		.dout(new_net_1254)
	);

	bfr new_net_1256_bfr_before (
		.din(new_net_1256),
		.dout(new_net_1255)
	);

	bfr new_net_1257_bfr_before (
		.din(new_net_1257),
		.dout(new_net_1256)
	);

	bfr new_net_1258_bfr_before (
		.din(new_net_1258),
		.dout(new_net_1257)
	);

	bfr new_net_1259_bfr_before (
		.din(new_net_1259),
		.dout(new_net_1258)
	);

	bfr new_net_1260_bfr_before (
		.din(new_net_1260),
		.dout(new_net_1259)
	);

	bfr new_net_1261_bfr_before (
		.din(new_net_1261),
		.dout(new_net_1260)
	);

	bfr new_net_1262_bfr_before (
		.din(new_net_1262),
		.dout(new_net_1261)
	);

	bfr new_net_1263_bfr_before (
		.din(new_net_1263),
		.dout(new_net_1262)
	);

	bfr new_net_1264_bfr_before (
		.din(new_net_1264),
		.dout(new_net_1263)
	);

	bfr new_net_1265_bfr_before (
		.din(new_net_1265),
		.dout(new_net_1264)
	);

	bfr new_net_1266_bfr_before (
		.din(new_net_1266),
		.dout(new_net_1265)
	);

	bfr new_net_1267_bfr_before (
		.din(new_net_1267),
		.dout(new_net_1266)
	);

	bfr new_net_1268_bfr_before (
		.din(new_net_1268),
		.dout(new_net_1267)
	);

	bfr new_net_1269_bfr_before (
		.din(new_net_1269),
		.dout(new_net_1268)
	);

	bfr new_net_1270_bfr_before (
		.din(new_net_1270),
		.dout(new_net_1269)
	);

	bfr new_net_1271_bfr_before (
		.din(new_net_1271),
		.dout(new_net_1270)
	);

	bfr new_net_1272_bfr_before (
		.din(new_net_1272),
		.dout(new_net_1271)
	);

	bfr new_net_1273_bfr_before (
		.din(new_net_1273),
		.dout(new_net_1272)
	);

	bfr new_net_1274_bfr_before (
		.din(new_net_1274),
		.dout(new_net_1273)
	);

	bfr new_net_1275_bfr_before (
		.din(new_net_1275),
		.dout(new_net_1274)
	);

	spl3L new_net_627_v_fanout (
		.a(new_net_627),
		.b(new_net_420),
		.c(new_net_424),
		.d(new_net_1275)
	);

	bfr new_net_1276_bfr_before (
		.din(new_net_1276),
		.dout(new_net_645)
	);

	bfr new_net_1277_bfr_before (
		.din(new_net_1277),
		.dout(new_net_1276)
	);

	bfr new_net_1278_bfr_before (
		.din(new_net_1278),
		.dout(new_net_1277)
	);

	bfr new_net_1279_bfr_before (
		.din(new_net_1279),
		.dout(new_net_1278)
	);

	bfr new_net_1280_bfr_before (
		.din(new_net_1280),
		.dout(new_net_1279)
	);

	bfr new_net_1281_bfr_before (
		.din(new_net_1281),
		.dout(new_net_1280)
	);

	bfr new_net_1282_bfr_before (
		.din(new_net_1282),
		.dout(new_net_1281)
	);

	bfr new_net_1283_bfr_before (
		.din(new_net_1283),
		.dout(new_net_1282)
	);

	bfr new_net_1284_bfr_before (
		.din(new_net_1284),
		.dout(new_net_1283)
	);

	bfr new_net_1285_bfr_before (
		.din(new_net_1285),
		.dout(new_net_1284)
	);

	bfr new_net_1286_bfr_before (
		.din(new_net_1286),
		.dout(new_net_1285)
	);

	bfr new_net_1287_bfr_before (
		.din(new_net_1287),
		.dout(new_net_1286)
	);

	bfr new_net_1288_bfr_before (
		.din(new_net_1288),
		.dout(new_net_1287)
	);

	bfr new_net_1289_bfr_before (
		.din(new_net_1289),
		.dout(new_net_1288)
	);

	bfr new_net_1290_bfr_before (
		.din(new_net_1290),
		.dout(new_net_1289)
	);

	bfr new_net_1291_bfr_before (
		.din(new_net_1291),
		.dout(new_net_1290)
	);

	bfr new_net_1292_bfr_before (
		.din(new_net_1292),
		.dout(new_net_1291)
	);

	bfr new_net_1293_bfr_before (
		.din(new_net_1293),
		.dout(new_net_1292)
	);

	bfr new_net_1294_bfr_before (
		.din(new_net_1294),
		.dout(new_net_1293)
	);

	bfr new_net_1295_bfr_before (
		.din(new_net_1295),
		.dout(new_net_1294)
	);

	bfr new_net_1296_bfr_before (
		.din(new_net_1296),
		.dout(new_net_1295)
	);

	bfr new_net_1297_bfr_before (
		.din(new_net_1297),
		.dout(new_net_1296)
	);

	bfr new_net_1298_bfr_before (
		.din(new_net_1298),
		.dout(new_net_1297)
	);

	bfr new_net_1299_bfr_before (
		.din(new_net_1299),
		.dout(new_net_1298)
	);

	bfr new_net_1300_bfr_before (
		.din(new_net_1300),
		.dout(new_net_1299)
	);

	spl3L new_net_647_v_fanout (
		.a(new_net_647),
		.b(new_net_50),
		.c(new_net_1300),
		.d(new_net_52)
	);

	bfr new_net_1301_bfr_before (
		.din(new_net_1301),
		.dout(new_net_609)
	);

	bfr new_net_1302_bfr_before (
		.din(new_net_1302),
		.dout(new_net_1301)
	);

	bfr new_net_1303_bfr_before (
		.din(new_net_1303),
		.dout(new_net_1302)
	);

	bfr new_net_1304_bfr_before (
		.din(new_net_1304),
		.dout(new_net_1303)
	);

	bfr new_net_1305_bfr_before (
		.din(new_net_1305),
		.dout(new_net_1304)
	);

	bfr new_net_1306_bfr_before (
		.din(new_net_1306),
		.dout(new_net_1305)
	);

	bfr new_net_1307_bfr_before (
		.din(new_net_1307),
		.dout(new_net_1306)
	);

	bfr new_net_1308_bfr_before (
		.din(new_net_1308),
		.dout(new_net_1307)
	);

	bfr new_net_1309_bfr_before (
		.din(new_net_1309),
		.dout(new_net_1308)
	);

	bfr new_net_1310_bfr_before (
		.din(new_net_1310),
		.dout(new_net_1309)
	);

	bfr new_net_1311_bfr_before (
		.din(new_net_1311),
		.dout(new_net_1310)
	);

	bfr new_net_1312_bfr_before (
		.din(new_net_1312),
		.dout(new_net_1311)
	);

	bfr new_net_1313_bfr_before (
		.din(new_net_1313),
		.dout(new_net_1312)
	);

	bfr new_net_1314_bfr_before (
		.din(new_net_1314),
		.dout(new_net_1313)
	);

	bfr new_net_1315_bfr_before (
		.din(new_net_1315),
		.dout(new_net_1314)
	);

	bfr new_net_1316_bfr_before (
		.din(new_net_1316),
		.dout(new_net_1315)
	);

	bfr new_net_1317_bfr_before (
		.din(new_net_1317),
		.dout(new_net_1316)
	);

	bfr new_net_1318_bfr_before (
		.din(new_net_1318),
		.dout(new_net_1317)
	);

	bfr new_net_1319_bfr_before (
		.din(new_net_1319),
		.dout(new_net_1318)
	);

	bfr new_net_1320_bfr_before (
		.din(new_net_1320),
		.dout(new_net_1319)
	);

	bfr new_net_1321_bfr_before (
		.din(new_net_1321),
		.dout(new_net_1320)
	);

	bfr new_net_1322_bfr_before (
		.din(new_net_1322),
		.dout(new_net_1321)
	);

	bfr new_net_1323_bfr_before (
		.din(new_net_1323),
		.dout(new_net_1322)
	);

	bfr new_net_1324_bfr_before (
		.din(new_net_1324),
		.dout(new_net_1323)
	);

	bfr new_net_1325_bfr_before (
		.din(new_net_1325),
		.dout(new_net_1324)
	);

	spl3L new_net_608_v_fanout (
		.a(new_net_608),
		.b(new_net_1325),
		.c(new_net_191),
		.d(new_net_189)
	);

	spl3L new_net_616_v_fanout (
		.a(new_net_616),
		.b(new_net_213),
		.c(new_net_212),
		.d(new_net_216)
	);

	bfr new_net_1326_bfr_before (
		.din(new_net_1326),
		.dout(new_net_593)
	);

	bfr new_net_1327_bfr_before (
		.din(new_net_1327),
		.dout(new_net_1326)
	);

	bfr new_net_1328_bfr_before (
		.din(new_net_1328),
		.dout(new_net_1327)
	);

	bfr new_net_1329_bfr_before (
		.din(new_net_1329),
		.dout(new_net_1328)
	);

	bfr new_net_1330_bfr_before (
		.din(new_net_1330),
		.dout(new_net_1329)
	);

	bfr new_net_1331_bfr_before (
		.din(new_net_1331),
		.dout(new_net_1330)
	);

	bfr new_net_1332_bfr_before (
		.din(new_net_1332),
		.dout(new_net_1331)
	);

	bfr new_net_1333_bfr_before (
		.din(new_net_1333),
		.dout(new_net_1332)
	);

	bfr new_net_1334_bfr_before (
		.din(new_net_1334),
		.dout(new_net_1333)
	);

	bfr new_net_1335_bfr_before (
		.din(new_net_1335),
		.dout(new_net_1334)
	);

	bfr new_net_1336_bfr_before (
		.din(new_net_1336),
		.dout(new_net_1335)
	);

	bfr new_net_1337_bfr_before (
		.din(new_net_1337),
		.dout(new_net_1336)
	);

	bfr new_net_1338_bfr_before (
		.din(new_net_1338),
		.dout(new_net_1337)
	);

	bfr new_net_1339_bfr_before (
		.din(new_net_1339),
		.dout(new_net_1338)
	);

	bfr new_net_1340_bfr_before (
		.din(new_net_1340),
		.dout(new_net_1339)
	);

	bfr new_net_1341_bfr_before (
		.din(new_net_1341),
		.dout(new_net_1340)
	);

	bfr new_net_1342_bfr_before (
		.din(new_net_1342),
		.dout(new_net_1341)
	);

	bfr new_net_1343_bfr_before (
		.din(new_net_1343),
		.dout(new_net_1342)
	);

	bfr new_net_1344_bfr_before (
		.din(new_net_1344),
		.dout(new_net_1343)
	);

	bfr new_net_1345_bfr_before (
		.din(new_net_1345),
		.dout(new_net_1344)
	);

	bfr new_net_1346_bfr_before (
		.din(new_net_1346),
		.dout(new_net_1345)
	);

	bfr new_net_1347_bfr_before (
		.din(new_net_1347),
		.dout(new_net_1346)
	);

	bfr new_net_1348_bfr_before (
		.din(new_net_1348),
		.dout(new_net_1347)
	);

	bfr new_net_1349_bfr_before (
		.din(new_net_1349),
		.dout(new_net_1348)
	);

	bfr new_net_1350_bfr_before (
		.din(new_net_1350),
		.dout(new_net_1349)
	);

	spl3L new_net_595_v_fanout (
		.a(new_net_595),
		.b(new_net_299),
		.c(new_net_1350),
		.d(new_net_297)
	);

	spl2 new_net_578_v_fanout (
		.a(new_net_578),
		.b(new_net_114),
		.c(new_net_113)
	);

	bfr new_net_1351_bfr_before (
		.din(new_net_1351),
		.dout(new_net_614)
	);

	bfr new_net_1352_bfr_before (
		.din(new_net_1352),
		.dout(new_net_1351)
	);

	bfr new_net_1353_bfr_before (
		.din(new_net_1353),
		.dout(new_net_1352)
	);

	bfr new_net_1354_bfr_before (
		.din(new_net_1354),
		.dout(new_net_1353)
	);

	bfr new_net_1355_bfr_before (
		.din(new_net_1355),
		.dout(new_net_1354)
	);

	bfr new_net_1356_bfr_before (
		.din(new_net_1356),
		.dout(new_net_1355)
	);

	bfr new_net_1357_bfr_before (
		.din(new_net_1357),
		.dout(new_net_1356)
	);

	bfr new_net_1358_bfr_before (
		.din(new_net_1358),
		.dout(new_net_1357)
	);

	bfr new_net_1359_bfr_before (
		.din(new_net_1359),
		.dout(new_net_1358)
	);

	bfr new_net_1360_bfr_before (
		.din(new_net_1360),
		.dout(new_net_1359)
	);

	bfr new_net_1361_bfr_before (
		.din(new_net_1361),
		.dout(new_net_1360)
	);

	bfr new_net_1362_bfr_before (
		.din(new_net_1362),
		.dout(new_net_1361)
	);

	bfr new_net_1363_bfr_before (
		.din(new_net_1363),
		.dout(new_net_1362)
	);

	bfr new_net_1364_bfr_before (
		.din(new_net_1364),
		.dout(new_net_1363)
	);

	bfr new_net_1365_bfr_before (
		.din(new_net_1365),
		.dout(new_net_1364)
	);

	bfr new_net_1366_bfr_before (
		.din(new_net_1366),
		.dout(new_net_1365)
	);

	bfr new_net_1367_bfr_before (
		.din(new_net_1367),
		.dout(new_net_1366)
	);

	bfr new_net_1368_bfr_before (
		.din(new_net_1368),
		.dout(new_net_1367)
	);

	bfr new_net_1369_bfr_before (
		.din(new_net_1369),
		.dout(new_net_1368)
	);

	bfr new_net_1370_bfr_before (
		.din(new_net_1370),
		.dout(new_net_1369)
	);

	bfr new_net_1371_bfr_before (
		.din(new_net_1371),
		.dout(new_net_1370)
	);

	bfr new_net_1372_bfr_before (
		.din(new_net_1372),
		.dout(new_net_1371)
	);

	bfr new_net_1373_bfr_before (
		.din(new_net_1373),
		.dout(new_net_1372)
	);

	bfr new_net_1374_bfr_before (
		.din(new_net_1374),
		.dout(new_net_1373)
	);

	bfr new_net_1375_bfr_before (
		.din(new_net_1375),
		.dout(new_net_1374)
	);

	bfr new_net_1376_bfr_before (
		.din(new_net_1376),
		.dout(new_net_1375)
	);

	spl2 new_net_615_v_fanout (
		.a(new_net_615),
		.b(new_net_215),
		.c(new_net_1376)
	);

	bfr new_net_1377_bfr_before (
		.din(new_net_1377),
		.dout(new_net_623)
	);

	bfr new_net_1378_bfr_before (
		.din(new_net_1378),
		.dout(new_net_1377)
	);

	bfr new_net_1379_bfr_before (
		.din(new_net_1379),
		.dout(new_net_1378)
	);

	bfr new_net_1380_bfr_before (
		.din(new_net_1380),
		.dout(new_net_1379)
	);

	bfr new_net_1381_bfr_before (
		.din(new_net_1381),
		.dout(new_net_1380)
	);

	bfr new_net_1382_bfr_before (
		.din(new_net_1382),
		.dout(new_net_1381)
	);

	bfr new_net_1383_bfr_before (
		.din(new_net_1383),
		.dout(new_net_1382)
	);

	bfr new_net_1384_bfr_before (
		.din(new_net_1384),
		.dout(new_net_1383)
	);

	bfr new_net_1385_bfr_before (
		.din(new_net_1385),
		.dout(new_net_1384)
	);

	bfr new_net_1386_bfr_before (
		.din(new_net_1386),
		.dout(new_net_1385)
	);

	bfr new_net_1387_bfr_before (
		.din(new_net_1387),
		.dout(new_net_1386)
	);

	bfr new_net_1388_bfr_before (
		.din(new_net_1388),
		.dout(new_net_1387)
	);

	bfr new_net_1389_bfr_before (
		.din(new_net_1389),
		.dout(new_net_1388)
	);

	bfr new_net_1390_bfr_before (
		.din(new_net_1390),
		.dout(new_net_1389)
	);

	bfr new_net_1391_bfr_before (
		.din(new_net_1391),
		.dout(new_net_1390)
	);

	bfr new_net_1392_bfr_before (
		.din(new_net_1392),
		.dout(new_net_1391)
	);

	bfr new_net_1393_bfr_before (
		.din(new_net_1393),
		.dout(new_net_1392)
	);

	bfr new_net_1394_bfr_before (
		.din(new_net_1394),
		.dout(new_net_1393)
	);

	bfr new_net_1395_bfr_before (
		.din(new_net_1395),
		.dout(new_net_1394)
	);

	bfr new_net_1396_bfr_before (
		.din(new_net_1396),
		.dout(new_net_1395)
	);

	bfr new_net_1397_bfr_before (
		.din(new_net_1397),
		.dout(new_net_1396)
	);

	bfr new_net_1398_bfr_before (
		.din(new_net_1398),
		.dout(new_net_1397)
	);

	bfr new_net_1399_bfr_before (
		.din(new_net_1399),
		.dout(new_net_1398)
	);

	bfr new_net_1400_bfr_before (
		.din(new_net_1400),
		.dout(new_net_1399)
	);

	bfr new_net_1401_bfr_before (
		.din(new_net_1401),
		.dout(new_net_1400)
	);

	spl3L new_net_622_v_fanout (
		.a(new_net_622),
		.b(new_net_1401),
		.c(new_net_368),
		.d(new_net_371)
	);

	bfr new_net_1402_bfr_before (
		.din(new_net_1402),
		.dout(new_net_618)
	);

	bfr new_net_1403_bfr_before (
		.din(new_net_1403),
		.dout(new_net_1402)
	);

	bfr new_net_1404_bfr_before (
		.din(new_net_1404),
		.dout(new_net_1403)
	);

	bfr new_net_1405_bfr_before (
		.din(new_net_1405),
		.dout(new_net_1404)
	);

	bfr new_net_1406_bfr_before (
		.din(new_net_1406),
		.dout(new_net_1405)
	);

	bfr new_net_1407_bfr_before (
		.din(new_net_1407),
		.dout(new_net_1406)
	);

	bfr new_net_1408_bfr_before (
		.din(new_net_1408),
		.dout(new_net_1407)
	);

	bfr new_net_1409_bfr_before (
		.din(new_net_1409),
		.dout(new_net_1408)
	);

	bfr new_net_1410_bfr_before (
		.din(new_net_1410),
		.dout(new_net_1409)
	);

	bfr new_net_1411_bfr_before (
		.din(new_net_1411),
		.dout(new_net_1410)
	);

	bfr new_net_1412_bfr_before (
		.din(new_net_1412),
		.dout(new_net_1411)
	);

	bfr new_net_1413_bfr_before (
		.din(new_net_1413),
		.dout(new_net_1412)
	);

	bfr new_net_1414_bfr_before (
		.din(new_net_1414),
		.dout(new_net_1413)
	);

	bfr new_net_1415_bfr_before (
		.din(new_net_1415),
		.dout(new_net_1414)
	);

	bfr new_net_1416_bfr_before (
		.din(new_net_1416),
		.dout(new_net_1415)
	);

	bfr new_net_1417_bfr_before (
		.din(new_net_1417),
		.dout(new_net_1416)
	);

	bfr new_net_1418_bfr_before (
		.din(new_net_1418),
		.dout(new_net_1417)
	);

	bfr new_net_1419_bfr_before (
		.din(new_net_1419),
		.dout(new_net_1418)
	);

	bfr new_net_1420_bfr_before (
		.din(new_net_1420),
		.dout(new_net_1419)
	);

	bfr new_net_1421_bfr_before (
		.din(new_net_1421),
		.dout(new_net_1420)
	);

	bfr new_net_1422_bfr_before (
		.din(new_net_1422),
		.dout(new_net_1421)
	);

	bfr new_net_1423_bfr_before (
		.din(new_net_1423),
		.dout(new_net_1422)
	);

	bfr new_net_1424_bfr_before (
		.din(new_net_1424),
		.dout(new_net_1423)
	);

	bfr new_net_1425_bfr_before (
		.din(new_net_1425),
		.dout(new_net_1424)
	);

	bfr new_net_1426_bfr_before (
		.din(new_net_1426),
		.dout(new_net_1425)
	);

	spl3L new_net_617_v_fanout (
		.a(new_net_617),
		.b(new_net_383),
		.c(new_net_1426),
		.d(new_net_380)
	);

	bfr new_net_1427_bfr_before (
		.din(new_net_1427),
		.dout(new_net_613)
	);

	bfr new_net_1428_bfr_before (
		.din(new_net_1428),
		.dout(new_net_1427)
	);

	bfr new_net_1429_bfr_before (
		.din(new_net_1429),
		.dout(new_net_1428)
	);

	bfr new_net_1430_bfr_before (
		.din(new_net_1430),
		.dout(new_net_1429)
	);

	bfr new_net_1431_bfr_before (
		.din(new_net_1431),
		.dout(new_net_1430)
	);

	bfr new_net_1432_bfr_before (
		.din(new_net_1432),
		.dout(new_net_1431)
	);

	bfr new_net_1433_bfr_before (
		.din(new_net_1433),
		.dout(new_net_1432)
	);

	bfr new_net_1434_bfr_before (
		.din(new_net_1434),
		.dout(new_net_1433)
	);

	bfr new_net_1435_bfr_before (
		.din(new_net_1435),
		.dout(new_net_1434)
	);

	bfr new_net_1436_bfr_before (
		.din(new_net_1436),
		.dout(new_net_1435)
	);

	bfr new_net_1437_bfr_before (
		.din(new_net_1437),
		.dout(new_net_1436)
	);

	bfr new_net_1438_bfr_before (
		.din(new_net_1438),
		.dout(new_net_1437)
	);

	bfr new_net_1439_bfr_before (
		.din(new_net_1439),
		.dout(new_net_1438)
	);

	bfr new_net_1440_bfr_before (
		.din(new_net_1440),
		.dout(new_net_1439)
	);

	bfr new_net_1441_bfr_before (
		.din(new_net_1441),
		.dout(new_net_1440)
	);

	bfr new_net_1442_bfr_before (
		.din(new_net_1442),
		.dout(new_net_1441)
	);

	bfr new_net_1443_bfr_before (
		.din(new_net_1443),
		.dout(new_net_1442)
	);

	bfr new_net_1444_bfr_before (
		.din(new_net_1444),
		.dout(new_net_1443)
	);

	bfr new_net_1445_bfr_before (
		.din(new_net_1445),
		.dout(new_net_1444)
	);

	bfr new_net_1446_bfr_before (
		.din(new_net_1446),
		.dout(new_net_1445)
	);

	bfr new_net_1447_bfr_before (
		.din(new_net_1447),
		.dout(new_net_1446)
	);

	bfr new_net_1448_bfr_before (
		.din(new_net_1448),
		.dout(new_net_1447)
	);

	bfr new_net_1449_bfr_before (
		.din(new_net_1449),
		.dout(new_net_1448)
	);

	bfr new_net_1450_bfr_before (
		.din(new_net_1450),
		.dout(new_net_1449)
	);

	bfr new_net_1451_bfr_before (
		.din(new_net_1451),
		.dout(new_net_1450)
	);

	bfr new_net_1452_bfr_before (
		.din(new_net_1452),
		.dout(new_net_1451)
	);

	spl3L new_net_612_v_fanout (
		.a(new_net_612),
		.b(new_net_97),
		.c(new_net_96),
		.d(new_net_1452)
	);

	bfr new_net_1453_bfr_before (
		.din(new_net_1453),
		.dout(new_net_571)
	);

	bfr new_net_1454_bfr_before (
		.din(new_net_1454),
		.dout(new_net_1453)
	);

	bfr new_net_1455_bfr_before (
		.din(new_net_1455),
		.dout(new_net_1454)
	);

	bfr new_net_1456_bfr_before (
		.din(new_net_1456),
		.dout(new_net_1455)
	);

	bfr new_net_1457_bfr_before (
		.din(new_net_1457),
		.dout(new_net_1456)
	);

	bfr new_net_1458_bfr_before (
		.din(new_net_1458),
		.dout(new_net_1457)
	);

	bfr new_net_1459_bfr_before (
		.din(new_net_1459),
		.dout(new_net_1458)
	);

	bfr new_net_1460_bfr_before (
		.din(new_net_1460),
		.dout(new_net_1459)
	);

	bfr new_net_1461_bfr_before (
		.din(new_net_1461),
		.dout(new_net_1460)
	);

	bfr new_net_1462_bfr_before (
		.din(new_net_1462),
		.dout(new_net_1461)
	);

	bfr new_net_1463_bfr_before (
		.din(new_net_1463),
		.dout(new_net_1462)
	);

	bfr new_net_1464_bfr_before (
		.din(new_net_1464),
		.dout(new_net_1463)
	);

	bfr new_net_1465_bfr_before (
		.din(new_net_1465),
		.dout(new_net_1464)
	);

	bfr new_net_1466_bfr_before (
		.din(new_net_1466),
		.dout(new_net_1465)
	);

	bfr new_net_1467_bfr_before (
		.din(new_net_1467),
		.dout(new_net_1466)
	);

	bfr new_net_1468_bfr_before (
		.din(new_net_1468),
		.dout(new_net_1467)
	);

	bfr new_net_1469_bfr_before (
		.din(new_net_1469),
		.dout(new_net_1468)
	);

	bfr new_net_1470_bfr_before (
		.din(new_net_1470),
		.dout(new_net_1469)
	);

	bfr new_net_1471_bfr_before (
		.din(new_net_1471),
		.dout(new_net_1470)
	);

	bfr new_net_1472_bfr_before (
		.din(new_net_1472),
		.dout(new_net_1471)
	);

	bfr new_net_1473_bfr_before (
		.din(new_net_1473),
		.dout(new_net_1472)
	);

	bfr new_net_1474_bfr_before (
		.din(new_net_1474),
		.dout(new_net_1473)
	);

	bfr new_net_1475_bfr_before (
		.din(new_net_1475),
		.dout(new_net_1474)
	);

	bfr new_net_1476_bfr_before (
		.din(new_net_1476),
		.dout(new_net_1475)
	);

	bfr new_net_1477_bfr_before (
		.din(new_net_1477),
		.dout(new_net_1476)
	);

	bfr new_net_1478_bfr_before (
		.din(new_net_1478),
		.dout(new_net_1477)
	);

	spl3L new_net_573_v_fanout (
		.a(new_net_573),
		.b(new_net_34),
		.c(new_net_1478),
		.d(new_net_32)
	);

	spl2 new_net_646_v_fanout (
		.a(new_net_646),
		.b(new_net_54),
		.c(new_net_49)
	);

	spl3L new_net_576_v_fanout (
		.a(new_net_576),
		.b(new_net_470),
		.c(new_net_469),
		.d(new_net_472)
	);

	bfr new_net_1479_bfr_before (
		.din(new_net_1479),
		.dout(new_net_574)
	);

	bfr new_net_1480_bfr_before (
		.din(new_net_1480),
		.dout(new_net_1479)
	);

	bfr new_net_1481_bfr_before (
		.din(new_net_1481),
		.dout(new_net_1480)
	);

	bfr new_net_1482_bfr_before (
		.din(new_net_1482),
		.dout(new_net_1481)
	);

	bfr new_net_1483_bfr_before (
		.din(new_net_1483),
		.dout(new_net_1482)
	);

	bfr new_net_1484_bfr_before (
		.din(new_net_1484),
		.dout(new_net_1483)
	);

	bfr new_net_1485_bfr_before (
		.din(new_net_1485),
		.dout(new_net_1484)
	);

	bfr new_net_1486_bfr_before (
		.din(new_net_1486),
		.dout(new_net_1485)
	);

	bfr new_net_1487_bfr_before (
		.din(new_net_1487),
		.dout(new_net_1486)
	);

	bfr new_net_1488_bfr_before (
		.din(new_net_1488),
		.dout(new_net_1487)
	);

	bfr new_net_1489_bfr_before (
		.din(new_net_1489),
		.dout(new_net_1488)
	);

	bfr new_net_1490_bfr_before (
		.din(new_net_1490),
		.dout(new_net_1489)
	);

	bfr new_net_1491_bfr_before (
		.din(new_net_1491),
		.dout(new_net_1490)
	);

	bfr new_net_1492_bfr_before (
		.din(new_net_1492),
		.dout(new_net_1491)
	);

	bfr new_net_1493_bfr_before (
		.din(new_net_1493),
		.dout(new_net_1492)
	);

	bfr new_net_1494_bfr_before (
		.din(new_net_1494),
		.dout(new_net_1493)
	);

	bfr new_net_1495_bfr_before (
		.din(new_net_1495),
		.dout(new_net_1494)
	);

	bfr new_net_1496_bfr_before (
		.din(new_net_1496),
		.dout(new_net_1495)
	);

	bfr new_net_1497_bfr_before (
		.din(new_net_1497),
		.dout(new_net_1496)
	);

	bfr new_net_1498_bfr_before (
		.din(new_net_1498),
		.dout(new_net_1497)
	);

	bfr new_net_1499_bfr_before (
		.din(new_net_1499),
		.dout(new_net_1498)
	);

	bfr new_net_1500_bfr_before (
		.din(new_net_1500),
		.dout(new_net_1499)
	);

	bfr new_net_1501_bfr_before (
		.din(new_net_1501),
		.dout(new_net_1500)
	);

	bfr new_net_1502_bfr_before (
		.din(new_net_1502),
		.dout(new_net_1501)
	);

	bfr new_net_1503_bfr_before (
		.din(new_net_1503),
		.dout(new_net_1502)
	);

	spl2 new_net_575_v_fanout (
		.a(new_net_575),
		.b(new_net_1503),
		.c(new_net_474)
	);

	bfr new_net_1504_bfr_before (
		.din(new_net_1504),
		.dout(new_net_592)
	);

	bfr new_net_1505_bfr_before (
		.din(new_net_1505),
		.dout(new_net_1504)
	);

	bfr new_net_1506_bfr_before (
		.din(new_net_1506),
		.dout(new_net_1505)
	);

	bfr new_net_1507_bfr_before (
		.din(new_net_1507),
		.dout(new_net_1506)
	);

	bfr new_net_1508_bfr_before (
		.din(new_net_1508),
		.dout(new_net_1507)
	);

	bfr new_net_1509_bfr_before (
		.din(new_net_1509),
		.dout(new_net_1508)
	);

	bfr new_net_1510_bfr_before (
		.din(new_net_1510),
		.dout(new_net_1509)
	);

	bfr new_net_1511_bfr_before (
		.din(new_net_1511),
		.dout(new_net_1510)
	);

	bfr new_net_1512_bfr_before (
		.din(new_net_1512),
		.dout(new_net_1511)
	);

	bfr new_net_1513_bfr_before (
		.din(new_net_1513),
		.dout(new_net_1512)
	);

	bfr new_net_1514_bfr_before (
		.din(new_net_1514),
		.dout(new_net_1513)
	);

	bfr new_net_1515_bfr_before (
		.din(new_net_1515),
		.dout(new_net_1514)
	);

	bfr new_net_1516_bfr_before (
		.din(new_net_1516),
		.dout(new_net_1515)
	);

	bfr new_net_1517_bfr_before (
		.din(new_net_1517),
		.dout(new_net_1516)
	);

	bfr new_net_1518_bfr_before (
		.din(new_net_1518),
		.dout(new_net_1517)
	);

	bfr new_net_1519_bfr_before (
		.din(new_net_1519),
		.dout(new_net_1518)
	);

	bfr new_net_1520_bfr_before (
		.din(new_net_1520),
		.dout(new_net_1519)
	);

	bfr new_net_1521_bfr_before (
		.din(new_net_1521),
		.dout(new_net_1520)
	);

	bfr new_net_1522_bfr_before (
		.din(new_net_1522),
		.dout(new_net_1521)
	);

	bfr new_net_1523_bfr_before (
		.din(new_net_1523),
		.dout(new_net_1522)
	);

	bfr new_net_1524_bfr_before (
		.din(new_net_1524),
		.dout(new_net_1523)
	);

	bfr new_net_1525_bfr_before (
		.din(new_net_1525),
		.dout(new_net_1524)
	);

	bfr new_net_1526_bfr_before (
		.din(new_net_1526),
		.dout(new_net_1525)
	);

	bfr new_net_1527_bfr_before (
		.din(new_net_1527),
		.dout(new_net_1526)
	);

	bfr new_net_1528_bfr_before (
		.din(new_net_1528),
		.dout(new_net_1527)
	);

	bfr new_net_1529_bfr_before (
		.din(new_net_1529),
		.dout(new_net_1528)
	);

	spl3L new_net_591_v_fanout (
		.a(new_net_591),
		.b(new_net_150),
		.c(new_net_147),
		.d(new_net_1529)
	);

	spl2 new_net_606_v_fanout (
		.a(new_net_606),
		.b(new_net_408),
		.c(new_net_406)
	);

	bfr new_net_1530_bfr_before (
		.din(new_net_1530),
		.dout(new_net_585)
	);

	bfr new_net_1531_bfr_before (
		.din(new_net_1531),
		.dout(new_net_1530)
	);

	bfr new_net_1532_bfr_before (
		.din(new_net_1532),
		.dout(new_net_1531)
	);

	bfr new_net_1533_bfr_before (
		.din(new_net_1533),
		.dout(new_net_1532)
	);

	bfr new_net_1534_bfr_before (
		.din(new_net_1534),
		.dout(new_net_1533)
	);

	bfr new_net_1535_bfr_before (
		.din(new_net_1535),
		.dout(new_net_1534)
	);

	bfr new_net_1536_bfr_before (
		.din(new_net_1536),
		.dout(new_net_1535)
	);

	bfr new_net_1537_bfr_before (
		.din(new_net_1537),
		.dout(new_net_1536)
	);

	bfr new_net_1538_bfr_before (
		.din(new_net_1538),
		.dout(new_net_1537)
	);

	bfr new_net_1539_bfr_before (
		.din(new_net_1539),
		.dout(new_net_1538)
	);

	bfr new_net_1540_bfr_before (
		.din(new_net_1540),
		.dout(new_net_1539)
	);

	bfr new_net_1541_bfr_before (
		.din(new_net_1541),
		.dout(new_net_1540)
	);

	bfr new_net_1542_bfr_before (
		.din(new_net_1542),
		.dout(new_net_1541)
	);

	bfr new_net_1543_bfr_before (
		.din(new_net_1543),
		.dout(new_net_1542)
	);

	bfr new_net_1544_bfr_before (
		.din(new_net_1544),
		.dout(new_net_1543)
	);

	bfr new_net_1545_bfr_before (
		.din(new_net_1545),
		.dout(new_net_1544)
	);

	bfr new_net_1546_bfr_before (
		.din(new_net_1546),
		.dout(new_net_1545)
	);

	bfr new_net_1547_bfr_before (
		.din(new_net_1547),
		.dout(new_net_1546)
	);

	bfr new_net_1548_bfr_before (
		.din(new_net_1548),
		.dout(new_net_1547)
	);

	bfr new_net_1549_bfr_before (
		.din(new_net_1549),
		.dout(new_net_1548)
	);

	bfr new_net_1550_bfr_before (
		.din(new_net_1550),
		.dout(new_net_1549)
	);

	bfr new_net_1551_bfr_before (
		.din(new_net_1551),
		.dout(new_net_1550)
	);

	bfr new_net_1552_bfr_before (
		.din(new_net_1552),
		.dout(new_net_1551)
	);

	bfr new_net_1553_bfr_before (
		.din(new_net_1553),
		.dout(new_net_1552)
	);

	bfr new_net_1554_bfr_before (
		.din(new_net_1554),
		.dout(new_net_1553)
	);

	bfr new_net_1555_bfr_before (
		.din(new_net_1555),
		.dout(new_net_1554)
	);

	spl3L new_net_587_v_fanout (
		.a(new_net_587),
		.b(new_net_344),
		.c(new_net_341),
		.d(new_net_1555)
	);

	bfr new_net_1556_bfr_before (
		.din(new_net_1556),
		.dout(new_net_648)
	);

	bfr new_net_1557_bfr_before (
		.din(new_net_1557),
		.dout(new_net_1556)
	);

	bfr new_net_1558_bfr_before (
		.din(new_net_1558),
		.dout(new_net_1557)
	);

	bfr new_net_1559_bfr_before (
		.din(new_net_1559),
		.dout(new_net_1558)
	);

	bfr new_net_1560_bfr_before (
		.din(new_net_1560),
		.dout(new_net_1559)
	);

	bfr new_net_1561_bfr_before (
		.din(new_net_1561),
		.dout(new_net_1560)
	);

	bfr new_net_1562_bfr_before (
		.din(new_net_1562),
		.dout(new_net_1561)
	);

	bfr new_net_1563_bfr_before (
		.din(new_net_1563),
		.dout(new_net_1562)
	);

	bfr new_net_1564_bfr_before (
		.din(new_net_1564),
		.dout(new_net_1563)
	);

	bfr new_net_1565_bfr_before (
		.din(new_net_1565),
		.dout(new_net_1564)
	);

	bfr new_net_1566_bfr_before (
		.din(new_net_1566),
		.dout(new_net_1565)
	);

	bfr new_net_1567_bfr_before (
		.din(new_net_1567),
		.dout(new_net_1566)
	);

	bfr new_net_1568_bfr_before (
		.din(new_net_1568),
		.dout(new_net_1567)
	);

	bfr new_net_1569_bfr_before (
		.din(new_net_1569),
		.dout(new_net_1568)
	);

	bfr new_net_1570_bfr_before (
		.din(new_net_1570),
		.dout(new_net_1569)
	);

	bfr new_net_1571_bfr_before (
		.din(new_net_1571),
		.dout(new_net_1570)
	);

	bfr new_net_1572_bfr_before (
		.din(new_net_1572),
		.dout(new_net_1571)
	);

	bfr new_net_1573_bfr_before (
		.din(new_net_1573),
		.dout(new_net_1572)
	);

	bfr new_net_1574_bfr_before (
		.din(new_net_1574),
		.dout(new_net_1573)
	);

	bfr new_net_1575_bfr_before (
		.din(new_net_1575),
		.dout(new_net_1574)
	);

	bfr new_net_1576_bfr_before (
		.din(new_net_1576),
		.dout(new_net_1575)
	);

	bfr new_net_1577_bfr_before (
		.din(new_net_1577),
		.dout(new_net_1576)
	);

	bfr new_net_1578_bfr_before (
		.din(new_net_1578),
		.dout(new_net_1577)
	);

	bfr new_net_1579_bfr_before (
		.din(new_net_1579),
		.dout(new_net_1578)
	);

	bfr new_net_1580_bfr_before (
		.din(new_net_1580),
		.dout(new_net_1579)
	);

	spl2 new_net_649_v_fanout (
		.a(new_net_649),
		.b(new_net_1580),
		.c(new_net_438)
	);

	spl3L new_net_650_v_fanout (
		.a(new_net_650),
		.b(new_net_442),
		.c(new_net_437),
		.d(new_net_440)
	);

	bfr new_net_1581_bfr_before (
		.din(new_net_1581),
		.dout(new_net_619)
	);

	bfr new_net_1582_bfr_before (
		.din(new_net_1582),
		.dout(new_net_1581)
	);

	bfr new_net_1583_bfr_before (
		.din(new_net_1583),
		.dout(new_net_1582)
	);

	bfr new_net_1584_bfr_before (
		.din(new_net_1584),
		.dout(new_net_1583)
	);

	bfr new_net_1585_bfr_before (
		.din(new_net_1585),
		.dout(new_net_1584)
	);

	bfr new_net_1586_bfr_before (
		.din(new_net_1586),
		.dout(new_net_1585)
	);

	bfr new_net_1587_bfr_before (
		.din(new_net_1587),
		.dout(new_net_1586)
	);

	bfr new_net_1588_bfr_before (
		.din(new_net_1588),
		.dout(new_net_1587)
	);

	bfr new_net_1589_bfr_before (
		.din(new_net_1589),
		.dout(new_net_1588)
	);

	bfr new_net_1590_bfr_before (
		.din(new_net_1590),
		.dout(new_net_1589)
	);

	bfr new_net_1591_bfr_before (
		.din(new_net_1591),
		.dout(new_net_1590)
	);

	bfr new_net_1592_bfr_before (
		.din(new_net_1592),
		.dout(new_net_1591)
	);

	bfr new_net_1593_bfr_before (
		.din(new_net_1593),
		.dout(new_net_1592)
	);

	bfr new_net_1594_bfr_before (
		.din(new_net_1594),
		.dout(new_net_1593)
	);

	bfr new_net_1595_bfr_before (
		.din(new_net_1595),
		.dout(new_net_1594)
	);

	bfr new_net_1596_bfr_before (
		.din(new_net_1596),
		.dout(new_net_1595)
	);

	bfr new_net_1597_bfr_before (
		.din(new_net_1597),
		.dout(new_net_1596)
	);

	bfr new_net_1598_bfr_before (
		.din(new_net_1598),
		.dout(new_net_1597)
	);

	bfr new_net_1599_bfr_before (
		.din(new_net_1599),
		.dout(new_net_1598)
	);

	bfr new_net_1600_bfr_before (
		.din(new_net_1600),
		.dout(new_net_1599)
	);

	bfr new_net_1601_bfr_before (
		.din(new_net_1601),
		.dout(new_net_1600)
	);

	bfr new_net_1602_bfr_before (
		.din(new_net_1602),
		.dout(new_net_1601)
	);

	bfr new_net_1603_bfr_before (
		.din(new_net_1603),
		.dout(new_net_1602)
	);

	bfr new_net_1604_bfr_before (
		.din(new_net_1604),
		.dout(new_net_1603)
	);

	bfr new_net_1605_bfr_before (
		.din(new_net_1605),
		.dout(new_net_1604)
	);

	spl3L new_net_621_v_fanout (
		.a(new_net_621),
		.b(new_net_1605),
		.c(new_net_206),
		.d(new_net_211)
	);

	spl2 new_net_638_v_fanout (
		.a(new_net_638),
		.b(new_net_234),
		.c(new_net_233)
	);

	spl3L new_net_601_v_fanout (
		.a(new_net_601),
		.b(new_net_248),
		.c(new_net_247),
		.d(new_net_249)
	);

	bfr new_net_1606_bfr_before (
		.din(new_net_1606),
		.dout(new_net_611)
	);

	bfr new_net_1607_bfr_before (
		.din(new_net_1607),
		.dout(new_net_1606)
	);

	bfr new_net_1608_bfr_before (
		.din(new_net_1608),
		.dout(new_net_1607)
	);

	bfr new_net_1609_bfr_before (
		.din(new_net_1609),
		.dout(new_net_1608)
	);

	bfr new_net_1610_bfr_before (
		.din(new_net_1610),
		.dout(new_net_1609)
	);

	bfr new_net_1611_bfr_before (
		.din(new_net_1611),
		.dout(new_net_1610)
	);

	bfr new_net_1612_bfr_before (
		.din(new_net_1612),
		.dout(new_net_1611)
	);

	bfr new_net_1613_bfr_before (
		.din(new_net_1613),
		.dout(new_net_1612)
	);

	bfr new_net_1614_bfr_before (
		.din(new_net_1614),
		.dout(new_net_1613)
	);

	bfr new_net_1615_bfr_before (
		.din(new_net_1615),
		.dout(new_net_1614)
	);

	bfr new_net_1616_bfr_before (
		.din(new_net_1616),
		.dout(new_net_1615)
	);

	bfr new_net_1617_bfr_before (
		.din(new_net_1617),
		.dout(new_net_1616)
	);

	bfr new_net_1618_bfr_before (
		.din(new_net_1618),
		.dout(new_net_1617)
	);

	bfr new_net_1619_bfr_before (
		.din(new_net_1619),
		.dout(new_net_1618)
	);

	bfr new_net_1620_bfr_before (
		.din(new_net_1620),
		.dout(new_net_1619)
	);

	bfr new_net_1621_bfr_before (
		.din(new_net_1621),
		.dout(new_net_1620)
	);

	bfr new_net_1622_bfr_before (
		.din(new_net_1622),
		.dout(new_net_1621)
	);

	bfr new_net_1623_bfr_before (
		.din(new_net_1623),
		.dout(new_net_1622)
	);

	bfr new_net_1624_bfr_before (
		.din(new_net_1624),
		.dout(new_net_1623)
	);

	bfr new_net_1625_bfr_before (
		.din(new_net_1625),
		.dout(new_net_1624)
	);

	bfr new_net_1626_bfr_before (
		.din(new_net_1626),
		.dout(new_net_1625)
	);

	bfr new_net_1627_bfr_before (
		.din(new_net_1627),
		.dout(new_net_1626)
	);

	bfr new_net_1628_bfr_before (
		.din(new_net_1628),
		.dout(new_net_1627)
	);

	bfr new_net_1629_bfr_before (
		.din(new_net_1629),
		.dout(new_net_1628)
	);

	bfr new_net_1630_bfr_before (
		.din(new_net_1630),
		.dout(new_net_1629)
	);

	spl3L new_net_610_v_fanout (
		.a(new_net_610),
		.b(new_net_1630),
		.c(new_net_260),
		.d(new_net_264)
	);

	spl3L new_net_570_v_fanout (
		.a(new_net_570),
		.b(new_net_181),
		.c(new_net_178),
		.d(new_net_182)
	);

	spl2 new_net_630_v_fanout (
		.a(new_net_630),
		.b(new_net_275),
		.c(new_net_274)
	);

	bfr new_net_1631_bfr_before (
		.din(new_net_1631),
		.dout(new_net_584)
	);

	bfr new_net_1632_bfr_before (
		.din(new_net_1632),
		.dout(new_net_1631)
	);

	bfr new_net_1633_bfr_before (
		.din(new_net_1633),
		.dout(new_net_1632)
	);

	bfr new_net_1634_bfr_before (
		.din(new_net_1634),
		.dout(new_net_1633)
	);

	bfr new_net_1635_bfr_before (
		.din(new_net_1635),
		.dout(new_net_1634)
	);

	bfr new_net_1636_bfr_before (
		.din(new_net_1636),
		.dout(new_net_1635)
	);

	bfr new_net_1637_bfr_before (
		.din(new_net_1637),
		.dout(new_net_1636)
	);

	bfr new_net_1638_bfr_before (
		.din(new_net_1638),
		.dout(new_net_1637)
	);

	bfr new_net_1639_bfr_before (
		.din(new_net_1639),
		.dout(new_net_1638)
	);

	bfr new_net_1640_bfr_before (
		.din(new_net_1640),
		.dout(new_net_1639)
	);

	bfr new_net_1641_bfr_before (
		.din(new_net_1641),
		.dout(new_net_1640)
	);

	bfr new_net_1642_bfr_before (
		.din(new_net_1642),
		.dout(new_net_1641)
	);

	bfr new_net_1643_bfr_before (
		.din(new_net_1643),
		.dout(new_net_1642)
	);

	bfr new_net_1644_bfr_before (
		.din(new_net_1644),
		.dout(new_net_1643)
	);

	bfr new_net_1645_bfr_before (
		.din(new_net_1645),
		.dout(new_net_1644)
	);

	bfr new_net_1646_bfr_before (
		.din(new_net_1646),
		.dout(new_net_1645)
	);

	bfr new_net_1647_bfr_before (
		.din(new_net_1647),
		.dout(new_net_1646)
	);

	bfr new_net_1648_bfr_before (
		.din(new_net_1648),
		.dout(new_net_1647)
	);

	bfr new_net_1649_bfr_before (
		.din(new_net_1649),
		.dout(new_net_1648)
	);

	bfr new_net_1650_bfr_before (
		.din(new_net_1650),
		.dout(new_net_1649)
	);

	bfr new_net_1651_bfr_before (
		.din(new_net_1651),
		.dout(new_net_1650)
	);

	bfr new_net_1652_bfr_before (
		.din(new_net_1652),
		.dout(new_net_1651)
	);

	bfr new_net_1653_bfr_before (
		.din(new_net_1653),
		.dout(new_net_1652)
	);

	bfr new_net_1654_bfr_before (
		.din(new_net_1654),
		.dout(new_net_1653)
	);

	bfr new_net_1655_bfr_before (
		.din(new_net_1655),
		.dout(new_net_1654)
	);

	spl3L new_net_583_v_fanout (
		.a(new_net_583),
		.b(new_net_282),
		.c(new_net_284),
		.d(new_net_1655)
	);

	spl3L new_net_590_v_fanout (
		.a(new_net_590),
		.b(new_net_222),
		.c(new_net_221),
		.d(new_net_223)
	);

	bfr new_net_1656_bfr_before (
		.din(new_net_1656),
		.dout(new_net_654)
	);

	bfr new_net_1657_bfr_before (
		.din(new_net_1657),
		.dout(new_net_1656)
	);

	bfr new_net_1658_bfr_before (
		.din(new_net_1658),
		.dout(new_net_1657)
	);

	bfr new_net_1659_bfr_before (
		.din(new_net_1659),
		.dout(new_net_1658)
	);

	bfr new_net_1660_bfr_before (
		.din(new_net_1660),
		.dout(new_net_1659)
	);

	bfr new_net_1661_bfr_before (
		.din(new_net_1661),
		.dout(new_net_1660)
	);

	bfr new_net_1662_bfr_before (
		.din(new_net_1662),
		.dout(new_net_1661)
	);

	bfr new_net_1663_bfr_before (
		.din(new_net_1663),
		.dout(new_net_1662)
	);

	bfr new_net_1664_bfr_before (
		.din(new_net_1664),
		.dout(new_net_1663)
	);

	bfr new_net_1665_bfr_before (
		.din(new_net_1665),
		.dout(new_net_1664)
	);

	bfr new_net_1666_bfr_before (
		.din(new_net_1666),
		.dout(new_net_1665)
	);

	bfr new_net_1667_bfr_before (
		.din(new_net_1667),
		.dout(new_net_1666)
	);

	bfr new_net_1668_bfr_before (
		.din(new_net_1668),
		.dout(new_net_1667)
	);

	bfr new_net_1669_bfr_before (
		.din(new_net_1669),
		.dout(new_net_1668)
	);

	bfr new_net_1670_bfr_before (
		.din(new_net_1670),
		.dout(new_net_1669)
	);

	bfr new_net_1671_bfr_before (
		.din(new_net_1671),
		.dout(new_net_1670)
	);

	bfr new_net_1672_bfr_before (
		.din(new_net_1672),
		.dout(new_net_1671)
	);

	bfr new_net_1673_bfr_before (
		.din(new_net_1673),
		.dout(new_net_1672)
	);

	bfr new_net_1674_bfr_before (
		.din(new_net_1674),
		.dout(new_net_1673)
	);

	bfr new_net_1675_bfr_before (
		.din(new_net_1675),
		.dout(new_net_1674)
	);

	bfr new_net_1676_bfr_before (
		.din(new_net_1676),
		.dout(new_net_1675)
	);

	bfr new_net_1677_bfr_before (
		.din(new_net_1677),
		.dout(new_net_1676)
	);

	bfr new_net_1678_bfr_before (
		.din(new_net_1678),
		.dout(new_net_1677)
	);

	bfr new_net_1679_bfr_before (
		.din(new_net_1679),
		.dout(new_net_1678)
	);

	bfr new_net_1680_bfr_before (
		.din(new_net_1680),
		.dout(new_net_1679)
	);

	spl3L new_net_656_v_fanout (
		.a(new_net_656),
		.b(new_net_398),
		.c(new_net_1680),
		.d(new_net_396)
	);

	spl2 new_net_652_v_fanout (
		.a(new_net_652),
		.b(new_net_351),
		.c(new_net_350)
	);

	spl2 new_net_581_v_fanout (
		.a(new_net_581),
		.b(new_net_317),
		.c(new_net_319)
	);

	bfr new_net_1681_bfr_before (
		.din(new_net_1681),
		.dout(new_net_602)
	);

	bfr new_net_1682_bfr_before (
		.din(new_net_1682),
		.dout(new_net_1681)
	);

	bfr new_net_1683_bfr_before (
		.din(new_net_1683),
		.dout(new_net_1682)
	);

	bfr new_net_1684_bfr_before (
		.din(new_net_1684),
		.dout(new_net_1683)
	);

	bfr new_net_1685_bfr_before (
		.din(new_net_1685),
		.dout(new_net_1684)
	);

	bfr new_net_1686_bfr_before (
		.din(new_net_1686),
		.dout(new_net_1685)
	);

	bfr new_net_1687_bfr_before (
		.din(new_net_1687),
		.dout(new_net_1686)
	);

	bfr new_net_1688_bfr_before (
		.din(new_net_1688),
		.dout(new_net_1687)
	);

	bfr new_net_1689_bfr_before (
		.din(new_net_1689),
		.dout(new_net_1688)
	);

	bfr new_net_1690_bfr_before (
		.din(new_net_1690),
		.dout(new_net_1689)
	);

	bfr new_net_1691_bfr_before (
		.din(new_net_1691),
		.dout(new_net_1690)
	);

	bfr new_net_1692_bfr_before (
		.din(new_net_1692),
		.dout(new_net_1691)
	);

	bfr new_net_1693_bfr_before (
		.din(new_net_1693),
		.dout(new_net_1692)
	);

	bfr new_net_1694_bfr_before (
		.din(new_net_1694),
		.dout(new_net_1693)
	);

	bfr new_net_1695_bfr_before (
		.din(new_net_1695),
		.dout(new_net_1694)
	);

	bfr new_net_1696_bfr_before (
		.din(new_net_1696),
		.dout(new_net_1695)
	);

	bfr new_net_1697_bfr_before (
		.din(new_net_1697),
		.dout(new_net_1696)
	);

	bfr new_net_1698_bfr_before (
		.din(new_net_1698),
		.dout(new_net_1697)
	);

	bfr new_net_1699_bfr_before (
		.din(new_net_1699),
		.dout(new_net_1698)
	);

	bfr new_net_1700_bfr_before (
		.din(new_net_1700),
		.dout(new_net_1699)
	);

	bfr new_net_1701_bfr_before (
		.din(new_net_1701),
		.dout(new_net_1700)
	);

	bfr new_net_1702_bfr_before (
		.din(new_net_1702),
		.dout(new_net_1701)
	);

	bfr new_net_1703_bfr_before (
		.din(new_net_1703),
		.dout(new_net_1702)
	);

	bfr new_net_1704_bfr_before (
		.din(new_net_1704),
		.dout(new_net_1703)
	);

	bfr new_net_1705_bfr_before (
		.din(new_net_1705),
		.dout(new_net_1704)
	);

	spl3L new_net_604_v_fanout (
		.a(new_net_604),
		.b(new_net_1705),
		.c(new_net_330),
		.d(new_net_326)
	);

	spl2 new_net_620_v_fanout (
		.a(new_net_620),
		.b(new_net_209),
		.c(new_net_207)
	);

	spl2 new_net_594_v_fanout (
		.a(new_net_594),
		.b(new_net_296),
		.c(new_net_300)
	);

	spl2 new_net_586_v_fanout (
		.a(new_net_586),
		.b(new_net_342),
		.c(new_net_345)
	);

	spl2 N37_v_fanout (
		.a(N37),
		.b(new_net_570),
		.c(new_net_569)
	);

	spl2 N17_v_fanout (
		.a(N17),
		.b(new_net_572),
		.c(new_net_573)
	);

	spl2 N69_v_fanout (
		.a(N69),
		.b(new_net_576),
		.c(new_net_575)
	);

	spl2 N29_v_fanout (
		.a(N29),
		.b(new_net_578),
		.c(new_net_579)
	);

	spl2 N5_v_fanout (
		.a(N5),
		.b(new_net_582),
		.c(new_net_581)
	);

	bfr new_net_1706_bfr_before (
		.din(new_net_1706),
		.dout(new_net_281)
	);

	bfr new_net_1707_bfr_before (
		.din(new_net_1707),
		.dout(new_net_283)
	);

	spl3L N85_v_fanout (
		.a(N85),
		.b(new_net_1706),
		.c(new_net_583),
		.d(new_net_1707)
	);

	spl2 N57_v_fanout (
		.a(N57),
		.b(new_net_586),
		.c(new_net_587)
	);

	spl2 N89_v_fanout (
		.a(N89),
		.b(new_net_590),
		.c(new_net_589)
	);

	bfr new_net_1708_bfr_before (
		.din(new_net_1708),
		.dout(new_net_149)
	);

	bfr new_net_1709_bfr_before (
		.din(new_net_1709),
		.dout(new_net_151)
	);

	spl3L N33_v_fanout (
		.a(N33),
		.b(new_net_1709),
		.c(new_net_1708),
		.d(new_net_591)
	);

	spl2 N117_v_fanout (
		.a(N117),
		.b(new_net_595),
		.c(new_net_594)
	);

	spl2 N21_v_fanout (
		.a(N21),
		.b(new_net_598),
		.c(new_net_597)
	);

	spl2 N45_v_fanout (
		.a(N45),
		.b(new_net_600),
		.c(new_net_601)
	);

	spl2 N121_v_fanout (
		.a(N121),
		.b(new_net_604),
		.c(new_net_603)
	);

	spl2 N61_v_fanout (
		.a(N61),
		.b(new_net_606),
		.c(new_net_607)
	);

	bfr new_net_1710_bfr_before (
		.din(new_net_1710),
		.dout(new_net_188)
	);

	bfr new_net_1711_bfr_before (
		.din(new_net_1711),
		.dout(new_net_193)
	);

	spl3L N105_v_fanout (
		.a(N105),
		.b(new_net_1711),
		.c(new_net_1710),
		.d(new_net_608)
	);

	bfr new_net_1712_bfr_before (
		.din(new_net_1712),
		.dout(new_net_261)
	);

	bfr new_net_1713_bfr_before (
		.din(new_net_1713),
		.dout(new_net_265)
	);

	spl3L N113_v_fanout (
		.a(N113),
		.b(new_net_1713),
		.c(new_net_1712),
		.d(new_net_610)
	);

	bfr new_net_1714_bfr_before (
		.din(new_net_1714),
		.dout(new_net_94)
	);

	bfr new_net_1715_bfr_before (
		.din(new_net_1715),
		.dout(new_net_98)
	);

	spl3L N25_v_fanout (
		.a(N25),
		.b(new_net_1715),
		.c(new_net_1714),
		.d(new_net_612)
	);

	spl2 N41_v_fanout (
		.a(N41),
		.b(new_net_615),
		.c(new_net_616)
	);

	bfr new_net_1716_bfr_before (
		.din(new_net_1716),
		.dout(new_net_379)
	);

	bfr new_net_1717_bfr_before (
		.din(new_net_1717),
		.dout(new_net_382)
	);

	spl3L N93_v_fanout (
		.a(N93),
		.b(new_net_1716),
		.c(new_net_617),
		.d(new_net_1717)
	);

	spl2 N77_v_fanout (
		.a(N77),
		.b(new_net_620),
		.c(new_net_621)
	);

	bfr new_net_1718_bfr_before (
		.din(new_net_1718),
		.dout(new_net_367)
	);

	bfr new_net_1719_bfr_before (
		.din(new_net_1719),
		.dout(new_net_370)
	);

	spl3L N125_v_fanout (
		.a(N125),
		.b(new_net_1719),
		.c(new_net_1718),
		.d(new_net_622)
	);

	spl2 N81_v_fanout (
		.a(N81),
		.b(new_net_625),
		.c(new_net_626)
	);

	bfr new_net_1720_bfr_before (
		.din(new_net_1720),
		.dout(new_net_419)
	);

	bfr new_net_1721_bfr_before (
		.din(new_net_1721),
		.dout(new_net_422)
	);

	spl3L N13_v_fanout (
		.a(N13),
		.b(new_net_1720),
		.c(new_net_627),
		.d(new_net_1721)
	);

	spl2 N49_v_fanout (
		.a(N49),
		.b(new_net_631),
		.c(new_net_630)
	);

	bfr new_net_1722_bfr_before (
		.din(new_net_1722),
		.dout(new_net_161)
	);

	bfr new_net_1723_bfr_before (
		.din(new_net_1723),
		.dout(new_net_163)
	);

	spl3L N101_v_fanout (
		.a(N101),
		.b(new_net_1723),
		.c(new_net_1722),
		.d(new_net_632)
	);

	spl2 N9_v_fanout (
		.a(N9),
		.b(new_net_635),
		.c(new_net_636)
	);

	spl2 N109_v_fanout (
		.a(N109),
		.b(new_net_638),
		.c(new_net_639)
	);

	spl2 N1_v_fanout (
		.a(N1),
		.b(new_net_642),
		.c(new_net_641)
	);

	spl2 N137_v_fanout (
		.a(N137),
		.b(new_net_643),
		.c(new_net_644)
	);

	spl2 N73_v_fanout (
		.a(N73),
		.b(new_net_646),
		.c(new_net_647)
	);

	spl2 N65_v_fanout (
		.a(N65),
		.b(new_net_650),
		.c(new_net_649)
	);

	spl2 N53_v_fanout (
		.a(N53),
		.b(new_net_652),
		.c(new_net_653)
	);

	spl2 N97_v_fanout (
		.a(N97),
		.b(new_net_656),
		.c(new_net_655)
	);

	bfr N750_bfr_after (
		.din(new_net_697),
		.dout(N750)
	);

	bfr N743_bfr_after (
		.din(new_net_709),
		.dout(N743)
	);

	bfr N753_bfr_after (
		.din(new_net_691),
		.dout(N753)
	);

	bfr N751_bfr_after (
		.din(new_net_699),
		.dout(N751)
	);

	bfr N741_bfr_after (
		.din(new_net_703),
		.dout(N741)
	);

	bfr N747_bfr_after (
		.din(new_net_711),
		.dout(N747)
	);

	bfr N744_bfr_after (
		.din(new_net_715),
		.dout(N744)
	);

	bfr new_net_1724_bfr_after (
		.din(N135),
		.dout(new_net_1724)
	);

	bfr new_net_672_bfr_after (
		.din(new_net_1724),
		.dout(new_net_672)
	);

	bfr new_net_1725_bfr_after (
		.din(N134),
		.dout(new_net_1725)
	);

	bfr new_net_681_bfr_after (
		.din(new_net_1725),
		.dout(new_net_681)
	);

	bfr new_net_1726_bfr_after (
		.din(_237_),
		.dout(new_net_1726)
	);

	bfr new_net_1727_bfr_after (
		.din(new_net_1726),
		.dout(new_net_1727)
	);

	bfr new_net_682_bfr_after (
		.din(new_net_1727),
		.dout(new_net_682)
	);

	bfr new_net_683_bfr_after (
		.din(_240_),
		.dout(new_net_683)
	);

	bfr new_net_684_bfr_after (
		.din(_241_),
		.dout(new_net_684)
	);

	bfr N740_bfr_after (
		.din(new_net_689),
		.dout(N740)
	);

	bfr N745_bfr_after (
		.din(new_net_693),
		.dout(N745)
	);

	bfr N746_bfr_after (
		.din(new_net_701),
		.dout(N746)
	);

	bfr N749_bfr_after (
		.din(new_net_705),
		.dout(N749)
	);

	bfr N755_bfr_after (
		.din(new_net_713),
		.dout(N755)
	);

	bfr new_net_1728_bfr_after (
		.din(N131),
		.dout(new_net_1728)
	);

	bfr new_net_671_bfr_after (
		.din(new_net_1728),
		.dout(new_net_671)
	);

	bfr N742_bfr_after (
		.din(new_net_685),
		.dout(N742)
	);

	bfr new_net_1729_bfr_after (
		.din(N136),
		.dout(new_net_1729)
	);

	bfr new_net_673_bfr_after (
		.din(new_net_1729),
		.dout(new_net_673)
	);

	bfr new_net_1730_bfr_after (
		.din(N129),
		.dout(new_net_1730)
	);

	bfr new_net_674_bfr_after (
		.din(new_net_1730),
		.dout(new_net_674)
	);

	bfr N748_bfr_after (
		.din(new_net_695),
		.dout(N748)
	);

	bfr N752_bfr_after (
		.din(new_net_707),
		.dout(N752)
	);

	bfr N754_bfr_after (
		.din(new_net_687),
		.dout(N754)
	);

	bfr new_net_1731_bfr_after (
		.din(N130),
		.dout(new_net_1731)
	);

	bfr new_net_675_bfr_after (
		.din(new_net_1731),
		.dout(new_net_675)
	);

	bfr new_net_1732_bfr_after (
		.din(N132),
		.dout(new_net_1732)
	);

	bfr new_net_676_bfr_after (
		.din(new_net_1732),
		.dout(new_net_676)
	);

	bfr new_net_677_bfr_after (
		.din(_172_),
		.dout(new_net_677)
	);

	bfr new_net_1733_bfr_after (
		.din(_174_),
		.dout(new_net_1733)
	);

	bfr new_net_678_bfr_after (
		.din(new_net_1733),
		.dout(new_net_678)
	);

	bfr new_net_1734_bfr_after (
		.din(_175_),
		.dout(new_net_1734)
	);

	bfr new_net_679_bfr_after (
		.din(new_net_1734),
		.dout(new_net_679)
	);

	bfr new_net_1735_bfr_after (
		.din(N133),
		.dout(new_net_1735)
	);

	bfr new_net_680_bfr_after (
		.din(new_net_1735),
		.dout(new_net_680)
	);

endmodule