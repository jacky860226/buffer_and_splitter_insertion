module c7552(N1,N164,N160,N82,N188,N152,N84,N174,N180,N55,N57,N65,N144,N343,N85,N41,N151,N211,N175,N183,N207,N210,N26,N162,N150,N346,N166,N319,N59,N156,N182,N38,N115,N337,N87,N219,N229,N289,N69,N352,N44,N133,N214,N109,N97,N240,N271,N88,N86,N242,N260,N189,N199,N186,N158,N198,N334,N118,N89,N212,N168,N205,N224,N64,N208,N155,N94,N9,N361,N195,N231,N124,N316,N293,N364,N232,N121,N78,N307,N245,N18,N179,N141,N280,N328,N358,N134,N239,N296,N81,N202,N29,N79,N163,N165,N217,N254,N193,N53,N80,N157,N154,N197,N218,N181,N196,N111,N167,N237,N112,N113,N172,N223,N106,N73,N263,N74,N203,N206,N76,N213,N135,N248,N32,N12,N226,N77,N201,N286,N170,N227,N236,N331,N184,N176,N310,N355,N173,N349,N190,N235,N47,N221,N153,N178,N191,N130,N257,N62,N200,N228,N230,N367,N66,N70,N185,N277,N233,N299,N234,N313,N83,N159,N177,N251,N103,N58,N216,N220,N241_I,N187,N60,N267,N204,N325,N15,N75,N303,N61,N171,N56,N340,N322,N138,N194,N23,N161,N54,N225,N283,N147,N127,N110,N274,N100,N222,N382,N238,N169,N35,N5,N114,N50,N209,N215,N192,N63);
    wire n_0944_;
    wire new_Jinkela_wire_9680;
    wire new_Jinkela_wire_5455;
    wire new_Jinkela_wire_6733;
    wire new_Jinkela_wire_8304;
    wire new_Jinkela_wire_5218;
    wire n_0045_;
    wire new_Jinkela_wire_8154;
    wire new_Jinkela_wire_8815;
    wire new_Jinkela_wire_7847;
    wire new_Jinkela_wire_10140;
    wire new_Jinkela_wire_6222;
    wire new_Jinkela_wire_9389;
    wire new_Jinkela_wire_4987;
    wire new_Jinkela_wire_884;
    wire new_Jinkela_wire_3243;
    wire new_Jinkela_wire_8951;
    wire n_0888_;
    wire n_0885_;
    wire new_Jinkela_wire_8919;
    wire new_Jinkela_wire_7138;
    wire new_Jinkela_wire_6116;
    wire new_Jinkela_wire_4404;
    wire new_Jinkela_wire_2254;
    wire new_Jinkela_wire_10287;
    wire n_0992_;
    wire new_Jinkela_wire_4160;
    wire new_Jinkela_wire_8623;
    wire new_Jinkela_wire_6529;
    wire new_Jinkela_wire_3574;
    wire new_Jinkela_wire_10629;
    wire new_Jinkela_wire_5235;
    wire new_Jinkela_wire_6729;
    wire new_Jinkela_wire_1753;
    wire new_Jinkela_wire_4979;
    wire new_Jinkela_wire_7319;
    wire new_Jinkela_wire_3709;
    wire new_Jinkela_wire_2145;
    wire new_Jinkela_wire_4966;
    wire new_Jinkela_wire_3893;
    wire new_Jinkela_wire_9733;
    wire new_Jinkela_wire_1062;
    wire new_Jinkela_wire_318;
    wire new_Jinkela_wire_14;
    wire new_Jinkela_wire_6487;
    wire new_Jinkela_wire_2795;
    wire n_1153_;
    wire new_Jinkela_wire_9783;
    wire new_Jinkela_wire_4056;
    wire new_Jinkela_wire_819;
    wire n_1066_;
    wire new_Jinkela_wire_10046;
    wire new_Jinkela_wire_7108;
    wire new_Jinkela_wire_7643;
    wire new_Jinkela_wire_8437;
    wire new_Jinkela_wire_978;
    wire new_Jinkela_wire_10437;
    wire new_Jinkela_wire_9811;
    wire new_Jinkela_wire_7706;
    wire new_Jinkela_wire_10035;
    wire new_Jinkela_wire_2104;
    wire new_Jinkela_wire_10085;
    wire new_Jinkela_wire_3335;
    wire new_Jinkela_wire_3086;
    wire new_Jinkela_wire_8286;
    wire new_Jinkela_wire_2660;
    wire new_Jinkela_wire_4821;
    wire new_Jinkela_wire_7077;
    wire new_Jinkela_wire_4957;
    wire new_Jinkela_wire_3706;
    wire n_0301_;
    wire new_Jinkela_wire_2808;
    wire n_0215_;
    wire new_Jinkela_wire_7945;
    wire new_Jinkela_wire_5655;
    wire new_Jinkela_wire_8436;
    wire new_Jinkela_wire_731;
    wire new_Jinkela_wire_6967;
    wire new_Jinkela_wire_2831;
    wire new_Jinkela_wire_3902;
    wire new_Jinkela_wire_7661;
    wire new_Jinkela_wire_9309;
    wire new_Jinkela_wire_9373;
    wire new_Jinkela_wire_9862;
    wire new_Jinkela_wire_324;
    wire new_Jinkela_wire_7368;
    wire new_Jinkela_wire_10627;
    wire new_Jinkela_wire_1795;
    wire new_Jinkela_wire_3020;
    wire new_Jinkela_wire_734;
    wire new_Jinkela_wire_8566;
    wire new_Jinkela_wire_2226;
    wire new_Jinkela_wire_6444;
    wire new_Jinkela_wire_1711;
    wire new_Jinkela_wire_6401;
    wire new_Jinkela_wire_5208;
    wire n_1149_;
    wire new_Jinkela_wire_9929;
    wire new_Jinkela_wire_7586;
    wire new_Jinkela_wire_8303;
    wire new_Jinkela_wire_2261;
    wire new_Jinkela_wire_4114;
    wire new_Jinkela_wire_3852;
    wire new_Jinkela_wire_8441;
    wire n_0010_;
    wire new_Jinkela_wire_1232;
    wire new_Jinkela_wire_7505;
    wire new_Jinkela_wire_476;
    wire new_Jinkela_wire_5301;
    wire new_Jinkela_wire_4865;
    wire new_Jinkela_wire_8405;
    wire new_Jinkela_wire_4010;
    wire new_Jinkela_wire_2803;
    wire new_Jinkela_wire_700;
    wire new_Jinkela_wire_5353;
    wire new_Jinkela_wire_1128;
    wire new_Jinkela_wire_3319;
    wire new_Jinkela_wire_113;
    wire new_Jinkela_wire_7009;
    wire new_Jinkela_wire_8221;
    wire new_Jinkela_wire_9252;
    wire new_Jinkela_wire_6845;
    wire new_Jinkela_wire_2887;
    wire new_Jinkela_wire_818;
    wire new_Jinkela_wire_3409;
    wire new_Jinkela_wire_3337;
    wire n_0373_;
    wire new_Jinkela_wire_3876;
    wire new_Jinkela_wire_1285;
    wire new_Jinkela_wire_6689;
    wire new_Jinkela_wire_8321;
    wire new_Jinkela_wire_5884;
    wire new_Jinkela_wire_9857;
    wire n_0745_;
    wire new_Jinkela_wire_8089;
    wire new_Jinkela_wire_4892;
    wire new_Jinkela_wire_6157;
    wire new_net_0;
    wire new_Jinkela_wire_9833;
    wire new_Jinkela_wire_1577;
    wire new_Jinkela_wire_6785;
    wire new_Jinkela_wire_7173;
    wire new_Jinkela_wire_32;
    wire new_Jinkela_wire_5253;
    wire new_Jinkela_wire_9584;
    wire new_Jinkela_wire_599;
    wire new_Jinkela_wire_3602;
    wire new_Jinkela_wire_8272;
    wire new_Jinkela_wire_2019;
    wire new_Jinkela_wire_1749;
    wire new_Jinkela_wire_9568;
    wire new_Jinkela_wire_2465;
    wire n_1290_;
    wire new_Jinkela_wire_3233;
    wire new_Jinkela_wire_1696;
    wire new_Jinkela_wire_8095;
    wire new_Jinkela_wire_10261;
    wire new_Jinkela_wire_8493;
    wire new_Jinkela_wire_369;
    wire new_Jinkela_wire_7157;
    wire new_Jinkela_wire_614;
    wire new_Jinkela_wire_3611;
    wire new_Jinkela_wire_845;
    wire new_Jinkela_wire_1744;
    wire new_Jinkela_wire_3502;
    wire new_Jinkela_wire_5490;
    wire new_Jinkela_wire_902;
    wire new_Jinkela_wire_9560;
    wire new_Jinkela_wire_900;
    wire n_0342_;
    wire new_Jinkela_wire_10243;
    wire new_Jinkela_wire_846;
    wire new_Jinkela_wire_1238;
    wire new_Jinkela_wire_7313;
    wire new_Jinkela_wire_9805;
    wire new_Jinkela_wire_3419;
    wire new_Jinkela_wire_5261;
    wire new_Jinkela_wire_4022;
    wire new_Jinkela_wire_2360;
    wire new_Jinkela_wire_6086;
    wire new_Jinkela_wire_716;
    wire new_Jinkela_wire_8634;
    wire new_Jinkela_wire_5338;
    wire new_Jinkela_wire_7100;
    wire new_Jinkela_wire_8857;
    wire new_Jinkela_wire_2911;
    wire new_Jinkela_wire_6706;
    wire n_1336_;
    wire new_Jinkela_wire_2054;
    wire new_Jinkela_wire_2575;
    wire new_Jinkela_wire_2307;
    wire new_Jinkela_wire_2579;
    wire new_Jinkela_wire_2823;
    wire new_Jinkela_wire_2169;
    wire new_Jinkela_wire_9894;
    wire new_Jinkela_wire_10380;
    wire new_Jinkela_wire_3497;
    wire new_Jinkela_wire_9220;
    wire new_Jinkela_wire_5706;
    wire new_Jinkela_wire_9117;
    wire new_Jinkela_wire_9203;
    wire n_1275_;
    wire n_0550_;
    wire new_Jinkela_wire_9493;
    wire new_Jinkela_wire_10186;
    wire new_Jinkela_wire_5377;
    wire new_Jinkela_wire_7179;
    wire new_Jinkela_wire_3862;
    wire new_Jinkela_wire_8027;
    wire new_Jinkela_wire_7091;
    wire new_Jinkela_wire_10337;
    wire new_Jinkela_wire_9210;
    wire new_Jinkela_wire_4947;
    wire new_Jinkela_wire_3965;
    wire new_Jinkela_wire_8137;
    wire new_Jinkela_wire_6616;
    wire new_Jinkela_wire_6955;
    wire new_Jinkela_wire_2427;
    wire new_Jinkela_wire_6188;
    wire new_Jinkela_wire_6379;
    wire new_Jinkela_wire_10177;
    wire new_Jinkela_wire_8677;
    wire new_Jinkela_wire_937;
    wire new_Jinkela_wire_8230;
    wire n_0561_;
    wire new_Jinkela_wire_1275;
    wire new_Jinkela_wire_7467;
    wire new_Jinkela_wire_1911;
    wire new_Jinkela_wire_3350;
    wire new_Jinkela_wire_6960;
    wire n_0897_;
    wire new_Jinkela_wire_4812;
    wire new_Jinkela_wire_5569;
    wire new_Jinkela_wire_7918;
    wire new_Jinkela_wire_9799;
    wire new_Jinkela_wire_8956;
    wire new_Jinkela_wire_6819;
    wire new_Jinkela_wire_6531;
    wire new_Jinkela_wire_1272;
    wire new_Jinkela_wire_7665;
    wire new_Jinkela_wire_684;
    wire new_Jinkela_wire_3705;
    wire n_0875_;
    wire new_Jinkela_wire_8052;
    wire new_Jinkela_wire_7898;
    wire n_0283_;
    wire new_Jinkela_wire_552;
    wire new_Jinkela_wire_3871;
    wire new_Jinkela_wire_5425;
    wire new_Jinkela_wire_3459;
    wire new_Jinkela_wire_98;
    wire new_Jinkela_wire_4603;
    wire new_Jinkela_wire_4696;
    wire new_Jinkela_wire_4911;
    wire new_Jinkela_wire_1763;
    wire new_Jinkela_wire_2685;
    wire new_Jinkela_wire_8684;
    wire new_Jinkela_wire_6011;
    wire new_Jinkela_wire_264;
    wire new_Jinkela_wire_2703;
    wire n_1201_;
    wire new_Jinkela_wire_5626;
    wire new_Jinkela_wire_9810;
    wire new_Jinkela_wire_390;
    wire new_Jinkela_wire_7471;
    wire new_Jinkela_wire_5685;
    wire new_Jinkela_wire_253;
    wire new_Jinkela_wire_8450;
    wire new_Jinkela_wire_9550;
    wire new_Jinkela_wire_8266;
    wire new_Jinkela_wire_5076;
    wire new_Jinkela_wire_7893;
    wire n_1176_;
    wire new_Jinkela_wire_1236;
    wire n_0573_;
    wire new_Jinkela_wire_8739;
    wire new_Jinkela_wire_1005;
    wire new_Jinkela_wire_10463;
    wire new_Jinkela_wire_370;
    wire new_Jinkela_wire_9784;
    wire new_Jinkela_wire_8480;
    wire new_Jinkela_wire_1207;
    wire new_Jinkela_wire_8442;
    wire new_Jinkela_wire_6288;
    wire new_Jinkela_wire_5787;
    wire new_Jinkela_wire_6194;
    wire new_Jinkela_wire_4978;
    wire new_Jinkela_wire_3578;
    wire new_Jinkela_wire_7535;
    wire new_Jinkela_wire_2603;
    wire new_Jinkela_wire_1598;
    wire new_Jinkela_wire_9551;
    wire new_Jinkela_wire_8967;
    wire new_Jinkela_wire_10003;
    wire new_Jinkela_wire_6899;
    wire new_Jinkela_wire_2988;
    wire new_Jinkela_wire_1220;
    wire new_Jinkela_wire_8625;
    wire new_Jinkela_wire_1142;
    wire new_Jinkela_wire_40;
    wire new_Jinkela_wire_6266;
    wire new_Jinkela_wire_51;
    wire new_Jinkela_wire_3390;
    wire new_Jinkela_wire_7215;
    wire new_Jinkela_wire_8123;
    wire new_Jinkela_wire_2820;
    wire new_Jinkela_wire_10250;
    wire n_0064_;
    wire new_Jinkela_wire_6408;
    wire new_Jinkela_wire_4650;
    wire n_1158_;
    wire new_Jinkela_wire_5497;
    wire new_Jinkela_wire_2880;
    wire new_Jinkela_wire_7614;
    wire new_Jinkela_wire_6773;
    wire new_Jinkela_wire_1333;
    wire n_0007_;
    wire new_Jinkela_wire_7111;
    wire n_0708_;
    wire new_Jinkela_wire_4789;
    wire new_Jinkela_wire_6981;
    wire new_Jinkela_wire_9677;
    wire new_Jinkela_wire_3078;
    wire n_0317_;
    wire new_Jinkela_wire_8531;
    wire n_1371_;
    wire new_Jinkela_wire_7705;
    wire new_Jinkela_wire_5758;
    wire new_Jinkela_wire_7843;
    wire n_0304_;
    wire new_Jinkela_wire_8273;
    wire new_Jinkela_wire_4576;
    wire new_Jinkela_wire_10398;
    wire new_Jinkela_wire_2679;
    wire new_Jinkela_wire_6508;
    wire n_1285_;
    wire n_0463_;
    wire new_Jinkela_wire_1258;
    wire new_Jinkela_wire_196;
    wire new_Jinkela_wire_6510;
    wire n_0900_;
    wire new_Jinkela_wire_1554;
    wire new_Jinkela_wire_1454;
    wire new_Jinkela_wire_10490;
    wire new_Jinkela_wire_6132;
    wire new_Jinkela_wire_9119;
    wire new_Jinkela_wire_2406;
    wire n_0080_;
    wire new_Jinkela_wire_5546;
    wire new_Jinkela_wire_6566;
    wire n_0942_;
    wire new_Jinkela_wire_721;
    wire new_Jinkela_wire_5586;
    wire new_Jinkela_wire_299;
    wire new_Jinkela_wire_5834;
    wire new_Jinkela_wire_10461;
    wire new_Jinkela_wire_3532;
    wire new_Jinkela_wire_5726;
    wire new_Jinkela_wire_6929;
    wire new_Jinkela_wire_9124;
    wire new_Jinkela_wire_2070;
    wire n_0912_;
    wire new_Jinkela_wire_6811;
    wire new_Jinkela_wire_5198;
    wire new_Jinkela_wire_6470;
    wire new_Jinkela_wire_2443;
    wire new_Jinkela_wire_719;
    wire n_0866_;
    wire new_Jinkela_wire_7676;
    wire n_0450_;
    wire new_Jinkela_wire_7636;
    wire new_Jinkela_wire_9655;
    wire new_Jinkela_wire_3842;
    wire new_Jinkela_wire_8314;
    wire new_Jinkela_wire_2917;
    wire new_Jinkela_wire_6290;
    wire new_Jinkela_wire_232;
    wire new_Jinkela_wire_2620;
    wire new_Jinkela_wire_1417;
    wire new_Jinkela_wire_6662;
    wire new_Jinkela_wire_2742;
    wire new_Jinkela_wire_8646;
    wire new_Jinkela_wire_2905;
    wire new_Jinkela_wire_1459;
    wire new_Jinkela_wire_2256;
    wire n_1306_;
    wire new_Jinkela_wire_8582;
    wire new_Jinkela_wire_2001;
    wire n_0272_;
    wire n_1207_;
    wire new_Jinkela_wire_8990;
    wire new_Jinkela_wire_5239;
    wire n_1097_;
    wire new_Jinkela_wire_7678;
    wire new_Jinkela_wire_3289;
    wire new_Jinkela_wire_6059;
    wire new_Jinkela_wire_617;
    wire new_Jinkela_wire_5679;
    wire new_Jinkela_wire_9668;
    wire new_Jinkela_wire_10229;
    wire new_Jinkela_wire_7369;
    wire new_Jinkela_wire_1772;
    wire new_Jinkela_wire_6518;
    wire new_Jinkela_wire_3825;
    wire new_Jinkela_wire_7333;
    wire new_Jinkela_wire_8517;
    wire new_Jinkela_wire_4343;
    wire new_Jinkela_wire_4327;
    wire new_Jinkela_wire_10570;
    wire new_Jinkela_wire_6622;
    wire new_Jinkela_wire_7832;
    wire new_Jinkela_wire_9581;
    wire new_Jinkela_wire_9228;
    wire new_Jinkela_wire_101;
    wire new_Jinkela_wire_7696;
    wire new_Jinkela_wire_10567;
    wire new_Jinkela_wire_4848;
    wire new_Jinkela_wire_4899;
    wire new_Jinkela_wire_5290;
    wire new_Jinkela_wire_2334;
    wire new_Jinkela_wire_6407;
    wire new_Jinkela_wire_1727;
    wire new_Jinkela_wire_7592;
    wire new_Jinkela_wire_490;
    wire new_Jinkela_wire_4918;
    wire n_0569_;
    wire new_Jinkela_wire_7704;
    wire new_Jinkela_wire_9038;
    wire new_Jinkela_wire_1355;
    wire new_Jinkela_wire_7714;
    wire new_Jinkela_wire_6355;
    wire new_Jinkela_wire_10346;
    wire new_Jinkela_wire_5742;
    wire new_Jinkela_wire_8848;
    wire new_Jinkela_wire_5719;
    wire new_Jinkela_wire_224;
    wire new_Jinkela_wire_4658;
    wire new_Jinkela_wire_259;
    wire new_Jinkela_wire_5611;
    wire new_Jinkela_wire_3353;
    wire new_Jinkela_wire_6264;
    wire n_1346_;
    wire new_Jinkela_wire_2107;
    wire new_Jinkela_wire_9869;
    wire new_Jinkela_wire_8828;
    wire new_Jinkela_wire_1054;
    wire new_Jinkela_wire_5542;
    wire n_0528_;
    wire new_Jinkela_wire_9594;
    wire n_0170_;
    wire new_Jinkela_wire_6499;
    wire new_Jinkela_wire_9899;
    wire new_Jinkela_wire_3364;
    wire new_Jinkela_wire_6574;
    wire new_Jinkela_wire_9616;
    wire new_Jinkela_wire_6377;
    wire n_1314_;
    wire n_0600_;
    wire new_Jinkela_wire_3771;
    wire new_Jinkela_wire_7201;
    wire new_Jinkela_wire_5465;
    wire new_Jinkela_wire_7825;
    wire n_0331_;
    wire new_Jinkela_wire_3470;
    wire new_Jinkela_wire_6415;
    wire new_Jinkela_wire_1383;
    wire new_Jinkela_wire_2504;
    wire new_Jinkela_wire_395;
    wire new_Jinkela_wire_9269;
    wire new_Jinkela_wire_9916;
    wire new_Jinkela_wire_9096;
    wire new_Jinkela_wire_5937;
    wire new_Jinkela_wire_6709;
    wire new_Jinkela_wire_8076;
    wire n_0534_;
    wire new_Jinkela_wire_5050;
    wire new_Jinkela_wire_8518;
    wire new_Jinkela_wire_8502;
    wire new_Jinkela_wire_291;
    wire new_Jinkela_wire_5745;
    wire new_Jinkela_wire_5150;
    wire new_Jinkela_wire_5737;
    wire new_Jinkela_wire_7709;
    wire new_Jinkela_wire_544;
    wire new_Jinkela_wire_7999;
    wire new_Jinkela_wire_250;
    wire new_Jinkela_wire_3682;
    wire new_Jinkela_wire_5199;
    wire new_Jinkela_wire_5574;
    wire new_Jinkela_wire_9271;
    wire new_Jinkela_wire_8906;
    wire new_Jinkela_wire_3413;
    wire new_Jinkela_wire_3219;
    wire new_Jinkela_wire_8981;
    wire new_Jinkela_wire_6242;
    wire new_Jinkela_wire_9287;
    wire n_0129_;
    wire new_Jinkela_wire_7141;
    wire new_Jinkela_wire_6972;
    wire new_Jinkela_wire_3410;
    wire n_0347_;
    wire new_Jinkela_wire_448;
    wire new_Jinkela_wire_10073;
    wire new_Jinkela_wire_412;
    wire n_0478_;
    wire new_Jinkela_wire_10377;
    wire new_Jinkela_wire_10476;
    wire new_Jinkela_wire_5312;
    wire new_Jinkela_wire_5762;
    wire new_Jinkela_wire_807;
    wire new_Jinkela_wire_10319;
    wire new_Jinkela_wire_8193;
    wire new_Jinkela_wire_50;
    wire new_Jinkela_wire_5518;
    wire new_Jinkela_wire_8730;
    wire new_Jinkela_wire_10477;
    wire new_Jinkela_wire_2049;
    wire new_Jinkela_wire_4808;
    wire new_Jinkela_wire_2855;
    wire n_0328_;
    wire new_Jinkela_wire_6672;
    wire new_Jinkela_wire_5881;
    wire new_Jinkela_wire_8832;
    wire new_Jinkela_wire_3967;
    wire new_Jinkela_wire_6888;
    wire n_0542_;
    wire new_Jinkela_wire_10305;
    wire new_Jinkela_wire_7443;
    wire new_Jinkela_wire_6799;
    wire new_Jinkela_wire_2392;
    wire new_Jinkela_wire_8243;
    wire n_0635_;
    wire n_0877_;
    wire new_Jinkela_wire_2355;
    wire new_Jinkela_wire_2304;
    wire n_1172_;
    wire new_Jinkela_wire_7854;
    wire new_Jinkela_wire_4852;
    wire n_1227_;
    wire new_Jinkela_wire_9628;
    wire new_Jinkela_wire_7747;
    wire n_1205_;
    wire new_Jinkela_wire_3834;
    wire new_Jinkela_wire_9112;
    wire new_Jinkela_wire_8100;
    wire new_Jinkela_wire_1811;
    wire new_Jinkela_wire_7638;
    wire new_Jinkela_wire_5785;
    wire new_Jinkela_wire_9122;
    wire new_Jinkela_wire_8490;
    wire new_Jinkela_wire_8059;
    wire new_Jinkela_wire_4088;
    wire new_Jinkela_wire_3521;
    wire n_0271_;
    wire new_Jinkela_wire_4856;
    wire n_0926_;
    wire n_0486_;
    wire new_Jinkela_wire_306;
    wire new_Jinkela_wire_9874;
    wire new_Jinkela_wire_5205;
    wire new_Jinkela_wire_4019;
    wire n_0522_;
    wire new_Jinkela_wire_2172;
    wire new_Jinkela_wire_676;
    wire new_Jinkela_wire_4857;
    wire new_Jinkela_wire_5663;
    wire new_Jinkela_wire_843;
    wire new_Jinkela_wire_9240;
    wire new_Jinkela_wire_244;
    wire new_Jinkela_wire_2474;
    wire new_Jinkela_wire_5718;
    wire new_Jinkela_wire_4394;
    wire new_Jinkela_wire_6783;
    wire new_Jinkela_wire_1541;
    wire new_Jinkela_wire_4864;
    wire new_Jinkela_wire_3779;
    wire new_Jinkela_wire_8462;
    wire new_Jinkela_wire_3012;
    wire new_Jinkela_wire_6750;
    wire n_0290_;
    wire n_0899_;
    wire new_Jinkela_wire_8521;
    wire n_0699_;
    wire new_Jinkela_wire_2384;
    wire new_Jinkela_wire_3355;
    wire new_Jinkela_wire_3547;
    wire new_Jinkela_wire_9672;
    wire new_Jinkela_wire_4480;
    wire new_Jinkela_wire_2537;
    wire new_Jinkela_wire_10397;
    wire new_Jinkela_wire_9746;
    wire new_Jinkela_wire_4033;
    wire new_Jinkela_wire_4231;
    wire n_0107_;
    wire new_Jinkela_wire_8445;
    wire new_Jinkela_wire_4244;
    wire new_Jinkela_wire_4965;
    wire new_Jinkela_wire_1560;
    wire new_Jinkela_wire_1444;
    wire new_Jinkela_wire_1155;
    wire new_Jinkela_wire_4230;
    wire new_Jinkela_wire_597;
    wire new_Jinkela_wire_4525;
    wire new_Jinkela_wire_2025;
    wire new_Jinkela_wire_9860;
    wire new_Jinkela_wire_3235;
    wire new_Jinkela_wire_9767;
    wire new_Jinkela_wire_6277;
    wire new_Jinkela_wire_9482;
    wire new_Jinkela_wire_3313;
    wire new_Jinkela_wire_4945;
    wire new_Jinkela_wire_5659;
    wire new_Jinkela_wire_3926;
    wire new_Jinkela_wire_781;
    wire new_Jinkela_wire_4392;
    wire new_Jinkela_wire_4173;
    wire new_Jinkela_wire_9025;
    wire new_Jinkela_wire_8529;
    wire new_Jinkela_wire_8880;
    wire new_Jinkela_wire_6949;
    wire new_Jinkela_wire_7023;
    wire n_1098_;
    wire new_Jinkela_wire_8203;
    wire new_Jinkela_wire_2448;
    wire new_Jinkela_wire_2325;
    wire n_0069_;
    wire new_Jinkela_wire_10394;
    wire new_Jinkela_wire_9849;
    wire n_1058_;
    wire new_Jinkela_wire_3155;
    wire new_Jinkela_wire_3156;
    wire new_Jinkela_wire_1650;
    wire new_Jinkela_wire_2976;
    wire n_0764_;
    wire new_Jinkela_wire_2758;
    wire new_Jinkela_wire_4921;
    wire new_Jinkela_wire_6087;
    wire new_Jinkela_wire_8367;
    wire new_Jinkela_wire_9687;
    wire new_Jinkela_wire_8574;
    wire new_Jinkela_wire_8269;
    wire new_Jinkela_wire_437;
    wire new_Jinkela_wire_1320;
    wire n_0818_;
    wire new_Jinkela_wire_241;
    wire new_Jinkela_wire_2223;
    wire new_Jinkela_wire_3028;
    wire new_Jinkela_wire_10326;
    wire new_Jinkela_wire_2190;
    wire new_Jinkela_wire_4323;
    wire new_Jinkela_wire_3822;
    wire new_Jinkela_wire_9786;
    wire n_0126_;
    wire new_Jinkela_wire_4756;
    wire new_Jinkela_wire_9383;
    wire new_Jinkela_wire_7923;
    wire new_Jinkela_wire_4508;
    wire new_Jinkela_wire_6630;
    wire new_Jinkela_wire_7349;
    wire new_Jinkela_wire_8520;
    wire new_Jinkela_wire_2036;
    wire new_Jinkela_wire_2011;
    wire new_Jinkela_wire_2408;
    wire new_Jinkela_wire_1852;
    wire new_Jinkela_wire_1124;
    wire new_Jinkela_wire_1051;
    wire new_Jinkela_wire_5658;
    wire new_Jinkela_wire_2550;
    wire new_Jinkela_wire_3585;
    wire new_Jinkela_wire_3462;
    wire new_Jinkela_wire_10547;
    wire new_Jinkela_wire_1378;
    wire new_Jinkela_wire_2541;
    wire new_Jinkela_wire_7561;
    wire new_Jinkela_wire_8936;
    wire new_Jinkela_wire_7293;
    wire new_Jinkela_wire_2449;
    wire new_Jinkela_wire_2616;
    wire n_1199_;
    wire new_Jinkela_wire_4397;
    wire new_Jinkela_wire_4407;
    wire new_Jinkela_wire_3473;
    wire new_Jinkela_wire_457;
    wire new_Jinkela_wire_3221;
    wire new_Jinkela_wire_806;
    wire new_Jinkela_wire_5641;
    wire new_Jinkela_wire_63;
    wire new_Jinkela_wire_635;
    wire new_Jinkela_wire_1467;
    wire new_Jinkela_wire_8339;
    wire new_Jinkela_wire_6323;
    wire new_Jinkela_wire_5677;
    wire new_Jinkela_wire_2813;
    wire new_Jinkela_wire_5398;
    wire new_Jinkela_wire_7776;
    wire new_Jinkela_wire_3043;
    wire new_Jinkela_wire_5615;
    wire new_Jinkela_wire_10175;
    wire new_Jinkela_wire_5154;
    wire new_Jinkela_wire_4213;
    wire new_Jinkela_wire_5575;
    wire new_Jinkela_wire_1116;
    wire n_0595_;
    wire new_Jinkela_wire_5624;
    wire new_Jinkela_wire_7559;
    wire new_Jinkela_wire_1974;
    wire new_Jinkela_wire_2565;
    wire new_Jinkela_wire_8156;
    wire new_Jinkela_wire_10221;
    wire new_Jinkela_wire_4541;
    wire new_Jinkela_wire_1901;
    wire new_Jinkela_wire_10575;
    wire new_Jinkela_wire_7083;
    wire n_0761_;
    wire new_Jinkela_wire_1359;
    wire new_Jinkela_wire_7380;
    wire new_Jinkela_wire_362;
    wire new_Jinkela_wire_5964;
    wire new_Jinkela_wire_8169;
    wire n_1262_;
    wire new_Jinkela_wire_7163;
    wire new_Jinkela_wire_1247;
    wire new_Jinkela_wire_2041;
    wire new_Jinkela_wire_8935;
    wire new_Jinkela_wire_10040;
    wire new_Jinkela_wire_1637;
    wire new_Jinkela_wire_6660;
    wire new_Jinkela_wire_7458;
    wire new_Jinkela_wire_7668;
    wire new_Jinkela_wire_1171;
    wire new_Jinkela_wire_6569;
    wire new_Jinkela_wire_10185;
    wire new_Jinkela_wire_2502;
    wire new_Jinkela_wire_5596;
    wire new_Jinkela_wire_1399;
    wire new_Jinkela_wire_756;
    wire n_0119_;
    wire new_Jinkela_wire_7974;
    wire new_Jinkela_wire_286;
    wire new_Jinkela_wire_236;
    wire new_Jinkela_wire_5236;
    wire new_Jinkela_wire_8066;
    wire new_Jinkela_wire_7619;
    wire new_Jinkela_wire_9132;
    wire new_Jinkela_wire_9356;
    wire new_Jinkela_wire_4683;
    wire new_Jinkela_wire_4101;
    wire new_Jinkela_wire_9331;
    wire new_Jinkela_wire_8870;
    wire new_Jinkela_wire_8852;
    wire new_Jinkela_wire_7842;
    wire n_1303_;
    wire new_Jinkela_wire_9270;
    wire new_net_2535;
    wire new_Jinkela_wire_2842;
    wire new_Jinkela_wire_2002;
    wire n_1311_;
    wire n_0366_;
    wire new_Jinkela_wire_5727;
    wire new_Jinkela_wire_7759;
    wire new_Jinkela_wire_10146;
    wire new_Jinkela_wire_7261;
    wire new_Jinkela_wire_6581;
    wire n_0587_;
    wire new_Jinkela_wire_3113;
    wire new_Jinkela_wire_8750;
    wire n_0663_;
    wire new_Jinkela_wire_1648;
    wire new_Jinkela_wire_8587;
    wire new_Jinkela_wire_8255;
    wire new_Jinkela_wire_9130;
    wire new_Jinkela_wire_3316;
    wire new_Jinkela_wire_7960;
    wire new_Jinkela_wire_6973;
    wire n_0767_;
    wire new_Jinkela_wire_4704;
    wire new_Jinkela_wire_3160;
    wire new_Jinkela_wire_2948;
    wire new_Jinkela_wire_4641;
    wire new_Jinkela_wire_6860;
    wire new_Jinkela_wire_7057;
    wire new_Jinkela_wire_4301;
    wire new_Jinkela_wire_715;
    wire new_Jinkela_wire_7254;
    wire new_Jinkela_wire_630;
    wire new_Jinkela_wire_5475;
    wire n_0951_;
    wire new_Jinkela_wire_3704;
    wire new_Jinkela_wire_10267;
    wire new_Jinkela_wire_5500;
    wire new_Jinkela_wire_8639;
    wire n_0812_;
    wire new_Jinkela_wire_2397;
    wire n_0199_;
    wire new_Jinkela_wire_5178;
    wire new_Jinkela_wire_6374;
    wire new_Jinkela_wire_959;
    wire new_Jinkela_wire_6115;
    wire n_0252_;
    wire new_Jinkela_wire_2188;
    wire new_Jinkela_wire_4004;
    wire new_Jinkela_wire_10282;
    wire new_Jinkela_wire_833;
    wire new_Jinkela_wire_7727;
    wire new_Jinkela_wire_1070;
    wire new_Jinkela_wire_2067;
    wire n_1204_;
    wire new_Jinkela_wire_970;
    wire n_1018_;
    wire new_Jinkela_wire_8836;
    wire n_0946_;
    wire new_Jinkela_wire_72;
    wire new_Jinkela_wire_5123;
    wire new_Jinkela_wire_2423;
    wire new_Jinkela_wire_8571;
    wire new_Jinkela_wire_1437;
    wire new_Jinkela_wire_561;
    wire new_Jinkela_wire_3836;
    wire new_Jinkela_wire_4553;
    wire new_net_2531;
    wire new_Jinkela_wire_1991;
    wire new_Jinkela_wire_4209;
    wire new_Jinkela_wire_6595;
    wire new_Jinkela_wire_2092;
    wire new_Jinkela_wire_3345;
    wire new_Jinkela_wire_10211;
    wire new_Jinkela_wire_1756;
    wire new_Jinkela_wire_2784;
    wire new_Jinkela_wire_4993;
    wire new_Jinkela_wire_718;
    wire new_Jinkela_wire_5501;
    wire new_Jinkela_wire_6890;
    wire new_Jinkela_wire_8264;
    wire new_Jinkela_wire_2997;
    wire new_Jinkela_wire_4330;
    wire new_Jinkela_wire_10128;
    wire new_Jinkela_wire_3541;
    wire new_Jinkela_wire_7927;
    wire new_Jinkela_wire_5856;
    wire n_1140_;
    wire new_Jinkela_wire_9496;
    wire new_Jinkela_wire_4123;
    wire new_Jinkela_wire_6505;
    wire new_Jinkela_wire_9091;
    wire new_Jinkela_wire_4374;
    wire new_Jinkela_wire_3568;
    wire new_Jinkela_wire_6137;
    wire new_Jinkela_wire_10404;
    wire new_Jinkela_wire_1832;
    wire new_Jinkela_wire_2840;
    wire new_Jinkela_wire_10270;
    wire n_0982_;
    wire new_Jinkela_wire_4023;
    wire new_Jinkela_wire_3123;
    wire new_Jinkela_wire_6335;
    wire new_Jinkela_wire_9159;
    wire new_Jinkela_wire_9488;
    wire n_0658_;
    wire new_Jinkela_wire_9962;
    wire n_0963_;
    wire new_Jinkela_wire_6614;
    wire new_Jinkela_wire_3479;
    wire n_0607_;
    wire new_Jinkela_wire_9497;
    wire n_0075_;
    wire new_Jinkela_wire_5296;
    wire new_Jinkela_wire_539;
    wire new_Jinkela_wire_9756;
    wire new_Jinkela_wire_7035;
    wire new_Jinkela_wire_4265;
    wire new_Jinkela_wire_6721;
    wire new_Jinkela_wire_503;
    wire new_Jinkela_wire_6107;
    wire new_Jinkela_wire_6442;
    wire new_Jinkela_wire_1602;
    wire n_0294_;
    wire new_Jinkela_wire_9741;
    wire new_Jinkela_wire_8276;
    wire new_Jinkela_wire_5670;
    wire new_Jinkela_wire_3391;
    wire new_Jinkela_wire_4513;
    wire new_Jinkela_wire_7408;
    wire new_Jinkela_wire_1792;
    wire new_Jinkela_wire_10205;
    wire new_Jinkela_wire_6650;
    wire new_Jinkela_wire_9104;
    wire new_Jinkela_wire_3217;
    wire new_Jinkela_wire_6006;
    wire n_0985_;
    wire new_Jinkela_wire_3056;
    wire new_Jinkela_wire_7131;
    wire new_Jinkela_wire_1088;
    wire new_Jinkela_wire_4883;
    wire new_Jinkela_wire_6802;
    wire new_Jinkela_wire_4006;
    wire n_0082_;
    wire new_Jinkela_wire_7949;
    wire new_Jinkela_wire_141;
    wire new_Jinkela_wire_10413;
    wire new_Jinkela_wire_7266;
    wire new_Jinkela_wire_3154;
    wire new_Jinkela_wire_5738;
    wire new_Jinkela_wire_3443;
    wire new_Jinkela_wire_8806;
    wire n_0776_;
    wire new_Jinkela_wire_9189;
    wire new_Jinkela_wire_192;
    wire new_Jinkela_wire_5894;
    wire new_Jinkela_wire_8559;
    wire new_Jinkela_wire_5968;
    wire new_Jinkela_wire_9031;
    wire new_Jinkela_wire_1886;
    wire new_Jinkela_wire_3527;
    wire new_Jinkela_wire_805;
    wire new_Jinkela_wire_3130;
    wire new_Jinkela_wire_9150;
    wire new_Jinkela_wire_8192;
    wire new_Jinkela_wire_2929;
    wire new_Jinkela_wire_3019;
    wire n_0721_;
    wire new_Jinkela_wire_5147;
    wire new_Jinkela_wire_5819;
    wire new_Jinkela_wire_1645;
    wire new_Jinkela_wire_7005;
    wire new_Jinkela_wire_6025;
    wire new_Jinkela_wire_774;
    wire new_Jinkela_wire_6769;
    wire new_Jinkela_wire_9466;
    wire new_Jinkela_wire_8885;
    wire new_Jinkela_wire_6324;
    wire new_Jinkela_wire_3618;
    wire new_Jinkela_wire_10468;
    wire new_Jinkela_wire_6483;
    wire new_Jinkela_wire_4902;
    wire new_Jinkela_wire_5774;
    wire new_Jinkela_wire_465;
    wire new_Jinkela_wire_187;
    wire new_Jinkela_wire_5608;
    wire n_0709_;
    wire new_Jinkela_wire_8309;
    wire new_Jinkela_wire_2928;
    wire new_Jinkela_wire_9557;
    wire new_Jinkela_wire_9543;
    wire new_Jinkela_wire_678;
    wire new_Jinkela_wire_4819;
    wire new_Jinkela_wire_5908;
    wire new_Jinkela_wire_7122;
    wire new_Jinkela_wire_2034;
    wire new_Jinkela_wire_9347;
    wire new_Jinkela_wire_6048;
    wire n_1059_;
    wire new_Jinkela_wire_3576;
    wire new_Jinkela_wire_1607;
    wire n_0343_;
    wire new_Jinkela_wire_1781;
    wire new_Jinkela_wire_8595;
    wire new_Jinkela_wire_5664;
    wire n_0316_;
    wire new_Jinkela_wire_4542;
    wire new_Jinkela_wire_7525;
    wire new_Jinkela_wire_8596;
    wire n_0454_;
    wire n_0844_;
    wire new_Jinkela_wire_9625;
    wire new_Jinkela_wire_400;
    wire new_Jinkela_wire_1686;
    wire new_Jinkela_wire_5167;
    wire new_Jinkela_wire_5292;
    wire n_0650_;
    wire new_Jinkela_wire_2451;
    wire new_Jinkela_wire_8789;
    wire new_Jinkela_wire_3819;
    wire new_Jinkela_wire_10093;
    wire new_Jinkela_wire_1990;
    wire new_Jinkela_wire_2458;
    wire new_Jinkela_wire_6240;
    wire new_Jinkela_wire_500;
    wire new_Jinkela_wire_1948;
    wire new_Jinkela_wire_4194;
    wire new_Jinkela_wire_887;
    wire new_Jinkela_wire_367;
    wire new_Jinkela_wire_9790;
    wire new_Jinkela_wire_9230;
    wire new_Jinkela_wire_939;
    wire n_1322_;
    wire new_Jinkela_wire_3352;
    wire new_Jinkela_wire_2110;
    wire new_Jinkela_wire_5948;
    wire new_Jinkela_wire_2966;
    wire new_Jinkela_wire_3016;
    wire new_Jinkela_wire_1782;
    wire new_Jinkela_wire_4174;
    wire n_0056_;
    wire new_Jinkela_wire_8393;
    wire new_Jinkela_wire_10498;
    wire new_Jinkela_wire_8475;
    wire new_Jinkela_wire_246;
    wire n_1216_;
    wire new_Jinkela_wire_6939;
    wire new_Jinkela_wire_9859;
    wire new_Jinkela_wire_135;
    wire new_Jinkela_wire_6053;
    wire new_Jinkela_wire_1386;
    wire new_Jinkela_wire_389;
    wire new_Jinkela_wire_2330;
    wire new_Jinkela_wire_1697;
    wire new_Jinkela_wire_5530;
    wire new_Jinkela_wire_3537;
    wire new_Jinkela_wire_2003;
    wire new_Jinkela_wire_1506;
    wire new_Jinkela_wire_116;
    wire new_Jinkela_wire_671;
    wire new_Jinkela_wire_905;
    wire new_Jinkela_wire_663;
    wire new_Jinkela_wire_9315;
    wire new_Jinkela_wire_7658;
    wire new_Jinkela_wire_1512;
    wire new_Jinkela_wire_9834;
    wire new_Jinkela_wire_8205;
    wire new_Jinkela_wire_9841;
    wire new_Jinkela_wire_7710;
    wire new_Jinkela_wire_1561;
    wire new_Jinkela_wire_3386;
    wire new_Jinkela_wire_7118;
    wire new_Jinkela_wire_8770;
    wire new_Jinkela_wire_5287;
    wire new_Jinkela_wire_10594;
    wire new_Jinkela_wire_6786;
    wire new_Jinkela_wire_5105;
    wire new_Jinkela_wire_2459;
    wire new_Jinkela_wire_10166;
    wire new_Jinkela_wire_10471;
    wire new_Jinkela_wire_3343;
    wire new_Jinkela_wire_1353;
    wire new_Jinkela_wire_5669;
    wire new_Jinkela_wire_8993;
    wire new_Jinkela_wire_6476;
    wire new_Jinkela_wire_4776;
    wire new_Jinkela_wire_9381;
    wire new_Jinkela_wire_513;
    wire new_Jinkela_wire_6176;
    wire new_Jinkela_wire_8790;
    wire new_Jinkela_wire_3052;
    wire new_Jinkela_wire_5721;
    wire new_Jinkela_wire_6265;
    wire new_Jinkela_wire_52;
    wire new_Jinkela_wire_10291;
    wire new_Jinkela_wire_582;
    wire new_Jinkela_wire_2714;
    wire n_0382_;
    wire new_Jinkela_wire_58;
    wire new_Jinkela_wire_9225;
    wire new_Jinkela_wire_9184;
    wire new_Jinkela_wire_5060;
    wire new_Jinkela_wire_7994;
    wire new_Jinkela_wire_9663;
    wire new_net_2507;
    wire new_Jinkela_wire_4803;
    wire new_Jinkela_wire_9729;
    wire new_Jinkela_wire_4345;
    wire n_1076_;
    wire new_Jinkela_wire_5636;
    wire new_Jinkela_wire_5340;
    wire new_Jinkela_wire_7932;
    wire new_Jinkela_wire_4332;
    wire new_Jinkela_wire_8009;
    wire n_0716_;
    wire new_Jinkela_wire_4888;
    wire new_Jinkela_wire_3817;
    wire new_Jinkela_wire_10527;
    wire new_Jinkela_wire_4790;
    wire n_0625_;
    wire new_Jinkela_wire_3961;
    wire n_0449_;
    wire new_Jinkela_wire_4876;
    wire new_Jinkela_wire_6687;
    wire new_Jinkela_wire_252;
    wire new_Jinkela_wire_5610;
    wire new_Jinkela_wire_7250;
    wire new_Jinkela_wire_1592;
    wire new_Jinkela_wire_2315;
    wire new_Jinkela_wire_7274;
    wire new_Jinkela_wire_5409;
    wire new_Jinkela_wire_6067;
    wire new_Jinkela_wire_6402;
    wire new_Jinkela_wire_5656;
    wire new_Jinkela_wire_9134;
    wire new_Jinkela_wire_8236;
    wire new_Jinkela_wire_5810;
    wire new_Jinkela_wire_8597;
    wire new_Jinkela_wire_4656;
    wire n_1168_;
    wire new_Jinkela_wire_8361;
    wire new_Jinkela_wire_4342;
    wire new_Jinkela_wire_751;
    wire new_Jinkela_wire_7589;
    wire new_Jinkela_wire_10242;
    wire new_Jinkela_wire_8552;
    wire new_Jinkela_wire_466;
    wire new_Jinkela_wire_8294;
    wire new_Jinkela_wire_4223;
    wire new_Jinkela_wire_10222;
    wire new_Jinkela_wire_3171;
    wire new_Jinkela_wire_4859;
    wire new_Jinkela_wire_7370;
    wire n_0185_;
    wire new_Jinkela_wire_2380;
    wire new_Jinkela_wire_7549;
    wire n_0849_;
    wire new_Jinkela_wire_8927;
    wire new_Jinkela_wire_1451;
    wire new_Jinkela_wire_2216;
    wire new_Jinkela_wire_1319;
    wire new_Jinkela_wire_1007;
    wire new_Jinkela_wire_9610;
    wire new_Jinkela_wire_6961;
    wire n_0536_;
    wire new_Jinkela_wire_7309;
    wire new_Jinkela_wire_9231;
    wire new_Jinkela_wire_8017;
    wire n_0956_;
    wire new_Jinkela_wire_8028;
    wire new_Jinkela_wire_6495;
    wire new_Jinkela_wire_2889;
    wire new_Jinkela_wire_8139;
    wire new_Jinkela_wire_8207;
    wire new_Jinkela_wire_10530;
    wire new_Jinkela_wire_1905;
    wire new_Jinkela_wire_9426;
    wire new_Jinkela_wire_7285;
    wire n_0255_;
    wire new_Jinkela_wire_4551;
    wire new_Jinkela_wire_6739;
    wire new_Jinkela_wire_10233;
    wire new_Jinkela_wire_7214;
    wire new_Jinkela_wire_3919;
    wire new_Jinkela_wire_7469;
    wire new_Jinkela_wire_2371;
    wire new_Jinkela_wire_1287;
    wire new_Jinkela_wire_1048;
    wire new_Jinkela_wire_5556;
    wire n_1267_;
    wire new_Jinkela_wire_440;
    wire new_Jinkela_wire_7746;
    wire n_0772_;
    wire new_Jinkela_wire_7024;
    wire new_Jinkela_wire_7973;
    wire new_Jinkela_wire_8747;
    wire new_Jinkela_wire_5868;
    wire new_Jinkela_wire_4178;
    wire new_Jinkela_wire_4946;
    wire new_Jinkela_wire_9191;
    wire new_Jinkela_wire_6390;
    wire new_Jinkela_wire_5835;
    wire new_Jinkela_wire_568;
    wire new_Jinkela_wire_5231;
    wire new_net_2552;
    wire new_Jinkela_wire_1486;
    wire new_Jinkela_wire_8741;
    wire n_1116_;
    wire new_Jinkela_wire_1767;
    wire new_Jinkela_wire_2938;
    wire new_Jinkela_wire_3374;
    wire new_Jinkela_wire_6005;
    wire new_Jinkela_wire_5000;
    wire new_Jinkela_wire_8569;
    wire new_Jinkela_wire_4321;
    wire new_Jinkela_wire_6931;
    wire new_Jinkela_wire_7738;
    wire new_Jinkela_wire_2508;
    wire new_Jinkela_wire_6420;
    wire new_Jinkela_wire_10531;
    wire new_Jinkela_wire_2238;
    wire new_Jinkela_wire_10429;
    wire new_Jinkela_wire_6861;
    wire new_Jinkela_wire_8633;
    wire new_Jinkela_wire_6089;
    wire new_Jinkela_wire_8580;
    wire new_Jinkela_wire_6228;
    wire new_Jinkela_wire_6759;
    wire new_Jinkela_wire_8391;
    wire new_Jinkela_wire_2681;
    wire new_Jinkela_wire_10534;
    wire n_0101_;
    wire new_Jinkela_wire_60;
    wire new_Jinkela_wire_10370;
    wire new_Jinkela_wire_4458;
    wire new_Jinkela_wire_1082;
    wire new_Jinkela_wire_5987;
    wire new_Jinkela_wire_10018;
    wire new_Jinkela_wire_7688;
    wire new_Jinkela_wire_10381;
    wire new_Jinkela_wire_2895;
    wire new_Jinkela_wire_2348;
    wire new_Jinkela_wire_4351;
    wire new_Jinkela_wire_6272;
    wire new_Jinkela_wire_4710;
    wire new_Jinkela_wire_3114;
    wire new_Jinkela_wire_4280;
    wire new_Jinkela_wire_10350;
    wire new_Jinkela_wire_8202;
    wire new_Jinkela_wire_5567;
    wire new_Jinkela_wire_1516;
    wire new_Jinkela_wire_4923;
    wire new_Jinkela_wire_10470;
    wire new_Jinkela_wire_5071;
    wire new_Jinkela_wire_6887;
    wire new_Jinkela_wire_6847;
    wire n_1154_;
    wire n_0051_;
    wire new_Jinkela_wire_9384;
    wire new_Jinkela_wire_5016;
    wire new_Jinkela_wire_5983;
    wire new_Jinkela_wire_5690;
    wire new_Jinkela_wire_4928;
    wire new_Jinkela_wire_6100;
    wire new_Jinkela_wire_267;
    wire new_Jinkela_wire_9728;
    wire new_Jinkela_wire_9454;
    wire new_Jinkela_wire_770;
    wire n_0672_;
    wire new_Jinkela_wire_3490;
    wire n_0172_;
    wire new_Jinkela_wire_4750;
    wire new_Jinkela_wire_6178;
    wire new_Jinkela_wire_1099;
    wire new_Jinkela_wire_31;
    wire new_Jinkela_wire_3013;
    wire n_1054_;
    wire new_Jinkela_wire_517;
    wire n_0110_;
    wire n_0293_;
    wire new_Jinkela_wire_6898;
    wire new_Jinkela_wire_1163;
    wire new_Jinkela_wire_4050;
    wire new_Jinkela_wire_8594;
    wire new_Jinkela_wire_10424;
    wire new_Jinkela_wire_3041;
    wire new_Jinkela_wire_3282;
    wire new_Jinkela_wire_2557;
    wire new_Jinkela_wire_10024;
    wire new_Jinkela_wire_8447;
    wire new_Jinkela_wire_4532;
    wire new_Jinkela_wire_5260;
    wire new_Jinkela_wire_282;
    wire new_Jinkela_wire_4449;
    wire new_Jinkela_wire_1835;
    wire new_Jinkela_wire_1338;
    wire new_Jinkela_wire_7785;
    wire new_Jinkela_wire_5328;
    wire new_Jinkela_wire_3711;
    wire new_Jinkela_wire_9027;
    wire new_Jinkela_wire_1892;
    wire new_Jinkela_wire_6015;
    wire new_Jinkela_wire_5345;
    wire new_Jinkela_wire_6952;
    wire new_Jinkela_wire_4304;
    wire new_Jinkela_wire_8550;
    wire new_Jinkela_wire_1535;
    wire new_Jinkela_wire_1427;
    wire new_Jinkela_wire_1166;
    wire new_Jinkela_wire_1069;
    wire new_Jinkela_wire_6018;
    wire new_Jinkela_wire_9851;
    wire new_Jinkela_wire_6204;
    wire new_Jinkela_wire_478;
    wire new_Jinkela_wire_3870;
    wire new_Jinkela_wire_7647;
    wire new_Jinkela_wire_5279;
    wire new_Jinkela_wire_8291;
    wire new_Jinkela_wire_4882;
    wire new_Jinkela_wire_9022;
    wire new_Jinkela_wire_6844;
    wire new_Jinkela_wire_5848;
    wire new_Jinkela_wire_2396;
    wire new_Jinkela_wire_7386;
    wire new_Jinkela_wire_10197;
    wire new_Jinkela_wire_9676;
    wire new_net_2556;
    wire new_Jinkela_wire_335;
    wire new_Jinkela_wire_5303;
    wire new_Jinkela_wire_2519;
    wire new_Jinkela_wire_5403;
    wire new_Jinkela_wire_3304;
    wire new_Jinkela_wire_8689;
    wire new_Jinkela_wire_3627;
    wire new_Jinkela_wire_4181;
    wire n_0521_;
    wire new_net_2521;
    wire new_Jinkela_wire_214;
    wire new_Jinkela_wire_1148;
    wire new_Jinkela_wire_849;
    wire n_0003_;
    wire n_1308_;
    wire new_Jinkela_wire_8706;
    wire new_Jinkela_wire_3071;
    wire new_Jinkela_wire_3157;
    wire new_Jinkela_wire_1130;
    wire new_Jinkela_wire_7859;
    wire new_Jinkela_wire_6814;
    wire new_Jinkela_wire_5616;
    wire new_Jinkela_wire_8943;
    wire new_Jinkela_wire_4844;
    wire new_Jinkela_wire_8928;
    wire new_Jinkela_wire_1472;
    wire new_Jinkela_wire_8248;
    wire new_Jinkela_wire_7268;
    wire n_1120_;
    wire n_0793_;
    wire n_0216_;
    wire new_Jinkela_wire_3614;
    wire new_Jinkela_wire_2137;
    wire new_Jinkela_wire_973;
    wire n_0759_;
    wire new_Jinkela_wire_154;
    wire new_Jinkela_wire_10122;
    wire new_Jinkela_wire_10617;
    wire new_Jinkela_wire_3115;
    wire new_Jinkela_wire_7355;
    wire new_Jinkela_wire_3274;
    wire new_Jinkela_wire_7441;
    wire new_Jinkela_wire_2582;
    wire new_Jinkela_wire_3126;
    wire new_Jinkela_wire_1891;
    wire new_Jinkela_wire_7780;
    wire new_Jinkela_wire_2667;
    wire n_0151_;
    wire new_Jinkela_wire_7167;
    wire new_Jinkela_wire_4337;
    wire new_Jinkela_wire_8173;
    wire new_Jinkela_wire_7591;
    wire new_Jinkela_wire_7881;
    wire new_Jinkela_wire_1279;
    wire new_Jinkela_wire_7692;
    wire new_Jinkela_wire_5373;
    wire new_Jinkela_wire_2467;
    wire n_0169_;
    wire new_Jinkela_wire_7878;
    wire new_Jinkela_wire_2021;
    wire new_Jinkela_wire_2659;
    wire new_Jinkela_wire_4640;
    wire new_Jinkela_wire_9222;
    wire new_net_2549;
    wire n_0164_;
    wire n_0136_;
    wire new_Jinkela_wire_3354;
    wire new_Jinkela_wire_1794;
    wire new_Jinkela_wire_2564;
    wire new_Jinkela_wire_4339;
    wire n_0969_;
    wire new_Jinkela_wire_7953;
    wire new_Jinkela_wire_3848;
    wire new_Jinkela_wire_6613;
    wire new_Jinkela_wire_7406;
    wire new_Jinkela_wire_9633;
    wire n_0072_;
    wire new_Jinkela_wire_4769;
    wire new_Jinkela_wire_5589;
    wire new_Jinkela_wire_1641;
    wire new_Jinkela_wire_8227;
    wire new_Jinkela_wire_1337;
    wire new_Jinkela_wire_6337;
    wire n_1217_;
    wire new_Jinkela_wire_8617;
    wire new_Jinkela_wire_4451;
    wire new_Jinkela_wire_417;
    wire new_Jinkela_wire_5164;
    wire new_Jinkela_wire_5383;
    wire new_Jinkela_wire_9548;
    wire new_Jinkela_wire_5886;
    wire new_Jinkela_wire_5996;
    wire new_Jinkela_wire_4400;
    wire new_Jinkela_wire_9502;
    wire new_Jinkela_wire_7788;
    wire new_Jinkela_wire_862;
    wire new_Jinkela_wire_4686;
    wire new_Jinkela_wire_4545;
    wire n_1335_;
    wire new_Jinkela_wire_1326;
    wire new_Jinkela_wire_1264;
    wire new_Jinkela_wire_6122;
    wire new_Jinkela_wire_8312;
    wire new_Jinkela_wire_9657;
    wire new_Jinkela_wire_2274;
    wire new_Jinkela_wire_4405;
    wire n_0031_;
    wire new_Jinkela_wire_8801;
    wire new_Jinkela_wire_1276;
    wire new_Jinkela_wire_7837;
    wire new_Jinkela_wire_1138;
    wire new_Jinkela_wire_7058;
    wire new_Jinkela_wire_1679;
    wire new_Jinkela_wire_9596;
    wire new_Jinkela_wire_5766;
    wire new_Jinkela_wire_2081;
    wire new_Jinkela_wire_1387;
    wire new_Jinkela_wire_7867;
    wire new_Jinkela_wire_10632;
    wire new_Jinkela_wire_926;
    wire new_Jinkela_wire_272;
    wire new_Jinkela_wire_8208;
    wire new_Jinkela_wire_5116;
    wire new_net_2570;
    wire new_Jinkela_wire_7116;
    wire new_Jinkela_wire_9409;
    wire new_Jinkela_wire_441;
    wire new_Jinkela_wire_1847;
    wire new_Jinkela_wire_2308;
    wire new_Jinkela_wire_6497;
    wire new_Jinkela_wire_1289;
    wire new_Jinkela_wire_10347;
    wire new_Jinkela_wire_9675;
    wire new_Jinkela_wire_9397;
    wire new_Jinkela_wire_2418;
    wire n_0147_;
    wire new_Jinkela_wire_8732;
    wire new_Jinkela_wire_5332;
    wire new_Jinkela_wire_4514;
    wire n_0430_;
    wire new_Jinkela_wire_4284;
    wire new_Jinkela_wire_6226;
    wire new_Jinkela_wire_5713;
    wire new_Jinkela_wire_6855;
    wire new_Jinkela_wire_7791;
    wire new_Jinkela_wire_3519;
    wire new_Jinkela_wire_2614;
    wire new_Jinkela_wire_8158;
    wire new_Jinkela_wire_8075;
    wire new_Jinkela_wire_2507;
    wire new_Jinkela_wire_1308;
    wire new_Jinkela_wire_10389;
    wire new_Jinkela_wire_7224;
    wire new_Jinkela_wire_256;
    wire new_Jinkela_wire_5237;
    wire new_Jinkela_wire_4482;
    wire new_Jinkela_wire_10473;
    wire new_Jinkela_wire_5228;
    wire new_Jinkela_wire_1531;
    wire new_Jinkela_wire_5498;
    wire new_Jinkela_wire_1789;
    wire new_Jinkela_wire_8892;
    wire new_Jinkela_wire_295;
    wire new_Jinkela_wire_1841;
    wire new_Jinkela_wire_3324;
    wire new_Jinkela_wire_1844;
    wire new_Jinkela_wire_3080;
    wire new_Jinkela_wire_6634;
    wire new_Jinkela_wire_347;
    wire new_Jinkela_wire_9431;
    wire new_Jinkela_wire_7605;
    wire new_Jinkela_wire_8189;
    wire new_Jinkela_wire_10196;
    wire new_Jinkela_wire_1518;
    wire new_Jinkela_wire_6576;
    wire new_Jinkela_wire_8307;
    wire new_Jinkela_wire_1826;
    wire new_Jinkela_wire_8456;
    wire new_Jinkela_wire_4639;
    wire new_Jinkela_wire_4085;
    wire new_Jinkela_wire_3814;
    wire new_Jinkela_wire_9656;
    wire new_Jinkela_wire_2269;
    wire new_Jinkela_wire_9621;
    wire n_0634_;
    wire new_Jinkela_wire_3193;
    wire new_Jinkela_wire_7587;
    wire new_Jinkela_wire_4341;
    wire n_1108_;
    wire new_Jinkela_wire_156;
    wire new_Jinkela_wire_8342;
    wire new_Jinkela_wire_3063;
    wire new_Jinkela_wire_1364;
    wire new_Jinkela_wire_6328;
    wire new_Jinkela_wire_8198;
    wire new_Jinkela_wire_202;
    wire new_Jinkela_wire_3134;
    wire new_Jinkela_wire_8040;
    wire new_Jinkela_wire_5486;
    wire new_Jinkela_wire_9693;
    wire new_Jinkela_wire_3378;
    wire new_Jinkela_wire_8004;
    wire new_Jinkela_wire_10133;
    wire new_Jinkela_wire_8720;
    wire new_Jinkela_wire_3638;
    wire new_Jinkela_wire_5259;
    wire new_Jinkela_wire_8636;
    wire new_Jinkela_wire_1949;
    wire new_Jinkela_wire_2573;
    wire n_0734_;
    wire new_Jinkela_wire_345;
    wire new_Jinkela_wire_10025;
    wire new_Jinkela_wire_7622;
    wire new_Jinkela_wire_9428;
    wire new_Jinkela_wire_7625;
    wire new_Jinkela_wire_5314;
    wire new_Jinkela_wire_9259;
    wire new_Jinkela_wire_1064;
    wire new_Jinkela_wire_9419;
    wire new_Jinkela_wire_10489;
    wire new_Jinkela_wire_5678;
    wire new_Jinkela_wire_8955;
    wire new_Jinkela_wire_2271;
    wire new_Jinkela_wire_8614;
    wire n_1211_;
    wire n_0690_;
    wire new_Jinkela_wire_127;
    wire new_Jinkela_wire_8224;
    wire new_Jinkela_wire_488;
    wire new_Jinkela_wire_8757;
    wire new_Jinkela_wire_5869;
    wire new_Jinkela_wire_4338;
    wire new_Jinkela_wire_6883;
    wire new_Jinkela_wire_3360;
    wire new_Jinkela_wire_3678;
    wire new_Jinkela_wire_8484;
    wire n_0664_;
    wire new_Jinkela_wire_6245;
    wire new_Jinkela_wire_410;
    wire new_Jinkela_wire_1001;
    wire new_Jinkela_wire_2005;
    wire new_Jinkela_wire_2082;
    wire n_1030_;
    wire new_Jinkela_wire_9743;
    wire new_Jinkela_wire_815;
    wire new_Jinkela_wire_507;
    wire new_Jinkela_wire_8389;
    wire new_Jinkela_wire_2786;
    wire new_Jinkela_wire_8157;
    wire new_Jinkela_wire_1342;
    wire new_Jinkela_wire_3634;
    wire new_Jinkela_wire_6121;
    wire new_Jinkela_wire_8014;
    wire new_Jinkela_wire_9804;
    wire new_Jinkela_wire_1256;
    wire new_Jinkela_wire_2937;
    wire new_Jinkela_wire_376;
    wire new_Jinkela_wire_2827;
    wire n_0677_;
    wire new_Jinkela_wire_6881;
    wire n_0886_;
    wire new_Jinkela_wire_2357;
    wire new_Jinkela_wire_4980;
    wire new_Jinkela_wire_3799;
    wire new_Jinkela_wire_9348;
    wire n_1014_;
    wire new_Jinkela_wire_6445;
    wire new_Jinkela_wire_10372;
    wire new_Jinkela_wire_7698;
    wire new_Jinkela_wire_4412;
    wire new_Jinkela_wire_10299;
    wire new_Jinkela_wire_9792;
    wire n_0002_;
    wire new_Jinkela_wire_2902;
    wire new_Jinkela_wire_4972;
    wire new_Jinkela_wire_7075;
    wire new_Jinkela_wire_5630;
    wire new_Jinkela_wire_8898;
    wire n_0270_;
    wire n_0769_;
    wire new_Jinkela_wire_7461;
    wire new_Jinkela_wire_10391;
    wire new_Jinkela_wire_7880;
    wire new_Jinkela_wire_5182;
    wire new_Jinkela_wire_1269;
    wire new_Jinkela_wire_6796;
    wire new_Jinkela_wire_8650;
    wire new_Jinkela_wire_7025;
    wire new_Jinkela_wire_7730;
    wire new_Jinkela_wire_5376;
    wire n_1162_;
    wire new_Jinkela_wire_1384;
    wire new_Jinkela_wire_7939;
    wire new_Jinkela_wire_8427;
    wire new_Jinkela_wire_7886;
    wire new_Jinkela_wire_9855;
    wire new_Jinkela_wire_2572;
    wire new_Jinkela_wire_616;
    wire n_0074_;
    wire new_Jinkela_wire_1162;
    wire new_Jinkela_wire_3166;
    wire n_0442_;
    wire new_Jinkela_wire_2546;
    wire new_Jinkela_wire_1643;
    wire new_Jinkela_wire_7382;
    wire new_Jinkela_wire_575;
    wire new_Jinkela_wire_5939;
    wire n_0868_;
    wire n_1195_;
    wire new_Jinkela_wire_5674;
    wire new_Jinkela_wire_6765;
    wire new_Jinkela_wire_2491;
    wire new_Jinkela_wire_7844;
    wire new_Jinkela_wire_6361;
    wire new_Jinkela_wire_2086;
    wire new_Jinkela_wire_9821;
    wire new_Jinkela_wire_3168;
    wire new_Jinkela_wire_9567;
    wire new_Jinkela_wire_4697;
    wire new_Jinkela_wire_1529;
    wire new_Jinkela_wire_3894;
    wire new_Jinkela_wire_4183;
    wire new_Jinkela_wire_10387;
    wire new_Jinkela_wire_6316;
    wire new_Jinkela_wire_6186;
    wire n_0053_;
    wire new_Jinkela_wire_9004;
    wire new_Jinkela_wire_3570;
    wire new_Jinkela_wire_4791;
    wire new_Jinkela_wire_8820;
    wire new_Jinkela_wire_3412;
    wire new_Jinkela_wire_2923;
    wire n_0809_;
    wire new_Jinkela_wire_4895;
    wire new_Jinkela_wire_10147;
    wire new_Jinkela_wire_3939;
    wire new_Jinkela_wire_8402;
    wire new_Jinkela_wire_5039;
    wire new_Jinkela_wire_542;
    wire new_Jinkela_wire_9394;
    wire new_Jinkela_wire_2362;
    wire new_Jinkela_wire_3699;
    wire new_Jinkela_wire_9943;
    wire new_Jinkela_wire_10264;
    wire new_Jinkela_wire_864;
    wire new_Jinkela_wire_6130;
    wire n_0488_;
    wire new_Jinkela_wire_5074;
    wire new_Jinkela_wire_9018;
    wire new_Jinkela_wire_3503;
    wire new_Jinkela_wire_2809;
    wire new_Jinkela_wire_1630;
    wire new_Jinkela_wire_8289;
    wire new_Jinkela_wire_2691;
    wire new_Jinkela_wire_10143;
    wire new_Jinkela_wire_7227;
    wire new_Jinkela_wire_9577;
    wire new_Jinkela_wire_907;
    wire new_Jinkela_wire_1517;
    wire new_Jinkela_wire_2854;
    wire new_Jinkela_wire_4592;
    wire new_Jinkela_wire_1104;
    wire new_Jinkela_wire_4861;
    wire new_Jinkela_wire_6358;
    wire n_0244_;
    wire new_Jinkela_wire_35;
    wire new_Jinkela_wire_6478;
    wire new_Jinkela_wire_340;
    wire new_Jinkela_wire_10039;
    wire new_Jinkela_wire_7849;
    wire new_Jinkela_wire_2830;
    wire new_Jinkela_wire_2048;
    wire new_Jinkela_wire_6817;
    wire new_net_2539;
    wire new_Jinkela_wire_8968;
    wire new_Jinkela_wire_3889;
    wire new_Jinkela_wire_6732;
    wire new_Jinkela_wire_1546;
    wire new_Jinkela_wire_6507;
    wire new_Jinkela_wire_8354;
    wire new_Jinkela_wire_9131;
    wire new_Jinkela_wire_5534;
    wire new_Jinkela_wire_5582;
    wire new_Jinkela_wire_4816;
    wire new_Jinkela_wire_6001;
    wire new_Jinkela_wire_6208;
    wire new_Jinkela_wire_185;
    wire n_0165_;
    wire n_1099_;
    wire n_0627_;
    wire new_Jinkela_wire_6491;
    wire new_Jinkela_wire_3059;
    wire new_Jinkela_wire_6368;
    wire new_Jinkela_wire_2087;
    wire new_Jinkela_wire_3980;
    wire new_Jinkela_wire_7751;
    wire n_0256_;
    wire new_Jinkela_wire_988;
    wire n_0805_;
    wire n_0208_;
    wire new_Jinkela_wire_10061;
    wire new_Jinkela_wire_2497;
    wire new_Jinkela_wire_3685;
    wire new_Jinkela_wire_5245;
    wire new_Jinkela_wire_8265;
    wire new_Jinkela_wire_7826;
    wire new_Jinkela_wire_7623;
    wire new_Jinkela_wire_2593;
    wire n_1343_;
    wire new_Jinkela_wire_611;
    wire new_Jinkela_wire_1327;
    wire new_Jinkela_wire_595;
    wire new_Jinkela_wire_8953;
    wire new_Jinkela_wire_760;
    wire new_Jinkela_wire_5944;
    wire new_Jinkela_wire_3393;
    wire new_Jinkela_wire_10415;
    wire n_0248_;
    wire new_Jinkela_wire_1871;
    wire new_Jinkela_wire_2217;
    wire new_Jinkela_wire_6224;
    wire new_Jinkela_wire_495;
    wire n_0532_;
    wire new_Jinkela_wire_2712;
    wire new_Jinkela_wire_9903;
    wire new_Jinkela_wire_7475;
    wire n_0851_;
    wire new_Jinkela_wire_1766;
    wire new_Jinkela_wire_7061;
    wire new_Jinkela_wire_1501;
    wire new_Jinkela_wire_10235;
    wire new_Jinkela_wire_8949;
    wire new_Jinkela_wire_7944;
    wire new_Jinkela_wire_5997;
    wire new_Jinkela_wire_4655;
    wire n_0434_;
    wire n_1020_;
    wire n_1170_;
    wire new_Jinkela_wire_9664;
    wire new_Jinkela_wire_73;
    wire new_Jinkela_wire_4298;
    wire new_Jinkela_wire_4560;
    wire new_Jinkela_wire_10430;
    wire new_Jinkela_wire_10105;
    wire n_0714_;
    wire new_Jinkela_wire_9563;
    wire n_1087_;
    wire new_Jinkela_wire_294;
    wire new_Jinkela_wire_5031;
    wire n_0636_;
    wire new_Jinkela_wire_7882;
    wire new_Jinkela_wire_1722;
    wire new_Jinkela_wire_4425;
    wire new_Jinkela_wire_10453;
    wire new_Jinkela_wire_10474;
    wire n_0710_;
    wire new_Jinkela_wire_5925;
    wire new_Jinkela_wire_1361;
    wire new_Jinkela_wire_9847;
    wire new_Jinkela_wire_7829;
    wire new_Jinkela_wire_6598;
    wire new_Jinkela_wire_9472;
    wire new_Jinkela_wire_1129;
    wire new_Jinkela_wire_4077;
    wire new_Jinkela_wire_4492;
    wire n_0660_;
    wire new_Jinkela_wire_2267;
    wire new_Jinkela_wire_3070;
    wire new_Jinkela_wire_6493;
    wire new_Jinkela_wire_5833;
    wire new_Jinkela_wire_493;
    wire new_Jinkela_wire_9775;
    wire new_Jinkela_wire_10352;
    wire new_Jinkela_wire_4645;
    wire new_Jinkela_wire_3048;
    wire new_Jinkela_wire_8547;
    wire new_Jinkela_wire_1025;
    wire new_Jinkela_wire_6951;
    wire new_Jinkela_wire_9601;
    wire new_Jinkela_wire_6064;
    wire new_Jinkela_wire_1213;
    wire new_Jinkela_wire_3681;
    wire new_Jinkela_wire_8600;
    wire new_Jinkela_wire_456;
    wire new_Jinkela_wire_612;
    wire new_Jinkela_wire_8201;
    wire new_Jinkela_wire_7875;
    wire new_Jinkela_wire_828;
    wire new_Jinkela_wire_9211;
    wire new_Jinkela_wire_8015;
    wire new_Jinkela_wire_4875;
    wire new_Jinkela_wire_4331;
    wire new_Jinkela_wire_5538;
    wire new_Jinkela_wire_3488;
    wire new_Jinkela_wire_9770;
    wire new_Jinkela_wire_5931;
    wire n_0715_;
    wire new_Jinkela_wire_5491;
    wire new_Jinkela_wire_7926;
    wire n_1210_;
    wire new_Jinkela_wire_68;
    wire new_Jinkela_wire_6591;
    wire n_0937_;
    wire n_0345_;
    wire new_Jinkela_wire_5059;
    wire new_Jinkela_wire_8555;
    wire new_Jinkela_wire_1492;
    wire new_Jinkela_wire_1672;
    wire new_Jinkela_wire_3199;
    wire new_Jinkela_wire_8068;
    wire new_Jinkela_wire_2768;
    wire new_Jinkela_wire_2419;
    wire new_Jinkela_wire_3481;
    wire n_0544_;
    wire new_Jinkela_wire_9392;
    wire new_Jinkela_wire_4049;
    wire new_Jinkela_wire_5356;
    wire new_Jinkela_wire_6501;
    wire new_Jinkela_wire_3062;
    wire new_Jinkela_wire_39;
    wire new_Jinkela_wire_8404;
    wire new_Jinkela_wire_7101;
    wire new_Jinkela_wire_6771;
    wire n_0592_;
    wire new_Jinkela_wire_7371;
    wire new_Jinkela_wire_3643;
    wire n_0168_;
    wire new_Jinkela_wire_9326;
    wire new_Jinkela_wire_6585;
    wire new_Jinkela_wire_9034;
    wire new_net_2568;
    wire new_Jinkela_wire_730;
    wire new_Jinkela_wire_1440;
    wire new_Jinkela_wire_4526;
    wire new_Jinkela_wire_5805;
    wire new_Jinkela_wire_7235;
    wire n_0852_;
    wire n_1362_;
    wire new_Jinkela_wire_2656;
    wire new_Jinkela_wire_4673;
    wire n_0134_;
    wire new_Jinkela_wire_856;
    wire new_Jinkela_wire_8537;
    wire new_Jinkela_wire_1733;
    wire new_Jinkela_wire_2683;
    wire new_Jinkela_wire_2734;
    wire new_Jinkela_wire_9061;
    wire new_Jinkela_wire_5381;
    wire new_Jinkela_wire_1685;
    wire new_Jinkela_wire_1182;
    wire new_Jinkela_wire_5122;
    wire new_Jinkela_wire_3066;
    wire new_Jinkela_wire_3504;
    wire n_0653_;
    wire new_Jinkela_wire_1126;
    wire new_Jinkela_wire_2727;
    wire new_Jinkela_wire_28;
    wire new_Jinkela_wire_5859;
    wire new_Jinkela_wire_505;
    wire new_Jinkela_wire_1600;
    wire new_Jinkela_wire_8907;
    wire n_0404_;
    wire new_Jinkela_wire_7466;
    wire new_Jinkela_wire_5729;
    wire new_Jinkela_wire_7565;
    wire new_Jinkela_wire_786;
    wire new_Jinkela_wire_1165;
    wire new_Jinkela_wire_5357;
    wire new_Jinkela_wire_2883;
    wire new_Jinkela_wire_4747;
    wire new_Jinkela_wire_4196;
    wire new_Jinkela_wire_2535;
    wire new_net_2533;
    wire new_Jinkela_wire_4210;
    wire new_Jinkela_wire_8713;
    wire new_Jinkela_wire_1810;
    wire new_Jinkela_wire_233;
    wire new_Jinkela_wire_6560;
    wire new_Jinkela_wire_9192;
    wire new_Jinkela_wire_10425;
    wire new_Jinkela_wire_5919;
    wire new_Jinkela_wire_1422;
    wire new_Jinkela_wire_10206;
    wire new_Jinkela_wire_9173;
    wire new_Jinkela_wire_2682;
    wire new_Jinkela_wire_6161;
    wire new_Jinkela_wire_2285;
    wire n_0220_;
    wire new_Jinkela_wire_8034;
    wire new_Jinkela_wire_3765;
    wire new_Jinkela_wire_8134;
    wire new_Jinkela_wire_6215;
    wire new_Jinkela_wire_3867;
    wire new_Jinkela_wire_268;
    wire new_Jinkela_wire_9788;
    wire new_Jinkela_wire_9522;
    wire new_Jinkela_wire_3117;
    wire new_Jinkela_wire_3263;
    wire n_0323_;
    wire new_Jinkela_wire_3260;
    wire new_Jinkela_wire_8733;
    wire new_Jinkela_wire_3538;
    wire new_Jinkela_wire_9212;
    wire new_Jinkela_wire_1723;
    wire n_1283_;
    wire new_Jinkela_wire_5949;
    wire new_Jinkela_wire_10456;
    wire new_Jinkela_wire_2004;
    wire new_net_7;
    wire new_Jinkela_wire_2028;
    wire n_0166_;
    wire new_Jinkela_wire_4318;
    wire new_Jinkela_wire_6389;
    wire new_Jinkela_wire_8147;
    wire new_Jinkela_wire_2788;
    wire new_Jinkela_wire_10006;
    wire new_Jinkela_wire_3908;
    wire new_Jinkela_wire_725;
    wire new_Jinkela_wire_1055;
    wire new_Jinkela_wire_3129;
    wire n_0645_;
    wire new_Jinkela_wire_3559;
    wire new_Jinkela_wire_9509;
    wire new_Jinkela_wire_6210;
    wire n_1248_;
    wire new_Jinkela_wire_4881;
    wire new_Jinkela_wire_7422;
    wire n_1007_;
    wire new_Jinkela_wire_9250;
    wire new_Jinkela_wire_8025;
    wire new_Jinkela_wire_1553;
    wire n_0739_;
    wire new_Jinkela_wire_7502;
    wire new_Jinkela_wire_4792;
    wire new_Jinkela_wire_9640;
    wire n_0298_;
    wire new_Jinkela_wire_5462;
    wire new_Jinkela_wire_2549;
    wire n_0207_;
    wire new_Jinkela_wire_6088;
    wire new_Jinkela_wire_9535;
    wire new_Jinkela_wire_5269;
    wire new_Jinkela_wire_533;
    wire new_Jinkela_wire_2811;
    wire new_Jinkela_wire_475;
    wire new_Jinkela_wire_118;
    wire new_Jinkela_wire_5485;
    wire n_0321_;
    wire new_Jinkela_wire_7868;
    wire new_Jinkela_wire_5369;
    wire n_0479_;
    wire new_Jinkela_wire_3061;
    wire new_Jinkela_wire_9968;
    wire new_Jinkela_wire_10433;
    wire new_Jinkela_wire_9726;
    wire n_0891_;
    wire new_Jinkela_wire_7985;
    wire new_Jinkela_wire_4534;
    wire n_0122_;
    wire new_Jinkela_wire_5495;
    wire n_0910_;
    wire new_Jinkela_wire_3897;
    wire n_1160_;
    wire new_Jinkela_wire_1539;
    wire new_Jinkela_wire_2783;
    wire new_Jinkela_wire_3127;
    wire new_Jinkela_wire_5440;
    wire new_Jinkela_wire_5734;
    wire new_Jinkela_wire_640;
    wire new_Jinkela_wire_8290;
    wire new_Jinkela_wire_2637;
    wire new_Jinkela_wire_7267;
    wire new_Jinkela_wire_638;
    wire new_Jinkela_wire_1137;
    wire new_Jinkela_wire_834;
    wire new_Jinkela_wire_10395;
    wire new_Jinkela_wire_2731;
    wire new_Jinkela_wire_9400;
    wire new_Jinkela_wire_2205;
    wire n_0079_;
    wire new_Jinkela_wire_10529;
    wire new_Jinkela_wire_9447;
    wire new_Jinkela_wire_1779;
    wire new_Jinkela_wire_10344;
    wire new_Jinkela_wire_9562;
    wire new_Jinkela_wire_581;
    wire new_Jinkela_wire_7470;
    wire new_Jinkela_wire_9456;
    wire new_Jinkela_wire_6195;
    wire new_Jinkela_wire_5221;
    wire n_0401_;
    wire new_Jinkela_wire_4681;
    wire new_Jinkela_wire_4027;
    wire new_Jinkela_wire_5984;
    wire n_1366_;
    wire n_0980_;
    wire new_Jinkela_wire_4741;
    wire new_Jinkela_wire_4982;
    wire new_Jinkela_wire_1931;
    wire n_0490_;
    wire new_Jinkela_wire_776;
    wire new_Jinkela_wire_8296;
    wire new_Jinkela_wire_2926;
    wire new_Jinkela_wire_3101;
    wire new_Jinkela_wire_5879;
    wire new_Jinkela_wire_2531;
    wire n_1202_;
    wire new_Jinkela_wire_1409;
    wire new_Jinkela_wire_3449;
    wire n_0183_;
    wire new_Jinkela_wire_4348;
    wire n_1141_;
    wire new_Jinkela_wire_6308;
    wire new_Jinkela_wire_7066;
    wire new_Jinkela_wire_5932;
    wire new_Jinkela_wire_1584;
    wire new_Jinkela_wire_7053;
    wire new_Jinkela_wire_2796;
    wire new_Jinkela_wire_7773;
    wire new_Jinkela_wire_3722;
    wire new_Jinkela_wire_153;
    wire new_Jinkela_wire_2076;
    wire new_Jinkela_wire_2638;
    wire new_Jinkela_wire_8629;
    wire new_Jinkela_wire_9606;
    wire new_Jinkela_wire_1291;
    wire new_Jinkela_wire_1301;
    wire new_Jinkela_wire_7839;
    wire new_Jinkela_wire_2584;
    wire new_Jinkela_wire_5484;
    wire new_Jinkela_wire_9204;
    wire new_Jinkela_wire_1740;
    wire new_Jinkela_wire_1748;
    wire new_Jinkela_wire_4579;
    wire new_Jinkela_wire_10091;
    wire new_Jinkela_wire_7269;
    wire n_0178_;
    wire new_Jinkela_wire_4584;
    wire new_Jinkela_wire_7427;
    wire new_Jinkela_wire_9013;
    wire new_Jinkela_wire_9979;
    wire new_Jinkela_wire_7389;
    wire new_Jinkela_wire_10581;
    wire new_Jinkela_wire_3455;
    wire new_Jinkela_wire_2686;
    wire new_Jinkela_wire_164;
    wire new_Jinkela_wire_7750;
    wire new_Jinkela_wire_2627;
    wire new_Jinkela_wire_5989;
    wire new_Jinkela_wire_9479;
    wire new_Jinkela_wire_7000;
    wire new_Jinkela_wire_655;
    wire new_Jinkela_wire_5814;
    wire new_Jinkela_wire_688;
    wire new_Jinkela_wire_9436;
    wire new_Jinkela_wire_6307;
    wire new_Jinkela_wire_1400;
    wire new_Jinkela_wire_3081;
    wire new_Jinkela_wire_9824;
    wire new_Jinkela_wire_6471;
    wire new_Jinkela_wire_1283;
    wire new_Jinkela_wire_10288;
    wire new_Jinkela_wire_1664;
    wire new_Jinkela_wire_3992;
    wire new_Jinkela_wire_9430;
    wire new_net_2541;
    wire new_Jinkela_wire_7572;
    wire new_Jinkela_wire_1846;
    wire new_Jinkela_wire_9975;
    wire new_Jinkela_wire_3745;
    wire new_Jinkela_wire_2599;
    wire new_Jinkela_wire_5701;
    wire n_0621_;
    wire n_0747_;
    wire new_Jinkela_wire_414;
    wire new_Jinkela_wire_3936;
    wire new_Jinkela_wire_3487;
    wire new_Jinkela_wire_1482;
    wire new_Jinkela_wire_3740;
    wire new_Jinkela_wire_3191;
    wire new_Jinkela_wire_1926;
    wire new_Jinkela_wire_2581;
    wire new_Jinkela_wire_5197;
    wire new_Jinkela_wire_7176;
    wire new_Jinkela_wire_10062;
    wire new_Jinkela_wire_8844;
    wire new_Jinkela_wire_7522;
    wire new_Jinkela_wire_3209;
    wire new_Jinkela_wire_6779;
    wire new_Jinkela_wire_5930;
    wire new_Jinkela_wire_8120;
    wire new_Jinkela_wire_4509;
    wire new_Jinkela_wire_603;
    wire new_Jinkela_wire_1498;
    wire new_Jinkela_wire_1729;
    wire n_0730_;
    wire n_0945_;
    wire new_Jinkela_wire_6238;
    wire n_0599_;
    wire new_Jinkela_wire_5173;
    wire new_Jinkela_wire_6022;
    wire new_Jinkela_wire_6090;
    wire new_Jinkela_wire_6275;
    wire n_1233_;
    wire new_Jinkela_wire_8655;
    wire new_Jinkela_wire_3533;
    wire new_Jinkela_wire_9097;
    wire new_Jinkela_wire_1234;
    wire new_Jinkela_wire_6336;
    wire new_Jinkela_wire_4575;
    wire new_Jinkela_wire_10257;
    wire new_Jinkela_wire_3812;
    wire new_Jinkela_wire_2161;
    wire new_Jinkela_wire_3054;
    wire new_Jinkela_wire_5489;
    wire new_Jinkela_wire_3073;
    wire new_Jinkela_wire_8637;
    wire new_Jinkela_wire_5514;
    wire n_0893_;
    wire new_Jinkela_wire_1690;
    wire new_Jinkela_wire_6260;
    wire new_Jinkela_wire_5952;
    wire new_Jinkela_wire_10604;
    wire new_Jinkela_wire_2943;
    wire new_Jinkela_wire_5133;
    wire new_Jinkela_wire_9012;
    wire new_Jinkela_wire_10001;
    wire new_Jinkela_wire_7351;
    wire new_Jinkela_wire_1739;
    wire new_Jinkela_wire_1322;
    wire new_Jinkela_wire_1278;
    wire new_Jinkela_wire_3181;
    wire new_Jinkela_wire_4032;
    wire new_Jinkela_wire_8863;
    wire new_Jinkela_wire_4688;
    wire new_Jinkela_wire_7109;
    wire new_Jinkela_wire_1822;
    wire new_Jinkela_wire_277;
    wire n_0411_;
    wire new_Jinkela_wire_1985;
    wire n_0399_;
    wire new_Jinkela_wire_3509;
    wire new_Jinkela_wire_512;
    wire new_Jinkela_wire_9674;
    wire new_Jinkela_wire_726;
    wire new_Jinkela_wire_9446;
    wire new_Jinkela_wire_5043;
    wire new_Jinkela_wire_4281;
    wire new_Jinkela_wire_4568;
    wire new_Jinkela_wire_210;
    wire new_Jinkela_wire_8347;
    wire new_Jinkela_wire_473;
    wire n_1350_;
    wire new_Jinkela_wire_288;
    wire new_Jinkela_wire_2722;
    wire new_Jinkela_wire_8911;
    wire new_Jinkela_wire_5005;
    wire new_Jinkela_wire_6;
    wire new_Jinkela_wire_2297;
    wire new_Jinkela_wire_8159;
    wire new_Jinkela_wire_6049;
    wire n_0856_;
    wire new_Jinkela_wire_9707;
    wire new_Jinkela_wire_10281;
    wire new_Jinkela_wire_9267;
    wire n_0443_;
    wire new_Jinkela_wire_5554;
    wire new_Jinkela_wire_7744;
    wire new_Jinkela_wire_8183;
    wire new_Jinkela_wire_7442;
    wire new_Jinkela_wire_9525;
    wire new_Jinkela_wire_2127;
    wire new_Jinkela_wire_7084;
    wire new_Jinkela_wire_10126;
    wire new_Jinkela_wire_831;
    wire new_Jinkela_wire_4251;
    wire new_Jinkela_wire_1370;
    wire new_Jinkela_wire_9637;
    wire new_Jinkela_wire_2437;
    wire new_Jinkela_wire_2321;
    wire n_1142_;
    wire new_Jinkela_wire_2737;
    wire new_Jinkela_wire_4826;
    wire new_Jinkela_wire_1095;
    wire new_Jinkela_wire_5809;
    wire new_Jinkela_wire_5970;
    wire new_Jinkela_wire_5175;
    wire new_Jinkela_wire_5899;
    wire new_Jinkela_wire_3266;
    wire new_Jinkela_wire_6738;
    wire new_Jinkela_wire_83;
    wire new_Jinkela_wire_5960;
    wire new_Jinkela_wire_5709;
    wire new_Jinkela_wire_9071;
    wire new_Jinkela_wire_9280;
    wire new_Jinkela_wire_9697;
    wire new_Jinkela_wire_7218;
    wire new_Jinkela_wire_7255;
    wire new_Jinkela_wire_375;
    wire n_0670_;
    wire new_Jinkela_wire_8714;
    wire new_Jinkela_wire_2754;
    wire new_Jinkela_wire_1093;
    wire new_Jinkela_wire_6434;
    wire new_Jinkela_wire_2959;
    wire new_Jinkela_wire_4958;
    wire new_Jinkela_wire_3323;
    wire new_Jinkela_wire_2589;
    wire new_Jinkela_wire_1164;
    wire new_Jinkela_wire_1698;
    wire new_Jinkela_wire_8454;
    wire new_Jinkela_wire_2009;
    wire new_Jinkela_wire_6351;
    wire new_Jinkela_wire_2996;
    wire new_Jinkela_wire_8008;
    wire new_Jinkela_wire_7972;
    wire new_Jinkela_wire_5998;
    wire new_Jinkela_wire_1365;
    wire new_Jinkela_wire_9768;
    wire new_Jinkela_wire_1593;
    wire new_Jinkela_wire_9460;
    wire new_Jinkela_wire_7541;
    wire new_Jinkela_wire_499;
    wire new_Jinkela_wire_1642;
    wire new_Jinkela_wire_1536;
    wire new_Jinkela_wire_3579;
    wire n_0648_;
    wire new_Jinkela_wire_4805;
    wire new_Jinkela_wire_6300;
    wire new_Jinkela_wire_4919;
    wire new_Jinkela_wire_5379;
    wire new_Jinkela_wire_4464;
    wire new_Jinkela_wire_8652;
    wire new_Jinkela_wire_2764;
    wire new_Jinkela_wire_6788;
    wire new_Jinkela_wire_5746;
    wire new_Jinkela_wire_8811;
    wire n_0921_;
    wire new_Jinkela_wire_6843;
    wire new_Jinkela_wire_10084;
    wire new_Jinkela_wire_9933;
    wire new_Jinkela_wire_6997;
    wire new_Jinkela_wire_2130;
    wire new_Jinkela_wire_3457;
    wire new_Jinkela_wire_3203;
    wire new_Jinkela_wire_1827;
    wire new_Jinkela_wire_5069;
    wire new_Jinkela_wire_9546;
    wire new_Jinkela_wire_2899;
    wire new_Jinkela_wire_4225;
    wire new_Jinkela_wire_2209;
    wire new_Jinkela_wire_9216;
    wire new_Jinkela_wire_5169;
    wire n_0510_;
    wire new_Jinkela_wire_7012;
    wire new_net_2529;
    wire new_Jinkela_wire_3854;
    wire new_Jinkela_wire_9201;
    wire new_Jinkela_wire_1332;
    wire new_Jinkela_wire_3207;
    wire new_Jinkela_wire_7159;
    wire new_Jinkela_wire_4486;
    wire new_Jinkela_wire_6904;
    wire new_Jinkela_wire_8368;
    wire new_Jinkela_wire_9009;
    wire new_Jinkela_wire_2674;
    wire new_Jinkela_wire_4977;
    wire new_Jinkela_wire_3530;
    wire new_Jinkela_wire_9865;
    wire new_Jinkela_wire_8374;
    wire new_Jinkela_wire_8133;
    wire new_Jinkela_wire_4274;
    wire new_Jinkela_wire_7731;
    wire new_Jinkela_wire_8259;
    wire n_0365_;
    wire new_Jinkela_wire_6414;
    wire new_Jinkela_wire_5882;
    wire new_Jinkela_wire_2605;
    wire new_Jinkela_wire_2688;
    wire new_Jinkela_wire_2915;
    wire new_Jinkela_wire_2866;
    wire new_Jinkela_wire_7740;
    wire n_1024_;
    wire new_Jinkela_wire_120;
    wire n_0551_;
    wire new_Jinkela_wire_3024;
    wire new_Jinkela_wire_7129;
    wire new_Jinkela_wire_487;
    wire new_Jinkela_wire_2159;
    wire new_Jinkela_wire_7068;
    wire n_1067_;
    wire new_Jinkela_wire_7761;
    wire new_Jinkela_wire_8847;
    wire new_Jinkela_wire_6206;
    wire new_Jinkela_wire_8431;
    wire new_Jinkela_wire_4442;
    wire new_Jinkela_wire_651;
    wire new_Jinkela_wire_3590;
    wire new_Jinkela_wire_180;
    wire new_Jinkela_wire_3931;
    wire new_Jinkela_wire_9361;
    wire new_Jinkela_wire_2268;
    wire new_Jinkela_wire_10120;
    wire n_0237_;
    wire new_Jinkela_wire_10325;
    wire new_Jinkela_wire_5557;
    wire new_Jinkela_wire_2973;
    wire new_Jinkela_wire_423;
    wire new_Jinkela_wire_10516;
    wire new_Jinkela_wire_3925;
    wire new_Jinkela_wire_2490;
    wire new_Jinkela_wire_2284;
    wire new_Jinkela_wire_5207;
    wire new_Jinkela_wire_6681;
    wire n_0996_;
    wire new_Jinkela_wire_1673;
    wire new_Jinkela_wire_2568;
    wire new_Jinkela_wire_869;
    wire new_Jinkela_wire_6710;
    wire new_Jinkela_wire_4384;
    wire new_Jinkela_wire_3474;
    wire new_Jinkela_wire_8575;
    wire new_Jinkela_wire_4743;
    wire new_Jinkela_wire_7377;
    wire new_Jinkela_wire_7508;
    wire new_Jinkela_wire_7853;
    wire new_Jinkela_wire_8382;
    wire new_Jinkela_wire_10113;
    wire n_0218_;
    wire n_0426_;
    wire new_Jinkela_wire_4571;
    wire new_Jinkela_wire_2173;
    wire new_Jinkela_wire_1594;
    wire new_Jinkela_wire_4912;
    wire new_Jinkela_wire_7236;
    wire new_Jinkela_wire_7260;
    wire new_Jinkela_wire_5346;
    wire new_Jinkela_wire_5349;
    wire new_Jinkela_wire_1747;
    wire new_Jinkela_wire_209;
    wire new_Jinkela_wire_7401;
    wire n_0965_;
    wire new_Jinkela_wire_6747;
    wire new_Jinkela_wire_4960;
    wire new_Jinkela_wire_848;
    wire new_Jinkela_wire_6079;
    wire new_Jinkela_wire_8859;
    wire new_Jinkela_wire_3815;
    wire new_Jinkela_wire_2255;
    wire new_Jinkela_wire_8854;
    wire new_Jinkela_wire_10537;
    wire new_Jinkela_wire_5820;
    wire new_Jinkela_wire_2518;
    wire new_Jinkela_wire_9247;
    wire new_Jinkela_wire_6485;
    wire new_Jinkela_wire_10544;
    wire new_Jinkela_wire_5761;
    wire new_Jinkela_wire_9169;
    wire new_Jinkela_wire_238;
    wire new_Jinkela_wire_1888;
    wire new_Jinkela_wire_4907;
    wire new_Jinkela_wire_7410;
    wire new_Jinkela_wire_2982;
    wire n_0356_;
    wire new_Jinkela_wire_2527;
    wire new_Jinkela_wire_7119;
    wire new_Jinkela_wire_10067;
    wire new_Jinkela_wire_8918;
    wire new_Jinkela_wire_1609;
    wire new_Jinkela_wire_5411;
    wire n_0032_;
    wire new_Jinkela_wire_9086;
    wire new_Jinkela_wire_7284;
    wire new_Jinkela_wire_2677;
    wire new_Jinkela_wire_4120;
    wire new_Jinkela_wire_6452;
    wire new_Jinkela_wire_2767;
    wire new_Jinkela_wire_554;
    wire new_Jinkela_wire_2950;
    wire new_Jinkela_wire_10158;
    wire new_Jinkela_wire_1000;
    wire new_Jinkela_wire_6549;
    wire new_Jinkela_wire_8132;
    wire new_Jinkela_wire_3125;
    wire new_Jinkela_wire_10236;
    wire new_Jinkela_wire_7651;
    wire n_1274_;
    wire new_Jinkela_wire_506;
    wire new_Jinkela_wire_7896;
    wire new_Jinkela_wire_1366;
    wire new_Jinkela_wire_1718;
    wire new_Jinkela_wire_7200;
    wire new_Jinkela_wire_7259;
    wire new_Jinkela_wire_7998;
    wire new_Jinkela_wire_4636;
    wire new_Jinkela_wire_4607;
    wire new_Jinkela_wire_1919;
    wire new_Jinkela_wire_10327;
    wire new_Jinkela_wire_6975;
    wire n_0738_;
    wire new_Jinkela_wire_1085;
    wire n_0094_;
    wire new_Jinkela_wire_4835;
    wire new_Jinkela_wire_317;
    wire new_Jinkela_wire_9778;
    wire new_Jinkela_wire_1414;
    wire new_Jinkela_wire_2088;
    wire new_Jinkela_wire_9930;
    wire new_Jinkela_wire_4501;
    wire new_Jinkela_wire_261;
    wire n_0391_;
    wire new_Jinkela_wire_2141;
    wire new_Jinkela_wire_7760;
    wire new_Jinkela_wire_1244;
    wire new_Jinkela_wire_5782;
    wire new_Jinkela_wire_8486;
    wire new_Jinkela_wire_2222;
    wire new_Jinkela_wire_1017;
    wire new_Jinkela_wire_4610;
    wire new_Jinkela_wire_5327;
    wire new_Jinkela_wire_4169;
    wire new_Jinkela_wire_5916;
    wire new_Jinkela_wire_2444;
    wire new_Jinkela_wire_9760;
    wire new_Jinkela_wire_9365;
    wire new_Jinkela_wire_2259;
    wire new_Jinkela_wire_8256;
    wire new_Jinkela_wire_968;
    wire n_1019_;
    wire new_Jinkela_wire_4100;
    wire new_Jinkela_wire_4310;
    wire new_Jinkela_wire_5643;
    wire new_Jinkela_wire_5347;
    wire new_Jinkela_wire_5250;
    wire new_Jinkela_wire_5874;
    wire new_Jinkela_wire_8788;
    wire new_Jinkela_wire_1425;
    wire new_Jinkela_wire_3807;
    wire new_Jinkela_wire_3249;
    wire n_1135_;
    wire new_Jinkela_wire_7145;
    wire new_Jinkela_wire_5676;
    wire new_Jinkela_wire_6731;
    wire new_Jinkela_wire_6869;
    wire new_Jinkela_wire_3654;
    wire new_Jinkela_wire_3735;
    wire new_Jinkela_wire_7424;
    wire new_Jinkela_wire_8277;
    wire new_Jinkela_wire_4507;
    wire new_Jinkela_wire_10254;
    wire n_0361_;
    wire new_Jinkela_wire_9224;
    wire new_Jinkela_wire_7980;
    wire new_Jinkela_wire_7478;
    wire new_Jinkela_wire_8420;
    wire new_Jinkela_wire_320;
    wire new_Jinkela_wire_9393;
    wire new_Jinkela_wire_747;
    wire new_Jinkela_wire_2445;
    wire new_Jinkela_wire_6185;
    wire new_Jinkela_wire_6649;
    wire new_Jinkela_wire_5906;
    wire new_Jinkela_wire_931;
    wire new_Jinkela_wire_3549;
    wire new_Jinkela_wire_3845;
    wire new_Jinkela_wire_1513;
    wire new_Jinkela_wire_5442;
    wire new_Jinkela_wire_909;
    wire new_Jinkela_wire_7411;
    wire new_Jinkela_wire_10240;
    wire new_Jinkela_wire_8915;
    wire new_Jinkela_wire_1819;
    wire n_0326_;
    wire new_Jinkela_wire_1807;
    wire new_Jinkela_wire_10458;
    wire new_Jinkela_wire_1899;
    wire new_Jinkela_wire_1252;
    wire new_Jinkela_wire_5564;
    wire new_Jinkela_wire_10262;
    wire new_Jinkela_wire_3982;
    wire new_Jinkela_wire_2064;
    wire n_0291_;
    wire new_Jinkela_wire_8292;
    wire new_Jinkela_wire_9880;
    wire new_Jinkela_wire_7573;
    wire new_Jinkela_wire_3671;
    wire new_Jinkela_wire_8267;
    wire new_Jinkela_wire_1957;
    wire new_Jinkela_wire_4672;
    wire n_0832_;
    wire new_Jinkela_wire_1837;
    wire new_Jinkela_wire_502;
    wire new_Jinkela_wire_1884;
    wire new_Jinkela_wire_7186;
    wire new_Jinkela_wire_1947;
    wire new_Jinkela_wire_276;
    wire new_Jinkela_wire_5402;
    wire new_Jinkela_wire_4931;
    wire new_Jinkela_wire_9671;
    wire new_Jinkela_wire_10159;
    wire new_Jinkela_wire_1659;
    wire new_Jinkela_wire_1310;
    wire new_Jinkela_wire_1933;
    wire new_Jinkela_wire_7487;
    wire new_Jinkela_wire_6164;
    wire new_Jinkela_wire_2505;
    wire new_Jinkela_wire_820;
    wire n_1023_;
    wire new_Jinkela_wire_2353;
    wire new_Jinkela_wire_3670;
    wire new_Jinkela_wire_1790;
    wire new_Jinkela_wire_3447;
    wire new_Jinkela_wire_2552;
    wire new_Jinkela_wire_530;
    wire new_Jinkela_wire_1412;
    wire new_Jinkela_wire_339;
    wire new_Jinkela_wire_2975;
    wire new_Jinkela_wire_2013;
    wire new_Jinkela_wire_4083;
    wire new_Jinkela_wire_7348;
    wire new_Jinkela_wire_1189;
    wire new_Jinkela_wire_923;
    wire new_Jinkela_wire_7834;
    wire new_Jinkela_wire_6554;
    wire new_Jinkela_wire_7539;
    wire new_Jinkela_wire_4832;
    wire new_Jinkela_wire_5477;
    wire n_1361_;
    wire n_1145_;
    wire new_Jinkela_wire_3103;
    wire new_Jinkela_wire_7872;
    wire new_Jinkela_wire_9420;
    wire new_Jinkela_wire_197;
    wire n_0933_;
    wire new_Jinkela_wire_4311;
    wire new_Jinkela_wire_2;
    wire new_Jinkela_wire_5529;
    wire new_Jinkela_wire_1736;
    wire new_Jinkela_wire_8635;
    wire new_Jinkela_wire_5910;
    wire new_Jinkela_wire_9501;
    wire new_Jinkela_wire_3057;
    wire new_Jinkela_wire_92;
    wire new_Jinkela_wire_1079;
    wire new_Jinkela_wire_5969;
    wire new_Jinkela_wire_6838;
    wire n_1155_;
    wire new_Jinkela_wire_9569;
    wire new_Jinkela_wire_3784;
    wire new_Jinkela_wire_5993;
    wire new_Jinkela_wire_4903;
    wire new_Jinkela_wire_3292;
    wire new_Jinkela_wire_9207;
    wire n_1004_;
    wire new_Jinkela_wire_6989;
    wire new_Jinkela_wire_7887;
    wire new_Jinkela_wire_10540;
    wire new_Jinkela_wire_8179;
    wire new_Jinkela_wire_8197;
    wire new_Jinkela_wire_1335;
    wire new_Jinkela_wire_10315;
    wire new_Jinkela_wire_2970;
    wire new_Jinkela_wire_3370;
    wire new_Jinkela_wire_8856;
    wire new_Jinkela_wire_8738;
    wire new_Jinkela_wire_1726;
    wire new_Jinkela_wire_5644;
    wire new_Jinkela_wire_7528;
    wire new_Jinkela_wire_6256;
    wire new_Jinkela_wire_5386;
    wire new_Jinkela_wire_3674;
    wire new_Jinkela_wire_7889;
    wire new_Jinkela_wire_2797;
    wire new_Jinkela_wire_2745;
    wire new_Jinkela_wire_5375;
    wire new_Jinkela_wire_8602;
    wire new_Jinkela_wire_7337;
    wire new_Jinkela_wire_1667;
    wire new_Jinkela_wire_5190;
    wire new_Jinkela_wire_941;
    wire new_Jinkela_wire_1903;
    wire new_Jinkela_wire_3778;
    wire new_Jinkela_wire_6633;
    wire new_Jinkela_wire_8113;
    wire new_Jinkela_wire_1616;
    wire new_Jinkela_wire_3302;
    wire new_Jinkela_wire_5119;
    wire new_Jinkela_wire_10081;
    wire new_net_2527;
    wire new_Jinkela_wire_3467;
    wire n_1348_;
    wire new_Jinkela_wire_5131;
    wire n_0519_;
    wire n_0462_;
    wire n_1261_;
    wire new_Jinkela_wire_5735;
    wire new_Jinkela_wire_1586;
    wire new_Jinkela_wire_7287;
    wire new_Jinkela_wire_9817;
    wire n_1132_;
    wire new_Jinkela_wire_4989;
    wire new_Jinkela_wire_1376;
    wire new_Jinkela_wire_10383;
    wire new_Jinkela_wire_3212;
    wire new_Jinkela_wire_6480;
    wire new_Jinkela_wire_8895;
    wire n_0752_;
    wire new_Jinkela_wire_9399;
    wire new_Jinkela_wire_9046;
    wire new_Jinkela_wire_4117;
    wire new_Jinkela_wire_9484;
    wire new_Jinkela_wire_10178;
    wire new_Jinkela_wire_2695;
    wire new_Jinkela_wire_5057;
    wire n_0591_;
    wire new_Jinkela_wire_5027;
    wire new_Jinkela_wire_10272;
    wire new_Jinkela_wire_9136;
    wire new_Jinkela_wire_287;
    wire new_Jinkela_wire_300;
    wire new_Jinkela_wire_10422;
    wire n_1214_;
    wire new_Jinkela_wire_5600;
    wire new_Jinkela_wire_8657;
    wire new_Jinkela_wire_7154;
    wire new_Jinkela_wire_5114;
    wire new_Jinkela_wire_4099;
    wire n_0513_;
    wire new_Jinkela_wire_2457;
    wire new_Jinkela_wire_6878;
    wire new_Jinkela_wire_2121;
    wire new_Jinkela_wire_664;
    wire n_1181_;
    wire new_Jinkela_wire_4971;
    wire new_Jinkela_wire_6606;
    wire new_Jinkela_wire_5605;
    wire n_1223_;
    wire new_Jinkela_wire_10260;
    wire new_Jinkela_wire_7115;
    wire n_0034_;
    wire new_Jinkela_wire_4721;
    wire new_Jinkela_wire_10056;
    wire new_Jinkela_wire_4008;
    wire new_Jinkela_wire_10072;
    wire new_Jinkela_wire_10014;
    wire new_Jinkela_wire_8234;
    wire new_Jinkela_wire_8298;
    wire new_Jinkela_wire_6413;
    wire n_0076_;
    wire new_Jinkela_wire_6353;
    wire n_0726_;
    wire new_Jinkela_wire_1186;
    wire new_Jinkela_wire_5025;
    wire new_Jinkela_wire_3440;
    wire new_Jinkela_wire_9369;
    wire n_0938_;
    wire new_Jinkela_wire_2547;
    wire n_0117_;
    wire new_Jinkela_wire_3030;
    wire new_Jinkela_wire_1183;
    wire new_Jinkela_wire_4041;
    wire new_Jinkela_wire_8775;
    wire new_Jinkela_wire_9206;
    wire new_Jinkela_wire_8111;
    wire n_0976_;
    wire new_Jinkela_wire_3646;
    wire new_Jinkela_wire_4286;
    wire new_Jinkela_wire_1910;
    wire new_Jinkela_wire_8219;
    wire new_Jinkela_wire_2503;
    wire new_Jinkela_wire_1701;
    wire new_Jinkela_wire_2062;
    wire new_Jinkela_wire_7181;
    wire n_1157_;
    wire new_Jinkela_wire_7770;
    wire new_Jinkela_wire_9379;
    wire n_0758_;
    wire new_Jinkela_wire_3917;
    wire new_Jinkela_wire_10097;
    wire new_Jinkela_wire_2262;
    wire n_0408_;
    wire new_Jinkela_wire_5297;
    wire n_1088_;
    wire new_Jinkela_wire_5341;
    wire new_Jinkela_wire_6562;
    wire new_Jinkela_wire_5793;
    wire new_Jinkela_wire_9320;
    wire new_Jinkela_wire_7815;
    wire new_Jinkela_wire_4738;
    wire new_Jinkela_wire_2856;
    wire new_Jinkela_wire_9801;
    wire new_Jinkela_wire_7488;
    wire new_Jinkela_wire_1923;
    wire new_Jinkela_wire_8323;
    wire new_Jinkela_wire_10074;
    wire new_Jinkela_wire_9423;
    wire new_Jinkela_wire_9424;
    wire new_Jinkela_wire_215;
    wire new_Jinkela_wire_4635;
    wire new_Jinkela_wire_3000;
    wire n_0753_;
    wire new_Jinkela_wire_303;
    wire new_Jinkela_wire_289;
    wire new_Jinkela_wire_9605;
    wire new_Jinkela_wire_6042;
    wire n_0012_;
    wire n_0932_;
    wire new_Jinkela_wire_4282;
    wire new_Jinkela_wire_10208;
    wire new_Jinkela_wire_9722;
    wire new_Jinkela_wire_3004;
    wire new_Jinkela_wire_374;
    wire new_Jinkela_wire_10013;
    wire new_Jinkela_wire_4420;
    wire new_Jinkela_wire_1377;
    wire new_Jinkela_wire_133;
    wire new_Jinkela_wire_9631;
    wire new_Jinkela_wire_2077;
    wire new_Jinkela_wire_10286;
    wire new_Jinkela_wire_1639;
    wire n_0262_;
    wire new_Jinkela_wire_5660;
    wire new_Jinkela_wire_6333;
    wire new_Jinkela_wire_5145;
    wire new_Jinkela_wire_2022;
    wire new_Jinkela_wire_4189;
    wire new_Jinkela_wire_3396;
    wire new_Jinkela_wire_7292;
    wire new_Jinkela_wire_2908;
    wire new_Jinkela_wire_6835;
    wire n_0385_;
    wire n_0668_;
    wire new_Jinkela_wire_5351;
    wire new_Jinkela_wire_7639;
    wire new_Jinkela_wire_7080;
    wire new_Jinkela_wire_8751;
    wire new_Jinkela_wire_9607;
    wire new_Jinkela_wire_1898;
    wire new_Jinkela_wire_1999;
    wire new_Jinkela_wire_7375;
    wire new_Jinkela_wire_8631;
    wire new_Jinkela_wire_10049;
    wire new_Jinkela_wire_4431;
    wire new_Jinkela_wire_5521;
    wire new_Jinkela_wire_8802;
    wire new_Jinkela_wire_4887;
    wire new_Jinkela_wire_727;
    wire new_Jinkela_wire_2100;
    wire new_Jinkela_wire_7721;
    wire new_Jinkela_wire_855;
    wire new_Jinkela_wire_4;
    wire new_Jinkela_wire_6356;
    wire n_0276_;
    wire new_Jinkela_wire_10623;
    wire new_Jinkela_wire_4076;
    wire n_0364_;
    wire new_Jinkela_wire_5513;
    wire new_Jinkela_wire_7203;
    wire n_0878_;
    wire new_Jinkela_wire_1611;
    wire new_Jinkela_wire_4595;
    wire new_Jinkela_wire_6254;
    wire new_Jinkela_wire_3617;
    wire new_Jinkela_wire_1514;
    wire n_0524_;
    wire new_Jinkela_wire_1958;
    wire new_Jinkela_wire_9465;
    wire new_Jinkela_wire_1173;
    wire new_Jinkela_wire_7128;
    wire new_Jinkela_wire_3659;
    wire new_Jinkela_wire_7357;
    wire new_Jinkela_wire_6966;
    wire new_Jinkela_wire_1267;
    wire new_Jinkela_wire_3133;
    wire new_Jinkela_wire_1391;
    wire new_Jinkela_wire_7627;
    wire n_0285_;
    wire new_Jinkela_wire_8246;
    wire new_Jinkela_wire_5831;
    wire new_Jinkela_wire_2249;
    wire new_Jinkela_wire_6388;
    wire new_Jinkela_wire_9652;
    wire new_Jinkela_wire_4717;
    wire new_Jinkela_wire_4722;
    wire new_Jinkela_wire_5176;
    wire new_Jinkela_wire_2063;
    wire new_Jinkela_wire_5657;
    wire new_Jinkela_wire_813;
    wire new_Jinkela_wire_7900;
    wire new_Jinkela_wire_8358;
    wire new_Jinkela_wire_4375;
    wire new_Jinkela_wire_2476;
    wire n_0275_;
    wire new_Jinkela_wire_8350;
    wire new_Jinkela_wire_10135;
    wire n_1093_;
    wire new_Jinkela_wire_5627;
    wire new_Jinkela_wire_23;
    wire new_Jinkela_wire_9162;
    wire new_Jinkela_wire_8659;
    wire new_Jinkela_wire_7509;
    wire new_Jinkela_wire_2708;
    wire new_Jinkela_wire_3772;
    wire n_0341_;
    wire new_Jinkela_wire_4667;
    wire new_Jinkela_wire_7013;
    wire new_Jinkela_wire_2317;
    wire n_0198_;
    wire new_Jinkela_wire_1260;
    wire new_Jinkela_wire_1689;
    wire new_Jinkela_wire_2512;
    wire new_Jinkela_wire_9396;
    wire new_Jinkela_wire_9227;
    wire new_Jinkela_wire_9070;
    wire new_Jinkela_wire_6809;
    wire new_Jinkela_wire_6347;
    wire new_Jinkela_wire_643;
    wire new_Jinkela_wire_10407;
    wire new_Jinkela_wire_5285;
    wire new_Jinkela_wire_6435;
    wire new_Jinkela_wire_3015;
    wire new_Jinkela_wire_1179;
    wire new_Jinkela_wire_5302;
    wire new_Jinkela_wire_1061;
    wire new_Jinkela_wire_9906;
    wire new_Jinkela_wire_2749;
    wire new_Jinkela_wire_8683;
    wire new_Jinkela_wire_5673;
    wire new_Jinkela_wire_2156;
    wire new_Jinkela_wire_5888;
    wire new_Jinkela_wire_1240;
    wire new_Jinkela_wire_1596;
    wire new_Jinkela_wire_3993;
    wire new_Jinkela_wire_44;
    wire new_Jinkela_wire_543;
    wire new_Jinkela_wire_10124;
    wire new_Jinkela_wire_4527;
    wire new_Jinkela_wire_1913;
    wire new_Jinkela_wire_6216;
    wire new_Jinkela_wire_9405;
    wire n_0458_;
    wire new_Jinkela_wire_4293;
    wire new_Jinkela_wire_9634;
    wire new_Jinkela_wire_2432;
    wire new_Jinkela_wire_1259;
    wire new_Jinkela_wire_1934;
    wire new_Jinkela_wire_4028;
    wire n_0142_;
    wire new_Jinkela_wire_3886;
    wire new_Jinkela_wire_623;
    wire n_0335_;
    wire new_Jinkela_wire_1012;
    wire new_Jinkela_wire_3347;
    wire new_Jinkela_wire_2661;
    wire new_Jinkela_wire_59;
    wire new_Jinkela_wire_9571;
    wire new_Jinkela_wire_3995;
    wire new_Jinkela_wire_7183;
    wire new_Jinkela_wire_993;
    wire new_Jinkela_wire_3025;
    wire new_Jinkela_wire_2684;
    wire new_Jinkela_wire_9294;
    wire new_Jinkela_wire_1123;
    wire new_Jinkela_wire_4766;
    wire new_Jinkela_wire_8782;
    wire new_Jinkela_wire_9000;
    wire new_Jinkela_wire_6172;
    wire new_Jinkela_wire_8459;
    wire new_Jinkela_wire_4290;
    wire n_0822_;
    wire n_0953_;
    wire new_Jinkela_wire_3524;
    wire new_Jinkela_wire_10297;
    wire new_Jinkela_wire_9443;
    wire new_Jinkela_wire_3773;
    wire new_Jinkela_wire_3639;
    wire new_Jinkela_wire_10538;
    wire new_Jinkela_wire_8992;
    wire new_Jinkela_wire_10207;
    wire new_Jinkela_wire_7524;
    wire new_Jinkela_wire_10276;
    wire new_Jinkela_wire_7054;
    wire new_Jinkela_wire_686;
    wire new_Jinkela_wire_5171;
    wire new_Jinkela_wire_9735;
    wire new_Jinkela_wire_8763;
    wire new_Jinkela_wire_3279;
    wire new_Jinkela_wire_1833;
    wire new_Jinkela_wire_8127;
    wire new_Jinkela_wire_281;
    wire new_Jinkela_wire_8803;
    wire new_Jinkela_wire_4862;
    wire new_Jinkela_wire_7583;
    wire new_Jinkela_wire_4629;
    wire new_Jinkela_wire_2347;
    wire new_Jinkela_wire_3724;
    wire new_Jinkela_wire_4834;
    wire new_Jinkela_wire_1499;
    wire new_Jinkela_wire_177;
    wire new_Jinkela_wire_5317;
    wire new_Jinkela_wire_3461;
    wire new_Jinkela_wire_2955;
    wire new_Jinkela_wire_6350;
    wire new_Jinkela_wire_7249;
    wire new_Jinkela_wire_8029;
    wire new_Jinkela_wire_1127;
    wire new_Jinkela_wire_4261;
    wire new_Jinkela_wire_2898;
    wire new_Jinkela_wire_5844;
    wire n_0161_;
    wire new_Jinkela_wire_1745;
    wire new_Jinkela_wire_6283;
    wire new_Jinkela_wire_321;
    wire new_Jinkela_wire_4487;
    wire new_Jinkela_wire_3252;
    wire new_Jinkela_wire_3860;
    wire new_net_2503;
    wire new_Jinkela_wire_2501;
    wire new_Jinkela_wire_7347;
    wire n_0128_;
    wire new_Jinkela_wire_1818;
    wire new_Jinkela_wire_7611;
    wire new_Jinkela_wire_6081;
    wire new_Jinkela_wire_9999;
    wire new_Jinkela_wire_7626;
    wire new_Jinkela_wire_4433;
    wire new_Jinkela_wire_9966;
    wire new_Jinkela_wire_9781;
    wire new_Jinkela_wire_2112;
    wire new_Jinkela_wire_2160;
    wire new_Jinkela_wire_3762;
    wire new_Jinkela_wire_9627;
    wire new_Jinkela_wire_9187;
    wire new_Jinkela_wire_4474;
    wire new_Jinkela_wire_7641;
    wire n_0617_;
    wire n_0308_;
    wire new_Jinkela_wire_4191;
    wire new_Jinkela_wire_9771;
    wire n_0464_;
    wire new_Jinkela_wire_10359;
    wire n_0983_;
    wire new_Jinkela_wire_10188;
    wire new_Jinkela_wire_1830;
    wire new_Jinkela_wire_2479;
    wire new_Jinkela_wire_5006;
    wire new_Jinkela_wire_3436;
    wire new_Jinkela_wire_9064;
    wire new_Jinkela_wire_5021;
    wire n_0620_;
    wire new_Jinkela_wire_1680;
    wire new_Jinkela_wire_3909;
    wire n_1021_;
    wire new_Jinkela_wire_9316;
    wire n_1177_;
    wire new_Jinkela_wire_7824;
    wire new_Jinkela_wire_3454;
    wire new_Jinkela_wire_8302;
    wire new_Jinkela_wire_9248;
    wire new_Jinkela_wire_3426;
    wire new_Jinkela_wire_1859;
    wire new_Jinkela_wire_4814;
    wire new_Jinkela_wire_10256;
    wire new_Jinkela_wire_3708;
    wire new_Jinkela_wire_7981;
    wire new_Jinkela_wire_6971;
    wire new_Jinkela_wire_6016;
    wire new_Jinkela_wire_3318;
    wire new_Jinkela_wire_6504;
    wire new_Jinkela_wire_5493;
    wire new_Jinkela_wire_6866;
    wire new_Jinkela_wire_4489;
    wire new_Jinkela_wire_10411;
    wire new_Jinkela_wire_4057;
    wire new_Jinkela_wire_9737;
    wire new_Jinkela_wire_5764;
    wire new_Jinkela_wire_7874;
    wire new_Jinkela_wire_6366;
    wire new_Jinkela_wire_7914;
    wire new_Jinkela_wire_350;
    wire new_Jinkela_wire_263;
    wire new_Jinkela_wire_8908;
    wire new_Jinkela_wire_3959;
    wire n_0781_;
    wire new_Jinkela_wire_9618;
    wire new_Jinkela_wire_415;
    wire new_Jinkela_wire_4256;
    wire new_Jinkela_wire_2430;
    wire new_Jinkela_wire_5032;
    wire new_Jinkela_wire_4590;
    wire n_0881_;
    wire new_Jinkela_wire_9255;
    wire new_Jinkela_wire_7506;
    wire new_Jinkela_wire_10273;
    wire new_Jinkela_wire_3322;
    wire new_Jinkela_wire_2981;
    wire new_Jinkela_wire_3295;
    wire new_Jinkela_wire_3381;
    wire new_Jinkela_wire_3696;
    wire n_0703_;
    wire new_Jinkela_wire_10080;
    wire new_Jinkela_wire_2023;
    wire new_Jinkela_wire_279;
    wire n_1281_;
    wire new_Jinkela_wire_9495;
    wire new_Jinkela_wire_6640;
    wire new_Jinkela_wire_421;
    wire n_0740_;
    wire new_Jinkela_wire_7383;
    wire new_Jinkela_wire_881;
    wire new_Jinkela_wire_6083;
    wire new_Jinkela_wire_7213;
    wire new_Jinkela_wire_6893;
    wire new_Jinkela_wire_8681;
    wire new_Jinkela_wire_8377;
    wire new_Jinkela_wire_4976;
    wire n_0154_;
    wire new_Jinkela_wire_9272;
    wire new_Jinkela_wire_2798;
    wire new_Jinkela_wire_1121;
    wire new_Jinkela_wire_5273;
    wire new_Jinkela_wire_7620;
    wire new_Jinkela_wire_7156;
    wire new_Jinkela_wire_6652;
    wire new_Jinkela_wire_9145;
    wire new_Jinkela_wire_8819;
    wire new_Jinkela_wire_8872;
    wire new_net_2513;
    wire new_Jinkela_wire_7243;
    wire new_Jinkela_wire_4035;
    wire new_Jinkela_wire_7599;
    wire new_Jinkela_wire_13;
    wire new_Jinkela_wire_2382;
    wire new_Jinkela_wire_4245;
    wire new_Jinkela_wire_5370;
    wire new_Jinkela_wire_2655;
    wire new_Jinkela_wire_2958;
    wire new_Jinkela_wire_9066;
    wire new_Jinkela_wire_3072;
    wire new_Jinkela_wire_4402;
    wire new_Jinkela_wire_3139;
    wire new_Jinkela_wire_4644;
    wire new_Jinkela_wire_7247;
    wire new_Jinkela_wire_7416;
    wire new_Jinkela_wire_3044;
    wire n_1312_;
    wire new_Jinkela_wire_4600;
    wire new_Jinkela_wire_2224;
    wire new_Jinkela_wire_5781;
    wire new_Jinkela_wire_9503;
    wire new_Jinkela_wire_1808;
    wire new_Jinkela_wire_9654;
    wire new_Jinkela_wire_7006;
    wire new_Jinkela_wire_2387;
    wire new_Jinkela_wire_4588;
    wire new_Jinkela_wire_8262;
    wire new_Jinkela_wire_8306;
    wire new_Jinkela_wire_4147;
    wire n_0476_;
    wire new_Jinkela_wire_4390;
    wire n_0543_;
    wire new_Jinkela_wire_3277;
    wire new_Jinkela_wire_6996;
    wire new_Jinkela_wire_1507;
    wire new_Jinkela_wire_7795;
    wire new_Jinkela_wire_4363;
    wire new_Jinkela_wire_9717;
    wire new_Jinkela_wire_7251;
    wire new_Jinkela_wire_1396;
    wire new_Jinkela_wire_3766;
    wire new_Jinkela_wire_3944;
    wire new_Jinkela_wire_1483;
    wire new_Jinkela_wire_5084;
    wire new_Jinkela_wire_8680;
    wire new_Jinkela_wire_6465;
    wire n_1167_;
    wire new_Jinkela_wire_10307;
    wire new_Jinkela_wire_8175;
    wire new_Jinkela_wire_7189;
    wire new_Jinkela_wire_5825;
    wire new_Jinkela_wire_841;
    wire new_Jinkela_wire_2433;
    wire new_Jinkela_wire_8320;
    wire new_Jinkela_wire_7113;
    wire new_Jinkela_wire_521;
    wire n_0901_;
    wire new_Jinkela_wire_8318;
    wire new_Jinkela_wire_4867;
    wire new_Jinkela_wire_8471;
    wire new_Jinkela_wire_1426;
    wire new_Jinkela_wire_5247;
    wire new_Jinkela_wire_6919;
    wire new_Jinkela_wire_7548;
    wire new_Jinkela_wire_8253;
    wire new_Jinkela_wire_4675;
    wire new_Jinkela_wire_2978;
    wire new_Jinkela_wire_1774;
    wire n_0825_;
    wire new_Jinkela_wire_8913;
    wire n_1277_;
    wire new_Jinkela_wire_9762;
    wire n_1010_;
    wire new_Jinkela_wire_1381;
    wire new_Jinkela_wire_10417;
    wire new_Jinkela_wire_8619;
    wire new_Jinkela_wire_1815;
    wire new_Jinkela_wire_5788;
    wire new_Jinkela_wire_712;
    wire new_Jinkela_wire_4429;
    wire n_0789_;
    wire new_Jinkela_wire_6798;
    wire new_Jinkela_wire_2635;
    wire new_Jinkela_wire_9237;
    wire new_Jinkela_wire_6526;
    wire new_Jinkela_wire_8989;
    wire new_Jinkela_wire_6712;
    wire new_Jinkela_wire_3582;
    wire new_Jinkela_wire_5162;
    wire new_Jinkela_wire_3930;
    wire new_Jinkela_wire_3153;
    wire new_Jinkela_wire_1678;
    wire new_Jinkela_wire_3865;
    wire new_Jinkela_wire_8421;
    wire new_Jinkela_wire_8467;
    wire n_0008_;
    wire new_Jinkela_wire_1226;
    wire new_Jinkela_wire_6870;
    wire new_Jinkela_wire_9731;
    wire new_Jinkela_wire_9558;
    wire n_0452_;
    wire new_Jinkela_wire_7051;
    wire new_Jinkela_wire_600;
    wire new_Jinkela_wire_8171;
    wire new_Jinkela_wire_9324;
    wire new_Jinkela_wire_6579;
    wire new_Jinkela_wire_2741;
    wire new_Jinkela_wire_314;
    wire new_Jinkela_wire_10280;
    wire new_Jinkela_wire_3777;
    wire new_Jinkela_wire_181;
    wire new_Jinkela_wire_3026;
    wire new_Jinkela_wire_10020;
    wire n_0501_;
    wire new_Jinkela_wire_5249;
    wire new_Jinkela_wire_2215;
    wire new_Jinkela_wire_6469;
    wire new_Jinkela_wire_2718;
    wire new_Jinkela_wire_6910;
    wire new_Jinkela_wire_4797;
    wire new_Jinkela_wire_8107;
    wire new_Jinkela_wire_4564;
    wire new_Jinkela_wire_10142;
    wire n_1036_;
    wire new_Jinkela_wire_5827;
    wire new_Jinkela_wire_3033;
    wire new_Jinkela_wire_9039;
    wire new_Jinkela_wire_8119;
    wire new_Jinkela_wire_9716;
    wire new_Jinkela_wire_6946;
    wire new_Jinkela_wire_3733;
    wire n_1128_;
    wire new_Jinkela_wire_10563;
    wire n_1125_;
    wire new_Jinkela_wire_9062;
    wire new_Jinkela_wire_6677;
    wire new_Jinkela_wire_10376;
    wire new_Jinkela_wire_4677;
    wire new_Jinkela_wire_9193;
    wire new_Jinkela_wire_2469;
    wire new_Jinkela_wire_1952;
    wire new_Jinkela_wire_7036;
    wire new_Jinkela_wire_6722;
    wire new_Jinkela_wire_1636;
    wire new_Jinkela_wire_6766;
    wire new_Jinkela_wire_6459;
    wire new_Jinkela_wire_5368;
    wire new_Jinkela_wire_3351;
    wire new_Jinkela_wire_6200;
    wire new_Jinkela_wire_1469;
    wire new_Jinkela_wire_9319;
    wire new_Jinkela_wire_4855;
    wire new_Jinkela_wire_5092;
    wire n_0306_;
    wire new_Jinkela_wire_6189;
    wire new_Jinkela_wire_8783;
    wire new_Jinkela_wire_7621;
    wire new_Jinkela_wire_5034;
    wire new_Jinkela_wire_4016;
    wire new_Jinkela_wire_8378;
    wire new_Jinkela_wire_1280;
    wire new_Jinkela_wire_2598;
    wire new_Jinkela_wire_5854;
    wire n_0393_;
    wire new_Jinkela_wire_6994;
    wire n_0320_;
    wire new_Jinkela_wire_3746;
    wire new_Jinkela_wire_4969;
    wire new_Jinkela_wire_1768;
    wire new_Jinkela_wire_10600;
    wire new_Jinkela_wire_8417;
    wire n_0494_;
    wire new_Jinkela_wire_1046;
    wire new_Jinkela_wire_2341;
    wire new_Jinkela_wire_4504;
    wire new_Jinkela_wire_2296;
    wire new_Jinkela_wire_2613;
    wire new_Jinkela_wire_8387;
    wire new_Jinkela_wire_7501;
    wire new_Jinkela_wire_2454;
    wire new_Jinkela_wire_3626;
    wire new_Jinkela_wire_5414;
    wire new_Jinkela_wire_6426;
    wire new_Jinkela_wire_1006;
    wire new_Jinkela_wire_4250;
    wire new_Jinkela_wire_810;
    wire new_Jinkela_wire_8556;
    wire new_Jinkela_wire_2587;
    wire new_Jinkela_wire_4150;
    wire new_Jinkela_wire_3145;
    wire n_0687_;
    wire n_0084_;
    wire new_Jinkela_wire_5049;
    wire new_Jinkela_wire_9015;
    wire new_Jinkela_wire_2199;
    wire new_Jinkela_wire_5174;
    wire new_Jinkela_wire_1730;
    wire new_Jinkela_wire_10571;
    wire new_Jinkela_wire_8054;
    wire new_Jinkela_wire_580;
    wire new_Jinkela_wire_3701;
    wire new_Jinkela_wire_2287;
    wire new_Jinkela_wire_8835;
    wire new_Jinkela_wire_844;
    wire new_Jinkela_wire_2323;
    wire new_Jinkela_wire_3750;
    wire new_Jinkela_wire_10514;
    wire new_Jinkela_wire_1606;
    wire new_Jinkela_wire_9485;
    wire new_Jinkela_wire_9354;
    wire new_Jinkela_wire_6023;
    wire n_0043_;
    wire new_Jinkela_wire_7346;
    wire new_Jinkela_wire_9796;
    wire new_Jinkela_wire_7850;
    wire new_Jinkela_wire_9991;
    wire n_0665_;
    wire new_Jinkela_wire_9303;
    wire new_Jinkela_wire_5769;
    wire new_Jinkela_wire_10501;
    wire new_Jinkela_wire_6982;
    wire new_Jinkela_wire_10497;
    wire new_Jinkela_wire_6262;
    wire new_Jinkela_wire_4043;
    wire new_Jinkela_wire_647;
    wire new_Jinkela_wire_1044;
    wire new_Jinkela_wire_8479;
    wire new_Jinkela_wire_6656;
    wire new_Jinkela_wire_2953;
    wire new_Jinkela_wire_3656;
    wire new_Jinkela_wire_606;
    wire new_Jinkela_wire_7464;
    wire new_Jinkela_wire_9980;
    wire new_Jinkela_wire_3492;
    wire new_Jinkela_wire_6764;
    wire new_Jinkela_wire_1865;
    wire new_Jinkela_wire_4040;
    wire new_Jinkela_wire_7564;
    wire new_Jinkela_wire_9597;
    wire n_0027_;
    wire n_0310_;
    wire new_Jinkela_wire_2841;
    wire new_Jinkela_wire_3663;
    wire new_Jinkela_wire_1027;
    wire new_Jinkela_wire_1089;
    wire new_Jinkela_wire_2858;
    wire new_Jinkela_wire_5857;
    wire n_0867_;
    wire new_Jinkela_wire_4828;
    wire new_Jinkela_wire_4913;
    wire new_Jinkela_wire_2994;
    wire new_Jinkela_wire_10548;
    wire new_Jinkela_wire_7996;
    wire new_Jinkela_wire_8039;
    wire new_Jinkela_wire_3489;
    wire new_Jinkela_wire_2954;
    wire new_Jinkela_wire_7253;
    wire new_Jinkela_wire_442;
    wire new_Jinkela_wire_1937;
    wire new_Jinkela_wire_6038;
    wire new_net_8;
    wire new_Jinkela_wire_10238;
    wire new_Jinkela_wire_5543;
    wire new_Jinkela_wire_1692;
    wire new_Jinkela_wire_7206;
    wire new_Jinkela_wire_10266;
    wire new_Jinkela_wire_8369;
    wire new_Jinkela_wire_7139;
    wire new_Jinkela_wire_1669;
    wire new_Jinkela_wire_10421;
    wire new_Jinkela_wire_1022;
    wire new_Jinkela_wire_9055;
    wire new_Jinkela_wire_429;
    wire new_Jinkela_wire_2863;
    wire new_Jinkela_wire_4961;
    wire new_Jinkela_wire_8785;
    wire new_Jinkela_wire_1219;
    wire new_Jinkela_wire_9538;
    wire new_Jinkela_wire_9921;
    wire new_Jinkela_wire_6392;
    wire new_Jinkela_wire_3175;
    wire new_Jinkela_wire_8886;
    wire new_Jinkela_wire_4015;
    wire new_Jinkela_wire_657;
    wire new_Jinkela_wire_7852;
    wire new_Jinkela_wire_6727;
    wire new_Jinkela_wire_6134;
    wire new_Jinkela_wire_10583;
    wire new_Jinkela_wire_5929;
    wire new_Jinkela_wire_1389;
    wire new_Jinkela_wire_3014;
    wire new_Jinkela_wire_560;
    wire new_Jinkela_wire_3201;
    wire new_Jinkela_wire_9275;
    wire new_Jinkela_wire_4413;
    wire new_Jinkela_wire_76;
    wire new_Jinkela_wire_10324;
    wire new_Jinkela_wire_6319;
    wire new_Jinkela_wire_4372;
    wire new_Jinkela_wire_1349;
    wire new_Jinkela_wire_5683;
    wire n_0058_;
    wire new_Jinkela_wire_3420;
    wire new_Jinkela_wire_9057;
    wire new_Jinkela_wire_10275;
    wire new_Jinkela_wire_5441;
    wire new_Jinkela_wire_9391;
    wire new_Jinkela_wire_8498;
    wire new_Jinkela_wire_9257;
    wire new_Jinkela_wire_2868;
    wire new_Jinkela_wire_8875;
    wire new_Jinkela_wire_3797;
    wire new_Jinkela_wire_1713;
    wire new_Jinkela_wire_1045;
    wire new_Jinkela_wire_9407;
    wire new_Jinkela_wire_4258;
    wire new_Jinkela_wire_2517;
    wire new_Jinkela_wire_9969;
    wire new_Jinkela_wire_9101;
    wire new_Jinkela_wire_8476;
    wire new_Jinkela_wire_6789;
    wire new_Jinkela_wire_8359;
    wire new_Jinkela_wire_27;
    wire new_Jinkela_wire_9011;
    wire new_Jinkela_wire_10227;
    wire new_Jinkela_wire_765;
    wire new_Jinkela_wire_10331;
    wire new_Jinkela_wire_2851;
    wire new_Jinkela_wire_8904;
    wire new_Jinkela_wire_4818;
    wire new_Jinkela_wire_9342;
    wire n_0656_;
    wire new_Jinkela_wire_8041;
    wire new_Jinkela_wire_3045;
    wire new_Jinkela_wire_2554;
    wire new_Jinkela_wire_6728;
    wire new_Jinkela_wire_5802;
    wire n_0861_;
    wire new_Jinkela_wire_1221;
    wire new_Jinkela_wire_7617;
    wire new_Jinkela_wire_6906;
    wire new_Jinkela_wire_66;
    wire new_Jinkela_wire_8121;
    wire new_Jinkela_wire_7836;
    wire new_Jinkela_wire_526;
    wire new_Jinkela_wire_4360;
    wire n_0642_;
    wire new_Jinkela_wire_7316;
    wire new_Jinkela_wire_3150;
    wire new_Jinkela_wire_3607;
    wire new_Jinkela_wire_7153;
    wire new_Jinkela_wire_439;
    wire new_Jinkela_wire_8887;
    wire new_Jinkela_wire_4909;
    wire new_Jinkela_wire_997;
    wire new_Jinkela_wire_8897;
    wire new_Jinkela_wire_4901;
    wire new_net_2558;
    wire new_Jinkela_wire_3592;
    wire new_Jinkela_wire_7444;
    wire new_Jinkela_wire_6191;
    wire new_Jinkela_wire_3937;
    wire n_1269_;
    wire new_Jinkela_wire_4141;
    wire new_Jinkela_wire_9684;
    wire new_Jinkela_wire_8301;
    wire new_Jinkela_wire_2873;
    wire new_Jinkela_wire_10029;
    wire new_Jinkela_wire_872;
    wire new_Jinkela_wire_3435;
    wire new_Jinkela_wire_10232;
    wire new_Jinkela_wire_7202;
    wire new_Jinkela_wire_2799;
    wire new_Jinkela_wire_5920;
    wire new_Jinkela_wire_2016;
    wire new_Jinkela_wire_8495;
    wire n_0362_;
    wire new_Jinkela_wire_4227;
    wire n_1198_;
    wire new_Jinkela_wire_2405;
    wire new_Jinkela_wire_6698;
    wire new_Jinkela_wire_4148;
    wire new_Jinkela_wire_7669;
    wire n_0855_;
    wire new_Jinkela_wire_10290;
    wire new_Jinkela_wire_3268;
    wire n_1055_;
    wire new_Jinkela_wire_4868;
    wire new_Jinkela_wire_5212;
    wire new_Jinkela_wire_10493;
    wire new_Jinkela_wire_4090;
    wire new_Jinkela_wire_2526;
    wire new_Jinkela_wire_1617;
    wire new_Jinkela_wire_917;
    wire new_Jinkela_wire_9886;
    wire new_Jinkela_wire_9155;
    wire new_Jinkela_wire_4840;
    wire new_Jinkela_wire_5473;
    wire new_Jinkela_wire_10562;
    wire new_Jinkela_wire_5044;
    wire new_Jinkela_wire_3174;
    wire new_Jinkela_wire_8760;
    wire new_Jinkela_wire_5281;
    wire n_1032_;
    wire new_Jinkela_wire_2413;
    wire new_Jinkela_wire_4156;
    wire new_Jinkela_wire_10009;
    wire n_1100_;
    wire new_Jinkela_wire_5893;
    wire n_0966_;
    wire new_Jinkela_wire_5195;
    wire new_Jinkela_wire_7716;
    wire new_Jinkela_wire_7417;
    wire new_Jinkela_wire_8532;
    wire new_Jinkela_wire_8185;
    wire new_Jinkela_wire_729;
    wire new_Jinkela_wire_9765;
    wire n_0517_;
    wire new_Jinkela_wire_9352;
    wire new_Jinkela_wire_7462;
    wire n_1194_;
    wire new_Jinkela_wire_10099;
    wire new_Jinkela_wire_7995;
    wire new_Jinkela_wire_9988;
    wire new_Jinkela_wire_9059;
    wire new_Jinkela_wire_6309;
    wire new_Jinkela_wire_8433;
    wire new_Jinkela_wire_5108;
    wire n_0357_;
    wire new_Jinkela_wire_211;
    wire n_0700_;
    wire new_Jinkela_wire_1357;
    wire new_Jinkela_wire_9785;
    wire new_Jinkela_wire_8601;
    wire n_0549_;
    wire new_Jinkela_wire_497;
    wire new_Jinkela_wire_9277;
    wire new_Jinkela_wire_1118;
    wire new_Jinkela_wire_6045;
    wire new_Jinkela_wire_8776;
    wire n_0149_;
    wire new_Jinkela_wire_8283;
    wire new_Jinkela_wire_1465;
    wire new_Jinkela_wire_3493;
    wire new_Jinkela_wire_2852;
    wire new_Jinkela_wire_4247;
    wire n_0202_;
    wire new_Jinkela_wire_10508;
    wire new_Jinkela_wire_5934;
    wire new_Jinkela_wire_274;
    wire new_Jinkela_wire_7630;
    wire n_0654_;
    wire new_Jinkela_wire_6827;
    wire new_Jinkela_wire_304;
    wire n_0104_;
    wire new_Jinkela_wire_10569;
    wire new_Jinkela_wire_10311;
    wire new_Jinkela_wire_8850;
    wire new_Jinkela_wire_1169;
    wire new_Jinkela_wire_4703;
    wire n_0995_;
    wire new_Jinkela_wire_6826;
    wire new_Jinkela_wire_3998;
    wire new_Jinkela_wire_5445;
    wire new_Jinkela_wire_10330;
    wire new_Jinkela_wire_3477;
    wire new_Jinkela_wire_7345;
    wire n_0609_;
    wire n_0869_;
    wire new_Jinkela_wire_4955;
    wire new_Jinkela_wire_7885;
    wire new_Jinkela_wire_10341;
    wire new_Jinkela_wire_7575;
    wire new_Jinkela_wire_9992;
    wire new_Jinkela_wire_5211;
    wire new_Jinkela_wire_3789;
    wire new_Jinkela_wire_8709;
    wire new_Jinkela_wire_4582;
    wire new_Jinkela_wire_919;
    wire new_Jinkela_wire_10464;
    wire new_Jinkela_wire_5633;
    wire new_Jinkela_wire_2411;
    wire new_Jinkela_wire_9807;
    wire new_Jinkela_wire_2869;
    wire new_Jinkela_wire_2435;
    wire new_Jinkela_wire_2370;
    wire new_Jinkela_wire_6854;
    wire new_Jinkela_wire_9564;
    wire n_0400_;
    wire new_Jinkela_wire_2352;
    wire new_Jinkela_wire_5421;
    wire new_Jinkela_wire_7520;
    wire new_Jinkela_wire_7654;
    wire new_Jinkela_wire_10109;
    wire new_Jinkela_wire_4981;
    wire n_0906_;
    wire new_Jinkela_wire_7011;
    wire new_Jinkela_wire_9822;
    wire new_Jinkela_wire_5748;
    wire new_Jinkela_wire_8799;
    wire new_Jinkela_wire_1094;
    wire new_Jinkela_wire_8214;
    wire new_Jinkela_wire_6118;
    wire new_Jinkela_wire_7144;
    wire new_Jinkela_wire_4389;
    wire new_Jinkela_wire_7455;
    wire new_Jinkela_wire_4356;
    wire new_Jinkela_wire_5479;
    wire new_Jinkela_wire_6258;
    wire new_Jinkela_wire_8174;
    wire n_0795_;
    wire n_1329_;
    wire new_Jinkela_wire_10582;
    wire new_Jinkela_wire_6131;
    wire new_Jinkela_wire_6391;
    wire new_Jinkela_wire_5740;
    wire new_Jinkela_wire_7434;
    wire new_Jinkela_wire_8411;
    wire new_Jinkela_wire_7120;
    wire new_net_2554;
    wire new_Jinkela_wire_6880;
    wire new_Jinkela_wire_2417;
    wire new_Jinkela_wire_5772;
    wire n_0913_;
    wire new_Jinkela_wire_4396;
    wire new_Jinkela_wire_7735;
    wire new_Jinkela_wire_7675;
    wire new_Jinkela_wire_2577;
    wire new_Jinkela_wire_6657;
    wire new_Jinkela_wire_6800;
    wire new_Jinkela_wire_4233;
    wire new_Jinkela_wire_5776;
    wire new_Jinkela_wire_1798;
    wire new_Jinkela_wire_4648;
    wire new_Jinkela_wire_3505;
    wire new_Jinkela_wire_5095;
    wire new_Jinkela_wire_2030;
    wire new_Jinkela_wire_201;
    wire new_Jinkela_wire_8163;
    wire new_Jinkela_wire_4110;
    wire new_Jinkela_wire_735;
    wire new_Jinkela_wire_8313;
    wire new_Jinkela_wire_8941;
    wire n_0131_;
    wire new_Jinkela_wire_7312;
    wire new_Jinkela_wire_8146;
    wire new_Jinkela_wire_9549;
    wire new_Jinkela_wire_8422;
    wire new_Jinkela_wire_2068;
    wire new_Jinkela_wire_10334;
    wire new_Jinkela_wire_5541;
    wire new_Jinkela_wire_3387;
    wire new_Jinkela_wire_4619;
    wire new_Jinkela_wire_5385;
    wire new_Jinkela_wire_10149;
    wire new_Jinkela_wire_4920;
    wire new_Jinkela_wire_1190;
    wire new_Jinkela_wire_4202;
    wire n_0250_;
    wire new_Jinkela_wire_6105;
    wire new_Jinkela_wire_9533;
    wire new_Jinkela_wire_4260;
    wire new_Jinkela_wire_9875;
    wire new_Jinkela_wire_545;
    wire new_Jinkela_wire_3158;
    wire new_Jinkela_wire_4950;
    wire new_Jinkela_wire_5298;
    wire new_Jinkela_wire_3776;
    wire n_0367_;
    wire new_Jinkela_wire_9209;
    wire new_Jinkela_wire_5200;
    wire new_Jinkela_wire_7707;
    wire new_Jinkela_wire_2450;
    wire new_Jinkela_wire_8932;
    wire new_Jinkela_wire_8451;
    wire new_Jinkela_wire_5528;
    wire new_Jinkela_wire_1540;
    wire new_Jinkela_wire_5109;
    wire n_0277_;
    wire new_Jinkela_wire_1360;
    wire new_Jinkela_wire_8275;
    wire new_Jinkela_wire_9803;
    wire new_Jinkela_wire_8724;
    wire new_Jinkela_wire_6294;
    wire new_Jinkela_wire_7065;
    wire new_Jinkela_wire_7538;
    wire new_Jinkela_wire_5444;
    wire new_Jinkela_wire_9073;
    wire new_Jinkela_wire_5775;
    wire new_Jinkela_wire_3731;
    wire new_Jinkela_wire_8062;
    wire new_Jinkela_wire_6519;
    wire new_Jinkela_wire_10495;
    wire new_Jinkela_wire_4463;
    wire new_Jinkela_wire_4536;
    wire new_Jinkela_wire_4806;
    wire new_Jinkela_wire_5124;
    wire n_0073_;
    wire new_Jinkela_wire_10507;
    wire new_Jinkela_wire_5367;
    wire new_Jinkela_wire_8645;
    wire new_Jinkela_wire_494;
    wire new_Jinkela_wire_832;
    wire new_Jinkela_wire_3534;
    wire new_Jinkela_wire_2059;
    wire n_0643_;
    wire new_Jinkela_wire_3754;
    wire new_Jinkela_wire_4638;
    wire new_Jinkela_wire_9914;
    wire new_Jinkela_wire_10131;
    wire new_Jinkela_wire_8543;
    wire new_Jinkela_wire_1737;
    wire n_0425_;
    wire new_Jinkela_wire_4932;
    wire new_Jinkela_wire_6004;
    wire new_Jinkela_wire_7004;
    wire n_0489_;
    wire n_0274_;
    wire new_Jinkela_wire_5571;
    wire new_Jinkela_wire_4775;
    wire new_Jinkela_wire_9385;
    wire new_Jinkela_wire_8808;
    wire new_Jinkela_wire_7655;
    wire new_Jinkela_wire_995;
    wire new_Jinkela_wire_9435;
    wire new_Jinkela_wire_1620;
    wire new_Jinkela_wire_8231;
    wire new_Jinkela_wire_1497;
    wire new_Jinkela_wire_4483;
    wire new_Jinkela_wire_9053;
    wire new_Jinkela_wire_7463;
    wire new_Jinkela_wire_9751;
    wire new_Jinkela_wire_9467;
    wire new_Jinkela_wire_3105;
    wire new_Jinkela_wire_5029;
    wire new_Jinkela_wire_10063;
    wire n_0962_;
    wire new_Jinkela_wire_2178;
    wire new_Jinkela_wire_45;
    wire n_1253_;
    wire n_0049_;
    wire new_Jinkela_wire_3037;
    wire new_Jinkela_wire_9953;
    wire new_Jinkela_wire_9740;
    wire new_Jinkela_wire_7680;
    wire new_Jinkela_wire_9995;
    wire new_Jinkela_wire_3427;
    wire new_Jinkela_wire_1227;
    wire new_Jinkela_wire_3642;
    wire n_1079_;
    wire new_Jinkela_wire_406;
    wire n_0009_;
    wire new_Jinkela_wire_758;
    wire new_Jinkela_wire_9302;
    wire new_Jinkela_wire_6692;
    wire new_Jinkela_wire_9378;
    wire new_Jinkela_wire_10500;
    wire n_0820_;
    wire new_Jinkela_wire_4967;
    wire new_Jinkela_wire_5214;
    wire new_Jinkela_wire_1430;
    wire new_net_2547;
    wire new_Jinkela_wire_4292;
    wire new_Jinkela_wire_1831;
    wire new_Jinkela_wire_9186;
    wire new_Jinkela_wire_9314;
    wire new_Jinkela_wire_4962;
    wire new_Jinkela_wire_7282;
    wire new_Jinkela_wire_7551;
    wire new_Jinkela_wire_7911;
    wire new_Jinkela_wire_6103;
    wire n_0089_;
    wire new_Jinkela_wire_10462;
    wire new_Jinkela_wire_767;
    wire new_Jinkela_wire_10034;
    wire new_Jinkela_wire_7052;
    wire new_Jinkela_wire_8793;
    wire new_Jinkela_wire_7846;
    wire new_Jinkela_wire_10058;
    wire new_Jinkela_wire_9641;
    wire new_Jinkela_wire_8679;
    wire new_Jinkela_wire_1887;
    wire new_Jinkela_wire_2892;
    wire new_Jinkela_wire_5023;
    wire new_Jinkela_wire_6926;
    wire new_Jinkela_wire_1728;
    wire new_Jinkela_wire_2671;
    wire new_Jinkela_wire_2622;
    wire new_Jinkela_wire_1257;
    wire new_Jinkela_wire_5921;
    wire n_0622_;
    wire new_Jinkela_wire_1784;
    wire new_Jinkela_wire_4742;
    wire new_Jinkela_wire_4218;
    wire new_Jinkela_wire_6371;
    wire new_Jinkela_wire_6777;
    wire new_Jinkela_wire_3775;
    wire new_Jinkela_wire_6548;
    wire new_Jinkela_wire_8995;
    wire new_Jinkela_wire_7229;
    wire new_Jinkela_wire_9163;
    wire new_Jinkela_wire_1520;
    wire new_Jinkela_wire_1170;
    wire new_Jinkela_wire_6292;
    wire new_Jinkela_wire_8356;
    wire new_Jinkela_wire_6441;
    wire new_Jinkela_wire_4441;
    wire new_Jinkela_wire_7415;
    wire new_Jinkela_wire_10558;
    wire new_Jinkela_wire_7171;
    wire n_0121_;
    wire new_Jinkela_wire_8630;
    wire new_Jinkela_wire_10300;
    wire new_Jinkela_wire_7578;
    wire new_Jinkela_wire_8167;
    wire new_Jinkela_wire_10329;
    wire new_Jinkela_wire_8965;
    wire new_Jinkela_wire_1311;
    wire new_Jinkela_wire_1314;
    wire new_Jinkela_wire_8295;
    wire new_Jinkela_wire_3485;
    wire new_Jinkela_wire_1206;
    wire new_Jinkela_wire_4621;
    wire new_Jinkela_wire_9321;
    wire n_0318_;
    wire new_Jinkela_wire_8721;
    wire new_Jinkela_wire_3231;
    wire new_Jinkela_wire_3180;
    wire new_Jinkela_wire_5104;
    wire new_Jinkela_wire_2146;
    wire new_Jinkela_wire_9103;
    wire new_Jinkela_wire_408;
    wire new_Jinkela_wire_2006;
    wire new_Jinkela_wire_8829;
    wire new_Jinkela_wire_3628;
    wire new_Jinkela_wire_7050;
    wire new_Jinkela_wire_10101;
    wire new_Jinkela_wire_230;
    wire new_Jinkela_wire_2992;
    wire new_Jinkela_wire_10136;
    wire n_0934_;
    wire new_Jinkela_wire_1398;
    wire n_0814_;
    wire new_Jinkela_wire_5264;
    wire new_Jinkela_wire_741;
    wire new_Jinkela_wire_10130;
    wire new_Jinkela_wire_7340;
    wire new_Jinkela_wire_6043;
    wire new_Jinkela_wire_2453;
    wire new_Jinkela_wire_10343;
    wire new_Jinkela_wire_6876;
    wire new_Jinkela_wire_450;
    wire new_Jinkela_wire_2085;
    wire new_Jinkela_wire_9343;
    wire new_Jinkela_wire_1941;
    wire new_Jinkela_wire_836;
    wire new_Jinkela_wire_10104;
    wire new_Jinkela_wire_8774;
    wire n_1317_;
    wire new_Jinkela_wire_9944;
    wire n_0112_;
    wire new_Jinkela_wire_7604;
    wire new_Jinkela_wire_7044;
    wire new_Jinkela_wire_9171;
    wire new_Jinkela_wire_6221;
    wire new_Jinkela_wire_6065;
    wire new_Jinkela_wire_3565;
    wire new_Jinkela_wire_9244;
    wire new_Jinkela_wire_1556;
    wire new_Jinkela_wire_2149;
    wire new_Jinkela_wire_7963;
    wire new_Jinkela_wire_2987;
    wire new_Jinkela_wire_1874;
    wire new_Jinkela_wire_7039;
    wire new_Jinkela_wire_3368;
    wire new_Jinkela_wire_6173;
    wire new_Jinkela_wire_2585;
    wire new_Jinkela_wire_6980;
    wire new_Jinkela_wire_793;
    wire new_Jinkela_wire_9262;
    wire new_Jinkela_wire_7055;
    wire new_Jinkela_wire_6639;
    wire n_0203_;
    wire new_Jinkela_wire_1547;
    wire new_Jinkela_wire_7954;
    wire new_Jinkela_wire_2769;
    wire new_Jinkela_wire_4299;
    wire new_Jinkela_wire_4628;
    wire new_Jinkela_wire_1388;
    wire new_Jinkela_wire_3885;
    wire new_Jinkela_wire_3720;
    wire new_Jinkela_wire_9021;
    wire n_0583_;
    wire new_Jinkela_wire_10156;
    wire new_Jinkela_wire_6274;
    wire new_net_11;
    wire new_Jinkela_wire_1591;
    wire n_0383_;
    wire n_0610_;
    wire new_Jinkela_wire_399;
    wire new_Jinkela_wire_4854;
    wire new_Jinkela_wire_6743;
    wire new_Jinkela_wire_7275;
    wire new_Jinkela_wire_8003;
    wire new_Jinkela_wire_5755;
    wire new_Jinkela_wire_7137;
    wire new_Jinkela_wire_5407;
    wire new_Jinkela_wire_5384;
    wire new_Jinkela_wire_6625;
    wire n_0833_;
    wire new_Jinkela_wire_7134;
    wire new_Jinkela_wire_4674;
    wire new_Jinkela_wire_5343;
    wire new_Jinkela_wire_10075;
    wire new_Jinkela_wire_10002;
    wire new_Jinkela_wire_2302;
    wire new_Jinkela_wire_7787;
    wire new_Jinkela_wire_6923;
    wire new_Jinkela_wire_1869;
    wire n_0138_;
    wire new_Jinkela_wire_10449;
    wire new_Jinkela_wire_7503;
    wire new_Jinkela_wire_9565;
    wire new_Jinkela_wire_2529;
    wire n_1047_;
    wire new_Jinkela_wire_2425;
    wire new_Jinkela_wire_778;
    wire n_0115_;
    wire new_Jinkela_wire_1168;
    wire new_Jinkela_wire_6988;
    wire new_Jinkela_wire_2031;
    wire new_Jinkela_wire_2119;
    wire new_Jinkela_wire_10148;
    wire new_Jinkela_wire_3173;
    wire new_Jinkela_wire_9976;
    wire n_0580_;
    wire new_Jinkela_wire_6207;
    wire new_Jinkela_wire_4221;
    wire n_0000_;
    wire new_Jinkela_wire_6167;
    wire new_Jinkela_wire_6984;
    wire new_Jinkela_wire_3584;
    wire new_Jinkela_wire_3091;
    wire n_1234_;
    wire new_Jinkela_wire_9266;
    wire new_Jinkela_wire_2814;
    wire new_Jinkela_wire_5714;
    wire new_Jinkela_wire_3195;
    wire new_Jinkela_wire_5423;
    wire new_Jinkela_wire_4664;
    wire new_Jinkela_wire_2281;
    wire new_Jinkela_wire_7175;
    wire n_0099_;
    wire new_Jinkela_wire_459;
    wire new_Jinkela_wire_10616;
    wire new_Jinkela_wire_6423;
    wire new_Jinkela_wire_5845;
    wire new_Jinkela_wire_4831;
    wire new_Jinkela_wire_4581;
    wire new_Jinkela_wire_9029;
    wire new_Jinkela_wire_4212;
    wire new_Jinkela_wire_3556;
    wire new_Jinkela_wire_5710;
    wire new_net_2574;
    wire new_Jinkela_wire_3924;
    wire new_Jinkela_wire_4668;
    wire new_Jinkela_wire_8383;
    wire new_Jinkela_wire_4017;
    wire new_Jinkela_wire_10107;
    wire new_Jinkela_wire_649;
    wire n_1333_;
    wire new_Jinkela_wire_10328;
    wire n_0671_;
    wire new_Jinkela_wire_221;
    wire new_Jinkela_wire_5456;
    wire new_Jinkela_wire_2555;
    wire n_0205_;
    wire new_Jinkela_wire_1608;
    wire new_Jinkela_wire_9033;
    wire new_Jinkela_wire_4565;
    wire new_Jinkela_wire_9366;
    wire new_Jinkela_wire_4625;
    wire new_Jinkela_wire_2857;
    wire new_Jinkela_wire_7172;
    wire new_Jinkela_wire_3929;
    wire new_Jinkela_wire_333;
    wire n_0194_;
    wire new_Jinkela_wire_10420;
    wire new_Jinkela_wire_4991;
    wire new_Jinkela_wire_10174;
    wire new_Jinkela_wire_2250;
    wire new_Jinkela_wire_6691;
    wire new_Jinkela_wire_2438;
    wire new_Jinkela_wire_6762;
    wire new_Jinkela_wire_5397;
    wire new_Jinkela_wire_989;
    wire new_Jinkela_wire_218;
    wire n_1263_;
    wire new_Jinkela_wire_7468;
    wire new_Jinkela_wire_8072;
    wire new_Jinkela_wire_131;
    wire new_Jinkela_wire_2363;
    wire new_Jinkela_wire_260;
    wire new_Jinkela_wire_6184;
    wire new_Jinkela_wire_1900;
    wire new_Jinkela_wire_5305;
    wire new_Jinkela_wire_10314;
    wire new_Jinkela_wire_5648;
    wire new_Jinkela_wire_7664;
    wire new_Jinkela_wire_962;
    wire new_Jinkela_wire_7102;
    wire new_Jinkela_wire_8715;
    wire new_Jinkela_wire_5612;
    wire new_Jinkela_wire_9837;
    wire new_Jinkela_wire_7890;
    wire n_0471_;
    wire new_Jinkela_wire_3035;
    wire n_0081_;
    wire new_Jinkela_wire_6979;
    wire new_Jinkela_wire_8701;
    wire new_Jinkela_wire_8468;
    wire new_Jinkela_wire_8128;
    wire new_Jinkela_wire_9258;
    wire new_Jinkela_wire_6620;
    wire n_0834_;
    wire new_Jinkela_wire_6359;
    wire new_Jinkela_wire_8110;
    wire n_0171_;
    wire new_Jinkela_wire_6818;
    wire n_0566_;
    wire new_Jinkela_wire_461;
    wire n_0722_;
    wire new_Jinkela_wire_8653;
    wire new_Jinkela_wire_5420;
    wire new_Jinkela_wire_5707;
    wire new_Jinkela_wire_2545;
    wire new_Jinkela_wire_8425;
    wire new_Jinkela_wire_409;
    wire new_Jinkela_wire_10313;
    wire new_Jinkela_wire_7965;
    wire new_Jinkela_wire_4850;
    wire new_Jinkela_wire_6429;
    wire new_Jinkela_wire_8150;
    wire n_0547_;
    wire new_Jinkela_wire_4080;
    wire new_Jinkela_wire_3453;
    wire new_Jinkela_wire_9037;
    wire n_1062_;
    wire new_Jinkela_wire_4317;
    wire new_Jinkela_wire_8478;
    wire new_Jinkela_wire_5747;
    wire new_Jinkela_wire_8021;
    wire new_Jinkela_wire_10561;
    wire new_Jinkela_wire_10519;
    wire new_Jinkela_wire_3736;
    wire new_Jinkela_wire_9889;
    wire new_Jinkela_wire_5763;
    wire n_1164_;
    wire new_Jinkela_wire_10586;
    wire new_Jinkela_wire_9450;
    wire new_Jinkela_wire_6403;
    wire new_Jinkela_wire_3594;
    wire new_Jinkela_wire_2979;
    wire new_Jinkela_wire_6718;
    wire new_Jinkela_wire_6384;
    wire new_Jinkela_wire_8140;
    wire new_Jinkela_wire_8972;
    wire new_Jinkela_wire_3512;
    wire n_1286_;
    wire new_Jinkela_wire_6047;
    wire new_Jinkela_wire_8734;
    wire new_Jinkela_wire_6453;
    wire new_Jinkela_wire_10379;
    wire n_1003_;
    wire n_0186_;
    wire new_Jinkela_wire_4566;
    wire new_Jinkela_wire_7327;
    wire new_Jinkela_wire_7216;
    wire new_Jinkela_wire_1857;
    wire new_Jinkela_wire_4939;
    wire new_Jinkela_wire_10506;
    wire new_Jinkela_wire_2180;
    wire new_Jinkela_wire_9235;
    wire new_Jinkela_wire_4633;
    wire new_Jinkela_wire_1302;
    wire new_Jinkela_wire_4249;
    wire new_Jinkela_wire_10191;
    wire new_Jinkela_wire_9217;
    wire new_Jinkela_wire_5242;
    wire new_Jinkela_wire_878;
    wire new_Jinkela_wire_10038;
    wire new_Jinkela_wire_877;
    wire new_Jinkela_wire_3739;
    wire n_1334_;
    wire new_Jinkela_wire_1362;
    wire new_Jinkela_wire_8622;
    wire n_0959_;
    wire new_Jinkela_wire_5448;
    wire new_Jinkela_wire_8866;
    wire new_Jinkela_wire_1662;
    wire new_Jinkela_wire_2812;
    wire new_Jinkela_wire_5336;
    wire new_Jinkela_wire_8685;
    wire new_Jinkela_wire_589;
    wire new_Jinkela_wire_7304;
    wire new_Jinkela_wire_6170;
    wire new_Jinkela_wire_7262;
    wire new_Jinkela_wire_8813;
    wire new_Jinkela_wire_1067;
    wire new_Jinkela_wire_1217;
    wire new_Jinkela_wire_4368;
    wire new_Jinkela_wire_2073;
    wire new_Jinkela_wire_10414;
    wire new_Jinkela_wire_4520;
    wire new_Jinkela_wire_6828;
    wire new_Jinkela_wire_3090;
    wire new_Jinkela_wire_7367;
    wire new_Jinkela_wire_713;
    wire new_Jinkela_wire_1848;
    wire new_Jinkela_wire_6683;
    wire new_Jinkela_wire_6443;
    wire new_Jinkela_wire_1158;
    wire new_Jinkela_wire_3922;
    wire n_0975_;
    wire new_Jinkela_wire_9827;
    wire new_Jinkela_wire_5394;
    wire new_Jinkela_wire_3110;
    wire new_Jinkela_wire_4620;
    wire new_Jinkela_wire_2721;
    wire new_Jinkela_wire_1605;
    wire new_Jinkela_wire_8853;
    wire new_Jinkela_wire_5206;
    wire new_Jinkela_wire_5099;
    wire new_Jinkela_wire_8504;
    wire new_Jinkela_wire_10252;
    wire n_0296_;
    wire new_Jinkela_wire_1270;
    wire new_Jinkela_wire_7001;
    wire n_0558_;
    wire new_Jinkela_wire_596;
    wire n_0106_;
    wire new_Jinkela_wire_1776;
    wire new_Jinkela_wire_1823;
    wire n_0905_;
    wire new_Jinkela_wire_1119;
    wire new_Jinkela_wire_4005;
    wire new_Jinkela_wire_10441;
    wire new_Jinkela_wire_4986;
    wire new_Jinkela_wire_4567;
    wire n_0456_;
    wire new_Jinkela_wire_10090;
    wire new_Jinkela_wire_6990;
    wire new_Jinkela_wire_6144;
    wire new_Jinkela_wire_7748;
    wire new_Jinkela_wire_1759;
    wire n_0497_;
    wire new_Jinkela_wire_455;
    wire new_Jinkela_wire_9050;
    wire new_Jinkela_wire_7067;
    wire new_Jinkela_wire_7936;
    wire n_1328_;
    wire new_Jinkela_wire_822;
    wire new_Jinkela_wire_7877;
    wire new_Jinkela_wire_7763;
    wire new_Jinkela_wire_5434;
    wire new_Jinkela_wire_9329;
    wire new_Jinkela_wire_97;
    wire new_Jinkela_wire_5220;
    wire new_Jinkela_wire_125;
    wire n_0392_;
    wire new_Jinkela_wire_861;
    wire new_Jinkela_wire_7659;
    wire new_Jinkela_wire_7220;
    wire new_Jinkela_wire_549;
    wire new_Jinkela_wire_4037;
    wire new_Jinkela_wire_927;
    wire new_Jinkela_wire_8165;
    wire new_Jinkela_wire_6193;
    wire new_Jinkela_wire_6578;
    wire new_Jinkela_wire_3065;
    wire new_Jinkela_wire_10363;
    wire new_Jinkela_wire_7943;
    wire new_Jinkela_wire_149;
    wire new_Jinkela_wire_9973;
    wire n_0545_;
    wire new_Jinkela_wire_1677;
    wire new_Jinkela_wire_5724;
    wire new_Jinkela_wire_4782;
    wire new_Jinkela_wire_8825;
    wire new_Jinkela_wire_269;
    wire new_Jinkela_wire_2825;
    wire new_Jinkela_wire_283;
    wire new_Jinkela_wire_1436;
    wire new_Jinkela_wire_4062;
    wire new_Jinkela_wire_2849;
    wire new_Jinkela_wire_797;
    wire new_Jinkela_wire_7851;
    wire new_Jinkela_wire_8678;
    wire new_Jinkela_wire_7209;
    wire new_Jinkela_wire_4355;
    wire new_Jinkela_wire_3805;
    wire new_Jinkela_wire_690;
    wire new_Jinkela_wire_7718;
    wire new_Jinkela_wire_705;
    wire new_Jinkela_wire_7597;
    wire new_Jinkela_wire_6246;
    wire new_Jinkela_wire_363;
    wire new_Jinkela_wire_56;
    wire n_0666_;
    wire new_Jinkela_wire_10505;
    wire new_Jinkela_wire_5126;
    wire new_Jinkela_wire_8749;
    wire new_Jinkela_wire_3373;
    wire new_Jinkela_wire_380;
    wire new_Jinkela_wire_7435;
    wire new_Jinkela_wire_6364;
    wire new_Jinkela_wire_9412;
    wire new_Jinkela_wire_9516;
    wire new_Jinkela_wire_4934;
    wire new_Jinkela_wire_8116;
    wire new_Jinkela_wire_4999;
    wire n_1228_;
    wire new_Jinkela_wire_7598;
    wire new_Jinkela_wire_1564;
    wire n_0139_;
    wire new_Jinkela_wire_158;
    wire new_Jinkela_wire_2980;
    wire new_Jinkela_wire_7391;
    wire new_Jinkela_wire_6836;
    wire new_Jinkela_wire_7090;
    wire new_Jinkela_wire_8258;
    wire new_Jinkela_wire_515;
    wire new_Jinkela_wire_7801;
    wire new_Jinkela_wire_9357;
    wire new_Jinkela_wire_8472;
    wire new_Jinkela_wire_4578;
    wire n_0624_;
    wire n_0838_;
    wire new_Jinkela_wire_9704;
    wire new_Jinkela_wire_2590;
    wire new_Jinkela_wire_7693;
    wire new_Jinkela_wire_453;
    wire n_0260_;
    wire new_Jinkela_wire_3273;
    wire new_Jinkela_wire_812;
    wire n_0560_;
    wire n_0258_;
    wire new_Jinkela_wire_8603;
    wire new_Jinkela_wire_3200;
    wire new_Jinkela_wire_3828;
    wire new_Jinkela_wire_952;
    wire new_Jinkela_wire_7016;
    wire new_Jinkela_wire_4264;
    wire new_Jinkela_wire_6325;
    wire new_Jinkela_wire_9739;
    wire new_Jinkela_wire_6296;
    wire new_Jinkela_wire_8357;
    wire new_Jinkela_wire_1623;
    wire new_Jinkela_wire_8460;
    wire new_Jinkela_wire_9718;
    wire n_0096_;
    wire new_Jinkela_wire_5512;
    wire n_0329_;
    wire n_1355_;
    wire new_Jinkela_wire_9578;
    wire n_0571_;
    wire new_Jinkela_wire_2366;
    wire n_0374_;
    wire new_Jinkela_wire_8212;
    wire new_Jinkela_wire_10193;
    wire new_Jinkela_wire_7450;
    wire new_Jinkela_wire_7930;
    wire new_Jinkela_wire_7606;
    wire new_Jinkela_wire_8370;
    wire new_Jinkela_wire_1953;
    wire new_Jinkela_wire_10619;
    wire new_Jinkela_wire_9168;
    wire new_Jinkela_wire_5985;
    wire new_Jinkela_wire_293;
    wire new_Jinkela_wire_10592;
    wire new_Jinkela_wire_4516;
    wire n_1354_;
    wire new_Jinkela_wire_620;
    wire new_Jinkela_wire_627;
    wire new_Jinkela_wire_2096;
    wire new_Jinkela_wire_1585;
    wire new_Jinkela_wire_2372;
    wire new_Jinkela_wire_6867;
    wire new_Jinkela_wire_6314;
    wire new_Jinkela_wire_2536;
    wire new_Jinkela_wire_9336;
    wire new_Jinkela_wire_7211;
    wire new_Jinkela_wire_5974;
    wire new_Jinkela_wire_4614;
    wire new_Jinkela_wire_6594;
    wire new_Jinkela_wire_10459;
    wire new_Jinkela_wire_1216;
    wire new_Jinkela_wire_7166;
    wire new_Jinkela_wire_8117;
    wire new_Jinkela_wire_7955;
    wire new_Jinkela_wire_9402;
    wire new_Jinkela_wire_4755;
    wire new_Jinkela_wire_8329;
    wire new_Jinkela_wire_3863;
    wire new_Jinkela_wire_10;
    wire n_0678_;
    wire n_1338_;
    wire new_Jinkela_wire_322;
    wire new_Jinkela_wire_5185;
    wire new_net_2564;
    wire new_Jinkela_wire_4383;
    wire new_Jinkela_wire_4851;
    wire new_Jinkela_wire_5324;
    wire n_0325_;
    wire new_Jinkela_wire_8966;
    wire n_0815_;
    wire n_0924_;
    wire new_Jinkela_wire_7921;
    wire n_0813_;
    wire new_Jinkela_wire_10016;
    wire new_Jinkela_wire_498;
    wire new_Jinkela_wire_10609;
    wire new_Jinkela_wire_602;
    wire new_Jinkela_wire_6424;
    wire new_Jinkela_wire_1106;
    wire new_Jinkela_wire_5146;
    wire new_Jinkela_wire_4243;
    wire new_Jinkela_wire_1545;
    wire new_Jinkela_wire_4780;
    wire n_0108_;
    wire new_Jinkela_wire_6506;
    wire new_net_2537;
    wire new_Jinkela_wire_7909;
    wire new_Jinkela_wire_4295;
    wire new_Jinkela_wire_4316;
    wire new_Jinkela_wire_1167;
    wire new_Jinkela_wire_2792;
    wire new_Jinkela_wire_3369;
    wire new_Jinkela_wire_2486;
    wire new_Jinkela_wire_443;
    wire new_Jinkela_wire_6310;
    wire new_Jinkela_wire_785;
    wire new_Jinkela_wire_1050;
    wire new_Jinkela_wire_2239;
    wire new_Jinkela_wire_8798;
    wire new_Jinkela_wire_7300;
    wire new_Jinkela_wire_1915;
    wire new_Jinkela_wire_7857;
    wire new_Jinkela_wire_7542;
    wire new_Jinkela_wire_4597;
    wire new_Jinkela_wire_6013;
    wire new_Jinkela_wire_1407;
    wire new_Jinkela_wire_5510;
    wire new_Jinkela_wire_753;
    wire new_Jinkela_wire_5912;
    wire new_Jinkela_wire_3247;
    wire new_Jinkela_wire_311;
    wire new_Jinkela_wire_206;
    wire new_Jinkela_wire_9541;
    wire new_Jinkela_wire_4364;
    wire n_1048_;
    wire new_Jinkela_wire_4896;
    wire n_0303_;
    wire n_0340_;
    wire new_Jinkela_wire_5572;
    wire new_Jinkela_wire_2723;
    wire n_0750_;
    wire new_Jinkela_wire_8429;
    wire new_Jinkela_wire_3438;
    wire new_Jinkela_wire_10447;
    wire new_Jinkela_wire_9850;
    wire new_Jinkela_wire_5947;
    wire new_Jinkela_wire_7021;
    wire new_Jinkela_wire_2906;
    wire new_Jinkela_wire_4187;
    wire new_Jinkela_wire_9910;
    wire new_Jinkela_wire_7125;
    wire new_Jinkela_wire_7217;
    wire new_Jinkela_wire_9626;
    wire new_Jinkela_wire_3550;
    wire new_Jinkela_wire_4476;
    wire new_Jinkela_wire_2765;
    wire n_0493_;
    wire new_Jinkela_wire_7961;
    wire new_Jinkela_wire_10059;
    wire new_Jinkela_wire_6741;
    wire new_Jinkela_wire_1408;
    wire new_Jinkela_wire_3769;
    wire new_Jinkela_wire_8910;
    wire new_Jinkela_wire_7593;
    wire n_0788_;
    wire n_1291_;
    wire n_1331_;
    wire new_Jinkela_wire_9639;
    wire new_Jinkela_wire_1942;
    wire new_Jinkela_wire_6317;
    wire n_1238_;
    wire new_Jinkela_wire_33;
    wire new_Jinkela_wire_6512;
    wire new_Jinkela_wire_1700;
    wire new_Jinkela_wire_8976;
    wire new_Jinkela_wire_1286;
    wire n_1095_;
    wire new_Jinkela_wire_7942;
    wire new_Jinkela_wire_3864;
    wire new_Jinkela_wire_7962;
    wire n_0468_;
    wire new_net_2560;
    wire new_Jinkela_wire_9489;
    wire new_Jinkela_wire_10356;
    wire n_0474_;
    wire new_Jinkela_wire_223;
    wire new_Jinkela_wire_5396;
    wire new_Jinkela_wire_2080;
    wire new_Jinkela_wire_8503;
    wire new_Jinkela_wire_5885;
    wire new_Jinkela_wire_3406;
    wire new_Jinkela_wire_1150;
    wire new_Jinkela_wire_9451;
    wire new_Jinkela_wire_4030;
    wire new_Jinkela_wire_9024;
    wire n_0594_;
    wire new_Jinkela_wire_9998;
    wire new_Jinkela_wire_8261;
    wire new_Jinkela_wire_5354;
    wire new_Jinkela_wire_2882;
    wire new_Jinkela_wire_4398;
    wire new_Jinkela_wire_7958;
    wire new_Jinkela_wire_7929;
    wire new_Jinkela_wire_9506;
    wire new_Jinkela_wire_10566;
    wire new_Jinkela_wire_4968;
    wire new_Jinkela_wire_5371;
    wire new_Jinkela_wire_8336;
    wire new_Jinkela_wire_15;
    wire new_Jinkela_wire_2147;
    wire new_Jinkela_wire_4830;
    wire n_1206_;
    wire new_Jinkela_wire_3499;
    wire new_Jinkela_wire_6273;
    wire new_Jinkela_wire_3317;
    wire n_0977_;
    wire new_Jinkela_wire_2558;
    wire new_Jinkela_wire_4736;
    wire new_Jinkela_wire_8947;
    wire new_Jinkela_wire_5577;
    wire new_Jinkela_wire_262;
    wire new_Jinkela_wire_7423;
    wire new_Jinkela_wire_6301;
    wire new_Jinkela_wire_667;
    wire new_Jinkela_wire_2175;
    wire n_0695_;
    wire new_Jinkela_wire_9844;
    wire new_Jinkela_wire_6241;
    wire n_0719_;
    wire new_Jinkela_wire_5427;
    wire new_Jinkela_wire_639;
    wire new_Jinkela_wire_1864;
    wire new_Jinkela_wire_1622;
    wire n_0639_;
    wire n_0831_;
    wire new_Jinkela_wire_4779;
    wire n_0616_;
    wire new_Jinkela_wire_10400;
    wire new_Jinkela_wire_7398;
    wire new_Jinkela_wire_7585;
    wire new_Jinkela_wire_704;
    wire new_Jinkela_wire_6682;
    wire new_Jinkela_wire_6772;
    wire new_Jinkela_wire_3346;
    wire new_Jinkela_wire_3111;
    wire new_Jinkela_wire_9738;
    wire new_Jinkela_wire_5401;
    wire new_Jinkela_wire_1473;
    wire n_0492_;
    wire new_Jinkela_wire_7272;
    wire new_Jinkela_wire_6937;
    wire new_Jinkela_wire_9949;
    wire new_Jinkela_wire_5052;
    wire new_Jinkela_wire_3838;
    wire new_Jinkela_wire_6768;
    wire new_Jinkela_wire_42;
    wire new_Jinkela_wire_7390;
    wire new_Jinkela_wire_2780;
    wire n_0732_;
    wire new_Jinkela_wire_5364;
    wire new_Jinkela_wire_2065;
    wire new_Jinkela_wire_3389;
    wire n_1117_;
    wire new_Jinkela_wire_7212;
    wire new_Jinkela_wire_10362;
    wire new_Jinkela_wire_1866;
    wire new_Jinkela_wire_9060;
    wire new_Jinkela_wire_1797;
    wire new_Jinkela_wire_8448;
    wire new_Jinkela_wire_7379;
    wire n_1033_;
    wire new_Jinkela_wire_3976;
    wire new_Jinkela_wire_6387;
    wire new_Jinkela_wire_3906;
    wire new_Jinkela_wire_3673;
    wire new_Jinkela_wire_10015;
    wire new_Jinkela_wire_4180;
    wire new_Jinkela_wire_9239;
    wire new_Jinkela_wire_2969;
    wire new_Jinkela_wire_9359;
    wire n_0647_;
    wire new_Jinkela_wire_2506;
    wire new_Jinkela_wire_8238;
    wire new_Jinkela_wire_2420;
    wire new_Jinkela_wire_6198;
    wire new_Jinkela_wire_7198;
    wire new_Jinkela_wire_7683;
    wire new_Jinkela_wire_8186;
    wire new_Jinkela_wire_4477;
    wire new_Jinkela_wire_6311;
    wire new_Jinkela_wire_5933;
    wire new_Jinkela_wire_6369;
    wire new_Jinkela_wire_8022;
    wire new_Jinkela_wire_5767;
    wire new_Jinkela_wire_7195;
    wire new_Jinkela_wire_6821;
    wire new_Jinkela_wire_9885;
    wire new_Jinkela_wire_3683;
    wire new_Jinkela_wire_6159;
    wire new_Jinkela_wire_703;
    wire new_Jinkela_wire_1140;
    wire new_Jinkela_wire_2876;
    wire new_Jinkela_wire_9552;
    wire new_Jinkela_wire_10224;
    wire new_Jinkela_wire_4784;
    wire new_Jinkela_wire_9100;
    wire new_Jinkela_wire_1218;
    wire new_Jinkela_wire_8945;
    wire new_Jinkela_wire_4662;
    wire new_Jinkela_wire_5446;
    wire new_Jinkela_wire_6477;
    wire new_Jinkela_wire_2867;
    wire new_Jinkela_wire_5563;
    wire new_Jinkela_wire_9828;
    wire new_net_2501;
    wire new_Jinkela_wire_2018;
    wire n_1187_;
    wire new_Jinkela_wire_7952;
    wire n_1041_;
    wire new_Jinkela_wire_8245;
    wire new_Jinkela_wire_9333;
    wire n_0659_;
    wire n_1196_;
    wire new_Jinkela_wire_8392;
    wire new_Jinkela_wire_5622;
    wire new_Jinkela_wire_9709;
    wire new_Jinkela_wire_2131;
    wire new_Jinkela_wire_2697;
    wire new_Jinkela_wire_6758;
    wire new_Jinkela_wire_8044;
    wire new_Jinkela_wire_5789;
    wire new_Jinkela_wire_7265;
    wire new_Jinkela_wire_3978;
    wire new_Jinkela_wire_6849;
    wire new_Jinkela_wire_4153;
    wire new_Jinkela_wire_8831;
    wire new_Jinkela_wire_10485;
    wire n_0791_;
    wire new_Jinkela_wire_1395;
    wire n_0972_;
    wire new_Jinkela_wire_6638;
    wire new_Jinkela_wire_1203;
    wire new_Jinkela_wire_5096;
    wire new_Jinkela_wire_3657;
    wire new_Jinkela_wire_8492;
    wire new_Jinkela_wire_1548;
    wire new_Jinkela_wire_4556;
    wire new_Jinkela_wire_4485;
    wire new_Jinkela_wire_1466;
    wire new_Jinkela_wire_1805;
    wire new_Jinkela_wire_2735;
    wire new_Jinkela_wire_852;
    wire new_Jinkela_wire_8397;
    wire n_1351_;
    wire new_Jinkela_wire_9878;
    wire new_Jinkela_wire_6263;
    wire n_0339_;
    wire n_0768_;
    wire new_Jinkela_wire_3366;
    wire new_Jinkela_wire_8282;
    wire new_Jinkela_wire_3832;
    wire new_Jinkela_wire_2377;
    wire new_Jinkela_wire_7437;
    wire new_Jinkela_wire_3348;
    wire new_Jinkela_wire_4254;
    wire n_1190_;
    wire new_Jinkela_wire_10173;
    wire new_Jinkela_wire_4975;
    wire new_Jinkela_wire_6913;
    wire n_0213_;
    wire new_Jinkela_wire_1793;
    wire new_Jinkela_wire_6749;
    wire new_Jinkela_wire_123;
    wire new_Jinkela_wire_4379;
    wire new_Jinkela_wire_8364;
    wire new_Jinkela_wire_3994;
    wire new_Jinkela_wire_9023;
    wire new_Jinkela_wire_3108;
    wire new_Jinkela_wire_5120;
    wire new_Jinkela_wire_7449;
    wire new_Jinkela_wire_2931;
    wire n_0898_;
    wire new_Jinkela_wire_1177;
    wire new_Jinkela_wire_5362;
    wire new_Jinkela_wire_6596;
    wire new_Jinkela_wire_8651;
    wire new_Jinkela_wire_2853;
    wire new_Jinkela_wire_3950;
    wire n_0023_;
    wire new_Jinkela_wire_4906;
    wire new_Jinkela_wire_8988;
    wire new_Jinkela_wire_6912;
    wire new_Jinkela_wire_9545;
    wire new_Jinkela_wire_553;
    wire new_Jinkela_wire_8731;
    wire new_Jinkela_wire_7130;
    wire new_Jinkela_wire_10545;
    wire n_0175_;
    wire new_net_2576;
    wire new_Jinkela_wire_489;
    wire new_Jinkela_wire_6422;
    wire n_0957_;
    wire new_Jinkela_wire_2047;
    wire new_Jinkela_wire_8605;
    wire new_Jinkela_wire_6066;
    wire new_Jinkela_wire_3498;
    wire new_Jinkela_wire_5682;
    wire new_Jinkela_wire_2117;
    wire new_Jinkela_wire_7808;
    wire new_Jinkela_wire_5337;
    wire new_Jinkela_wire_2187;
    wire new_Jinkela_wire_2294;
    wire new_Jinkela_wire_10125;
    wire new_Jinkela_wire_5535;
    wire new_Jinkela_wire_3977;
    wire new_Jinkela_wire_1909;
    wire new_Jinkela_wire_6740;
    wire n_0819_;
    wire new_Jinkela_wire_4475;
    wire new_Jinkela_wire_8624;
    wire new_Jinkela_wire_5504;
    wire new_Jinkela_wire_9300;
    wire new_Jinkela_wire_3226;
    wire new_Jinkela_wire_3428;
    wire new_Jinkela_wire_8145;
    wire new_Jinkela_wire_6174;
    wire new_Jinkela_wire_894;
    wire new_Jinkela_wire_7812;
    wire new_Jinkela_wire_3007;
    wire new_Jinkela_wire_4354;
    wire new_Jinkela_wire_803;
    wire new_Jinkela_wire_5865;
    wire new_Jinkela_wire_1817;
    wire new_Jinkela_wire_4763;
    wire new_Jinkela_wire_7436;
    wire new_Jinkela_wire_6534;
    wire n_1188_;
    wire new_Jinkela_wire_9291;
    wire n_0736_;
    wire new_Jinkela_wire_9950;
    wire new_Jinkela_wire_8787;
    wire new_Jinkela_wire_2608;
    wire new_Jinkela_wire_5225;
    wire new_Jinkela_wire_652;
    wire new_Jinkela_wire_5300;
    wire new_Jinkela_wire_4488;
    wire new_Jinkela_wire_6791;
    wire new_Jinkela_wire_1125;
    wire new_Jinkela_wire_6073;
    wire new_Jinkela_wire_4478;
    wire new_Jinkela_wire_2897;
    wire new_Jinkela_wire_4858;
    wire new_Jinkela_wire_1816;
    wire new_Jinkela_wire_9375;
    wire new_Jinkela_wire_2153;
    wire new_Jinkela_wire_2942;
    wire new_Jinkela_wire_6730;
    wire new_Jinkela_wire_7204;
    wire new_Jinkela_wire_10139;
    wire new_Jinkela_wire_1614;
    wire new_Jinkela_wire_3962;
    wire new_Jinkela_wire_10435;
    wire n_0850_;
    wire new_Jinkela_wire_9725;
    wire new_Jinkela_wire_8505;
    wire new_Jinkela_wire_9769;
    wire new_Jinkela_wire_10045;
    wire new_Jinkela_wire_7536;
    wire new_Jinkela_wire_1243;
    wire new_Jinkela_wire_6381;
    wire new_Jinkela_wire_6135;
    wire new_Jinkela_wire_4096;
    wire new_Jinkela_wire_7765;
    wire new_Jinkela_wire_229;
    wire new_Jinkela_wire_4395;
    wire new_Jinkela_wire_1145;
    wire n_0725_;
    wire new_Jinkela_wire_7722;
    wire new_Jinkela_wire_2597;
    wire new_Jinkela_wire_1040;
    wire n_1077_;
    wire new_Jinkela_wire_2904;
    wire new_Jinkela_wire_2781;
    wire new_Jinkela_wire_1092;
    wire new_Jinkela_wire_4036;
    wire new_Jinkela_wire_8001;
    wire new_Jinkela_wire_10000;
    wire n_0182_;
    wire new_Jinkela_wire_7043;
    wire new_Jinkela_wire_10551;
    wire new_Jinkela_wire_6805;
    wire new_Jinkela_wire_7097;
    wire new_Jinkela_wire_2829;
    wire new_Jinkela_wire_8330;
    wire new_Jinkela_wire_8759;
    wire new_Jinkela_wire_43;
    wire new_Jinkela_wire_6825;
    wire n_0712_;
    wire new_Jinkela_wire_4435;
    wire new_Jinkela_wire_329;
    wire new_Jinkela_wire_3728;
    wire new_Jinkela_wire_3010;
    wire new_Jinkela_wire_10078;
    wire new_Jinkela_wire_618;
    wire new_Jinkela_wire_6153;
    wire new_Jinkela_wire_9685;
    wire new_Jinkela_wire_5395;
    wire new_Jinkela_wire_5693;
    wire new_Jinkela_wire_7552;
    wire n_1313_;
    wire new_Jinkela_wire_8481;
    wire new_Jinkela_wire_7196;
    wire new_Jinkela_wire_2787;
    wire new_Jinkela_wire_697;
    wire new_Jinkela_wire_8728;
    wire new_Jinkela_wire_4314;
    wire new_Jinkela_wire_2845;
    wire new_Jinkela_wire_3087;
    wire new_Jinkela_wire_6563;
    wire new_Jinkela_wire_2974;
    wire n_1302_;
    wire new_Jinkela_wire_6930;
    wire new_Jinkela_wire_1971;
    wire new_Jinkela_wire_8160;
    wire new_Jinkela_wire_1960;
    wire new_Jinkela_wire_9951;
    wire new_Jinkela_wire_2740;
    wire new_Jinkela_wire_3411;
    wire new_Jinkela_wire_5840;
    wire n_0503_;
    wire new_Jinkela_wire_6330;
    wire new_Jinkela_wire_2337;
    wire new_Jinkela_wire_6669;
    wire new_Jinkela_wire_1791;
    wire new_Jinkela_wire_7192;
    wire new_Jinkela_wire_1889;
    wire new_Jinkela_wire_3018;
    wire new_Jinkela_wire_8761;
    wire new_Jinkela_wire_3540;
    wire new_Jinkela_wire_7165;
    wire new_Jinkela_wire_2743;
    wire new_Jinkela_wire_837;
    wire new_Jinkela_wire_6472;
    wire new_Jinkela_wire_3843;
    wire new_Jinkela_wire_7533;
    wire new_Jinkela_wire_8618;
    wire new_Jinkela_wire_5604;
    wire new_Jinkela_wire_971;
    wire new_Jinkela_wire_8933;
    wire n_0548_;
    wire new_Jinkela_wire_1699;
    wire new_Jinkela_wire_3380;
    wire new_Jinkela_wire_9180;
    wire new_Jinkela_wire_8964;
    wire new_Jinkela_wire_938;
    wire new_Jinkela_wire_4467;
    wire new_Jinkela_wire_5847;
    wire new_Jinkela_wire_9970;
    wire new_Jinkela_wire_9843;
    wire new_Jinkela_wire_8305;
    wire new_Jinkela_wire_9590;
    wire new_Jinkela_wire_531;
    wire new_Jinkela_wire_130;
    wire new_Jinkela_wire_8676;
    wire new_Jinkela_wire_3649;
    wire new_Jinkela_wire_4884;
    wire new_Jinkela_wire_5082;
    wire new_Jinkela_wire_166;
    wire new_Jinkela_wire_3307;
    wire n_0475_;
    wire n_1357_;
    wire new_Jinkela_wire_6007;
    wire new_Jinkela_wire_9174;
    wire new_Jinkela_wire_1317;
    wire new_net_2572;
    wire new_Jinkela_wire_6289;
    wire new_Jinkela_wire_5875;
    wire new_Jinkela_wire_2539;
    wire new_Jinkela_wire_3816;
    wire new_Jinkela_wire_1800;
    wire new_Jinkela_wire_9085;
    wire n_0091_;
    wire new_Jinkela_wire_5804;
    wire new_Jinkela_wire_906;
    wire new_Jinkela_wire_4369;
    wire new_Jinkela_wire_8905;
    wire new_Jinkela_wire_7894;
    wire new_Jinkela_wire_480;
    wire new_Jinkela_wire_3619;
    wire new_Jinkela_wire_569;
    wire new_Jinkela_wire_6754;
    wire new_Jinkela_wire_1984;
    wire new_Jinkela_wire_53;
    wire new_Jinkela_wire_6467;
    wire new_Jinkela_wire_5704;
    wire new_Jinkela_wire_108;
    wire new_Jinkela_wire_7903;
    wire new_Jinkela_wire_4167;
    wire new_Jinkela_wire_8845;
    wire new_Jinkela_wire_1066;
    wire new_Jinkela_wire_5365;
    wire n_0145_;
    wire new_Jinkela_wire_145;
    wire new_Jinkela_wire_4470;
    wire new_Jinkela_wire_7301;
    wire new_Jinkela_wire_5972;
    wire new_Jinkela_wire_7135;
    wire new_Jinkela_wire_1893;
    wire new_Jinkela_wire_9047;
    wire new_Jinkela_wire_1883;
    wire new_Jinkela_wire_3990;
    wire new_Jinkela_wire_3425;
    wire new_Jinkela_wire_3206;
    wire n_0174_;
    wire new_Jinkela_wire_6685;
    wire new_Jinkela_wire_3082;
    wire new_Jinkela_wire_7556;
    wire new_Jinkela_wire_641;
    wire n_0039_;
    wire new_Jinkela_wire_4589;
    wire new_Jinkela_wire_3563;
    wire new_Jinkela_wire_4649;
    wire new_Jinkela_wire_9608;
    wire new_Jinkela_wire_6012;
    wire new_Jinkela_wire_2563;
    wire new_Jinkela_wire_6340;
    wire n_0431_;
    wire new_Jinkela_wire_1572;
    wire new_Jinkela_wire_5;
    wire new_Jinkela_wire_4469;
    wire new_Jinkela_wire_9334;
    wire new_Jinkela_wire_6458;
    wire new_Jinkela_wire_9371;
    wire n_0396_;
    wire new_Jinkela_wire_8527;
    wire new_Jinkela_wire_4228;
    wire new_Jinkela_wire_2999;
    wire new_Jinkela_wire_5432;
    wire new_Jinkela_wire_2416;
    wire new_Jinkela_wire_6376;
    wire new_Jinkela_wire_1418;
    wire new_Jinkela_wire_8215;
    wire new_Jinkela_wire_8485;
    wire new_Jinkela_wire_759;
    wire n_1031_;
    wire new_Jinkela_wire_8925;
    wire new_Jinkela_wire_2877;
    wire new_Jinkela_wire_227;
    wire new_Jinkela_wire_8249;
    wire new_Jinkela_wire_4350;
    wire new_Jinkela_wire_8662;
    wire new_Jinkela_wire_954;
    wire new_Jinkela_wire_1566;
    wire new_Jinkela_wire_6745;
    wire new_Jinkela_wire_5986;
    wire new_Jinkela_wire_555;
    wire new_Jinkela_wire_4684;
    wire n_1185_;
    wire new_Jinkela_wire_5189;
    wire new_Jinkela_wire_10322;
    wire n_1298_;
    wire new_Jinkela_wire_1916;
    wire new_Jinkela_wire_880;
    wire new_Jinkela_wire_4171;
    wire new_Jinkela_wire_4866;
    wire new_Jinkela_wire_216;
    wire new_Jinkela_wire_95;
    wire new_Jinkela_wire_1172;
    wire new_Jinkela_wire_634;
    wire new_Jinkela_wire_998;
    wire new_Jinkela_wire_3284;
    wire new_Jinkela_wire_5262;
    wire new_Jinkela_wire_3442;
    wire new_Jinkela_wire_8921;
    wire n_0862_;
    wire new_Jinkela_wire_3553;
    wire new_Jinkela_wire_3932;
    wire new_Jinkela_wire_168;
    wire new_Jinkela_wire_3985;
    wire new_Jinkela_wire_1626;
    wire new_Jinkela_wire_9028;
    wire new_Jinkela_wire_1446;
    wire new_Jinkela_wire_3210;
    wire new_Jinkela_wire_646;
    wire new_Jinkela_wire_9109;
    wire new_Jinkela_wire_4715;
    wire new_Jinkela_wire_7987;
    wire new_Jinkela_wire_8250;
    wire new_Jinkela_wire_6921;
    wire new_Jinkela_wire_1631;
    wire n_0336_;
    wire n_0315_;
    wire new_Jinkela_wire_2744;
    wire new_Jinkela_wire_6243;
    wire new_Jinkela_wire_7105;
    wire new_Jinkela_wire_6457;
    wire new_Jinkela_wire_610;
    wire new_Jinkela_wire_2733;
    wire new_Jinkela_wire_6909;
    wire new_Jinkela_wire_2578;
    wire new_Jinkela_wire_6069;
    wire new_Jinkela_wire_10611;
    wire new_Jinkela_wire_1870;
    wire new_Jinkela_wire_6751;
    wire new_Jinkela_wire_5922;
    wire new_Jinkela_wire_220;
    wire n_0279_;
    wire new_Jinkela_wire_5977;
    wire new_Jinkela_wire_8669;
    wire new_Jinkela_wire_8530;
    wire new_Jinkela_wire_8082;
    wire n_1040_;
    wire new_Jinkela_wire_5590;
    wire new_Jinkela_wire_3679;
    wire new_Jinkela_wire_3331;
    wire new_Jinkela_wire_5681;
    wire new_Jinkela_wire_2090;
    wire new_Jinkela_wire_1114;
    wire new_Jinkela_wire_5750;
    wire new_Jinkela_wire_6295;
    wire new_Jinkela_wire_4119;
    wire new_Jinkela_wire_3625;
    wire new_Jinkela_wire_7197;
    wire new_Jinkela_wire_10247;
    wire new_Jinkela_wire_10502;
    wire new_Jinkela_wire_4626;
    wire new_Jinkela_wire_698;
    wire new_Jinkela_wire_6782;
    wire new_Jinkela_wire_6500;
    wire new_Jinkela_wire_6944;
    wire new_Jinkela_wire_3974;
    wire new_Jinkela_wire_9937;
    wire new_Jinkela_wire_801;
    wire new_Jinkela_wire_1299;
    wire new_Jinkela_wire_10088;
    wire new_Jinkela_wire_5957;
    wire new_Jinkela_wire_6586;
    wire new_Jinkela_wire_3241;
    wire new_Jinkela_wire_8948;
    wire new_Jinkela_wire_8325;
    wire new_Jinkela_wire_7049;
    wire new_Jinkela_wire_9989;
    wire new_Jinkela_wire_5728;
    wire new_Jinkela_wire_2320;
    wire new_Jinkela_wire_7451;
    wire new_Jinkela_wire_3394;
    wire n_1182_;
    wire new_Jinkela_wire_6987;
    wire new_Jinkela_wire_4898;
    wire new_Jinkela_wire_9020;
    wire new_Jinkela_wire_10004;
    wire new_Jinkela_wire_3311;
    wire new_Jinkela_wire_6559;
    wire new_Jinkela_wire_3417;
    wire new_Jinkela_wire_7069;
    wire new_Jinkela_wire_9175;
    wire new_Jinkela_wire_5915;
    wire new_Jinkela_wire_8144;
    wire new_net_2515;
    wire n_0727_;
    wire n_0970_;
    wire new_Jinkela_wire_883;
    wire new_Jinkela_wire_1612;
    wire new_Jinkela_wire_7439;
    wire new_Jinkela_wire_904;
    wire new_Jinkela_wire_8920;
    wire new_Jinkela_wire_4206;
    wire new_Jinkela_wire_4878;
    wire new_Jinkela_wire_5013;
    wire new_Jinkela_wire_8693;
    wire n_0239_;
    wire new_Jinkela_wire_2604;
    wire new_Jinkela_wire_8923;
    wire new_Jinkela_wire_1704;
    wire new_Jinkela_wire_7428;
    wire n_0001_;
    wire new_Jinkela_wire_9599;
    wire new_Jinkela_wire_6834;
    wire new_Jinkela_wire_82;
    wire new_Jinkela_wire_4778;
    wire n_0655_;
    wire new_Jinkela_wire_4995;
    wire new_Jinkela_wire_1568;
    wire new_Jinkela_wire_2500;
    wire new_Jinkela_wire_6523;
    wire n_0757_;
    wire new_Jinkela_wire_4753;
    wire new_Jinkela_wire_592;
    wire new_Jinkela_wire_5311;
    wire new_Jinkela_wire_343;
    wire n_0309_;
    wire new_Jinkela_wire_1640;
    wire new_Jinkela_wire_8326;
    wire new_Jinkela_wire_137;
    wire new_Jinkela_wire_7904;
    wire new_Jinkela_wire_4988;
    wire new_Jinkela_wire_2706;
    wire new_Jinkela_wire_5429;
    wire new_Jinkela_wire_1428;
    wire new_Jinkela_wire_1755;
    wire new_Jinkela_wire_3905;
    wire new_Jinkela_wire_3813;
    wire new_Jinkela_wire_9658;
    wire new_Jinkela_wire_6318;
    wire new_Jinkela_wire_7207;
    wire new_Jinkela_wire_5316;
    wire new_Jinkela_wire_9710;
    wire new_Jinkela_wire_8285;
    wire new_Jinkela_wire_1175;
    wire new_Jinkela_wire_6019;
    wire new_Jinkela_wire_2924;
    wire new_Jinkela_wire_10467;
    wire new_Jinkela_wire_7652;
    wire new_Jinkela_wire_10249;
    wire new_Jinkela_wire_179;
    wire n_1065_;
    wire new_Jinkela_wire_4211;
    wire new_Jinkela_wire_8718;
    wire new_Jinkela_wire_4558;
    wire new_Jinkela_wire_9422;
    wire new_Jinkela_wire_3666;
    wire new_Jinkela_wire_2098;
    wire new_Jinkela_wire_5559;
    wire new_Jinkela_wire_586;
    wire new_Jinkela_wire_8216;
    wire new_Jinkela_wire_6608;
    wire new_Jinkela_wire_1741;
    wire new_Jinkela_wire_5103;
    wire new_Jinkela_wire_4092;
    wire new_Jinkela_wire_7160;
    wire n_0914_;
    wire new_Jinkela_wire_9689;
    wire new_Jinkela_wire_10213;
    wire new_Jinkela_wire_1765;
    wire new_Jinkela_wire_2528;
    wire new_Jinkela_wire_6804;
    wire new_Jinkela_wire_3227;
    wire n_0988_;
    wire new_Jinkela_wire_1135;
    wire new_Jinkela_wire_7798;
    wire new_Jinkela_wire_9537;
    wire new_Jinkela_wire_7663;
    wire new_Jinkela_wire_5064;
    wire new_Jinkela_wire_8375;
    wire new_Jinkela_wire_7126;
    wire new_Jinkela_wire_7278;
    wire n_0674_;
    wire new_Jinkela_wire_2314;
    wire new_Jinkela_wire_5757;
    wire n_0960_;
    wire new_Jinkela_wire_7028;
    wire new_Jinkela_wire_9208;
    wire new_Jinkela_wire_6419;
    wire new_Jinkela_wire_1573;
    wire n_0484_;
    wire n_0612_;
    wire new_Jinkela_wire_1542;
    wire new_Jinkela_wire_9413;
    wire n_0156_;
    wire new_Jinkela_wire_591;
    wire new_Jinkela_wire_8067;
    wire n_0784_;
    wire new_Jinkela_wire_2114;
    wire new_Jinkela_wire_2038;
    wire n_0417_;
    wire new_Jinkela_wire_961;
    wire new_Jinkela_wire_4802;
    wire new_Jinkela_wire_3839;
    wire new_Jinkela_wire_5815;
    wire new_Jinkela_wire_9513;
    wire new_Jinkela_wire_10426;
    wire new_Jinkela_wire_4729;
    wire new_Jinkela_wire_1912;
    wire new_Jinkela_wire_6659;
    wire new_Jinkela_wire_7517;
    wire new_Jinkela_wire_10484;
    wire new_Jinkela_wire_1343;
    wire new_Jinkela_wire_2017;
    wire n_1215_;
    wire new_Jinkela_wire_7950;
    wire new_Jinkela_wire_8432;
    wire new_Jinkela_wire_3143;
    wire new_Jinkela_wire_1020;
    wire new_Jinkela_wire_6160;
    wire new_Jinkela_wire_8868;
    wire new_Jinkela_wire_2494;
    wire new_Jinkela_wire_74;
    wire new_Jinkela_wire_10121;
    wire new_Jinkela_wire_9757;
    wire new_Jinkela_wire_5791;
    wire new_Jinkela_wire_6345;
    wire new_Jinkela_wire_7239;
    wire new_Jinkela_wire_2818;
    wire new_Jinkela_wire_6212;
    wire n_0333_;
    wire new_Jinkela_wire_9205;
    wire new_Jinkela_wire_1443;
    wire new_Jinkela_wire_1421;
    wire n_1284_;
    wire new_Jinkela_wire_4182;
    wire new_Jinkela_wire_3272;
    wire n_0040_;
    wire new_Jinkela_wire_2185;
    wire n_0228_;
    wire new_Jinkela_wire_1977;
    wire new_Jinkela_wire_8315;
    wire new_Jinkela_wire_8675;
    wire n_0829_;
    wire new_Jinkela_wire_7813;
    wire new_Jinkela_wire_6907;
    wire new_Jinkela_wire_1205;
    wire new_Jinkela_wire_8252;
    wire new_Jinkela_wire_7271;
    wire new_Jinkela_wire_9121;
    wire new_Jinkela_wire_8077;
    wire new_Jinkela_wire_9830;
    wire new_Jinkela_wire_963;
    wire new_Jinkela_wire_1014;
    wire new_Jinkela_wire_7489;
    wire new_Jinkela_wire_8773;
    wire n_0030_;
    wire n_0264_;
    wire new_Jinkela_wire_413;
    wire new_Jinkela_wire_4563;
    wire n_0242_;
    wire new_Jinkela_wire_4519;
    wire new_Jinkela_wire_8581;
    wire new_Jinkela_wire_6629;
    wire new_Jinkela_wire_9332;
    wire n_1301_;
    wire new_Jinkela_wire_9113;
    wire new_Jinkela_wire_1799;
    wire new_Jinkela_wire_297;
    wire new_Jinkela_wire_3586;
    wire new_Jinkela_wire_5652;
    wire new_Jinkela_wire_7409;
    wire new_Jinkela_wire_7679;
    wire n_0247_;
    wire new_Jinkela_wire_6481;
    wire new_Jinkela_wire_9908;
    wire new_Jinkela_wire_5088;
    wire new_Jinkela_wire_5525;
    wire n_0280_;
    wire new_Jinkela_wire_8573;
    wire new_Jinkela_wire_9251;
    wire new_Jinkela_wire_6057;
    wire new_Jinkela_wire_4994;
    wire new_Jinkela_wire_2390;
    wire new_Jinkela_wire_4606;
    wire new_Jinkela_wire_2826;
    wire new_Jinkela_wire_10550;
    wire new_Jinkela_wire_5471;
    wire new_Jinkela_wire_5036;
    wire new_Jinkela_wire_1646;
    wire new_Jinkela_wire_9176;
    wire new_Jinkela_wire_142;
    wire new_Jinkela_wire_10399;
    wire new_Jinkela_wire_6305;
    wire n_1270_;
    wire new_Jinkela_wire_3698;
    wire new_Jinkela_wire_5579;
    wire new_Jinkela_wire_6521;
    wire new_Jinkela_wire_7915;
    wire n_0405_;
    wire new_Jinkela_wire_5322;
    wire new_Jinkela_wire_3732;
    wire new_Jinkela_wire_3237;
    wire new_Jinkela_wire_6974;
    wire new_Jinkela_wire_4647;
    wire new_Jinkela_wire_3339;
    wire new_Jinkela_wire_1758;
    wire new_Jinkela_wire_1610;
    wire new_Jinkela_wire_388;
    wire new_Jinkela_wire_9045;
    wire new_Jinkela_wire_8081;
    wire new_Jinkela_wire_1434;
    wire new_Jinkela_wire_7814;
    wire new_Jinkela_wire_354;
    wire new_Jinkela_wire_7917;
    wire n_0038_;
    wire new_Jinkela_wire_8092;
    wire n_0684_;
    wire new_Jinkela_wire_2383;
    wire new_Jinkela_wire_4012;
    wire new_Jinkela_wire_3562;
    wire new_Jinkela_wire_1918;
    wire new_Jinkela_wire_8667;
    wire new_Jinkela_wire_6199;
    wire new_Jinkela_wire_5330;
    wire new_Jinkela_wire_4535;
    wire new_Jinkela_wire_3859;
    wire n_1122_;
    wire new_Jinkela_wire_9679;
    wire new_Jinkela_wire_5902;
    wire new_Jinkela_wire_305;
    wire n_1193_;
    wire new_Jinkela_wire_1086;
    wire n_1203_;
    wire new_Jinkela_wire_1109;
    wire new_Jinkela_wire_151;
    wire new_Jinkela_wire_7544;
    wire new_Jinkela_wire_1709;
    wire new_Jinkela_wire_5723;
    wire new_Jinkela_wire_4446;
    wire new_Jinkela_wire_9026;
    wire new_Jinkela_wire_2580;
    wire new_Jinkela_wire_2431;
    wire new_Jinkela_wire_2615;
    wire new_Jinkela_wire_3809;
    wire new_Jinkela_wire_2678;
    wire n_0473_;
    wire new_Jinkela_wire_2368;
    wire new_Jinkela_wire_4727;
    wire new_Jinkela_wire_9941;
    wire new_Jinkela_wire_1813;
    wire new_Jinkela_wire_9290;
    wire new_Jinkela_wire_3520;
    wire new_Jinkela_wire_7840;
    wire new_Jinkela_wire_3290;
    wire new_Jinkela_wire_10573;
    wire new_Jinkela_wire_2532;
    wire new_Jinkela_wire_8143;
    wire new_Jinkela_wire_8510;
    wire new_Jinkela_wire_1940;
    wire new_Jinkela_wire_6490;
    wire new_Jinkela_wire_1108;
    wire new_Jinkela_wire_3610;
    wire new_Jinkela_wire_3548;
    wire new_Jinkela_wire_2881;
    wire new_Jinkela_wire_10106;
    wire new_Jinkela_wire_5335;
    wire new_Jinkela_wire_3001;
    wire new_Jinkela_wire_4963;
    wire new_Jinkela_wire_2208;
    wire new_Jinkela_wire_2947;
    wire n_0827_;
    wire new_Jinkela_wire_6902;
    wire new_Jinkela_wire_1312;
    wire n_0360_;
    wire new_Jinkela_wire_1978;
    wire new_Jinkela_wire_8961;
    wire new_Jinkela_wire_9153;
    wire new_Jinkela_wire_7644;
    wire new_Jinkela_wire_8300;
    wire new_Jinkela_wire_7782;
    wire new_Jinkela_wire_9178;
    wire n_0132_;
    wire new_Jinkela_wire_9519;
    wire new_Jinkela_wire_5720;
    wire new_Jinkela_wire_9499;
    wire new_Jinkela_wire_1992;
    wire new_Jinkela_wire_2496;
    wire new_Jinkela_wire_4737;
    wire new_Jinkela_wire_967;
    wire new_Jinkela_wire_2940;
    wire new_Jinkela_wire_7540;
    wire new_Jinkela_wire_2739;
    wire n_1133_;
    wire new_Jinkela_wire_2084;
    wire new_Jinkela_wire_7032;
    wire new_Jinkela_wire_9084;
    wire new_Jinkela_wire_5828;
    wire new_Jinkela_wire_6297;
    wire n_0016_;
    wire n_1123_;
    wire n_1341_;
    wire n_0606_;
    wire new_Jinkela_wire_8423;
    wire new_Jinkela_wire_4424;
    wire new_Jinkela_wire_9919;
    wire new_Jinkela_wire_2475;
    wire new_Jinkela_wire_9318;
    wire new_Jinkela_wire_7223;
    wire n_0289_;
    wire new_Jinkela_wire_2619;
    wire new_Jinkela_wire_7146;
    wire new_Jinkela_wire_419;
    wire new_Jinkela_wire_327;
    wire new_Jinkela_wire_4234;
    wire new_Jinkela_wire_7394;
    wire new_Jinkela_wire_10340;
    wire new_Jinkela_wire_1047;
    wire new_Jinkela_wire_6339;
    wire new_Jinkela_wire_10289;
    wire new_Jinkela_wire_403;
    wire new_Jinkela_wire_78;
    wire new_Jinkela_wire_3107;
    wire new_Jinkela_wire_9587;
    wire new_Jinkela_wire_10167;
    wire new_Jinkela_wire_2918;
    wire new_Jinkela_wire_10055;
    wire new_Jinkela_wire_6627;
    wire n_0231_;
    wire n_1046_;
    wire new_Jinkela_wire_5007;
    wire new_Jinkela_wire_3246;
    wire new_Jinkela_wire_1840;
    wire new_Jinkela_wire_1973;
    wire n_1022_;
    wire new_Jinkela_wire_1154;
    wire new_Jinkela_wire_8465;
    wire new_Jinkela_wire_1855;
    wire new_Jinkela_wire_5422;
    wire new_Jinkela_wire_6009;
    wire n_0153_;
    wire new_Jinkela_wire_2101;
    wire new_Jinkela_wire_6028;
    wire new_Jinkela_wire_5502;
    wire new_Jinkela_wire_9952;
    wire new_Jinkela_wire_2925;
    wire new_Jinkela_wire_7283;
    wire new_Jinkela_wire_8188;
    wire new_Jinkela_wire_5458;
    wire new_Jinkela_wire_434;
    wire new_Jinkela_wire_4713;
    wire n_1051_;
    wire new_Jinkela_wire_4357;
    wire new_Jinkela_wire_6168;
    wire new_Jinkela_wire_9149;
    wire new_Jinkela_wire_8401;
    wire new_Jinkela_wire_5870;
    wire new_Jinkela_wire_90;
    wire new_Jinkela_wire_1306;
    wire new_Jinkela_wire_6947;
    wire new_Jinkela_wire_1925;
    wire new_Jinkela_wire_8218;
    wire new_Jinkela_wire_3450;
    wire new_Jinkela_wire_3802;
    wire new_Jinkela_wire_1684;
    wire new_Jinkela_wire_2540;
    wire new_Jinkela_wire_4585;
    wire new_Jinkela_wire_7132;
    wire new_Jinkela_wire_6102;
    wire new_Jinkela_wire_2214;
    wire new_Jinkela_wire_2266;
    wire new_Jinkela_wire_7732;
    wire new_Jinkela_wire_4047;
    wire new_Jinkela_wire_10366;
    wire new_Jinkela_wire_2322;
    wire new_Jinkela_wire_9344;
    wire new_Jinkela_wire_7703;
    wire new_Jinkela_wire_1235;
    wire new_Jinkela_wire_3928;
    wire new_Jinkela_wire_743;
    wire new_Jinkela_wire_7429;
    wire new_Jinkela_wire_4847;
    wire new_Jinkela_wire_3573;
    wire new_Jinkela_wire_1049;
    wire new_Jinkela_wire_5603;
    wire new_Jinkela_wire_7567;
    wire new_Jinkela_wire_8986;
    wire new_Jinkela_wire_5246;
    wire new_Jinkela_wire_565;
    wire new_Jinkela_wire_6287;
    wire new_Jinkela_wire_2139;
    wire new_Jinkela_wire_331;
    wire new_Jinkela_wire_8740;
    wire new_Jinkela_wire_9816;
    wire new_Jinkela_wire_1139;
    wire n_0013_;
    wire n_0046_;
    wire n_0413_;
    wire n_1138_;
    wire new_Jinkela_wire_3303;
    wire new_Jinkela_wire_2165;
    wire new_Jinkela_wire_1352;
    wire new_Jinkela_wire_8244;
    wire new_Jinkela_wire_6879;
    wire new_Jinkela_wire_396;
    wire new_Jinkela_wire_2477;
    wire new_Jinkela_wire_4081;
    wire new_Jinkela_wire_5841;
    wire new_Jinkela_wire_2125;
    wire new_Jinkela_wire_8840;
    wire n_0652_;
    wire n_1242_;
    wire new_Jinkela_wire_4419;
    wire new_Jinkela_wire_9758;
    wire new_Jinkela_wire_8388;
    wire new_Jinkela_wire_3194;
    wire new_Jinkela_wire_1644;
    wire new_Jinkela_wire_3783;
    wire n_0723_;
    wire new_Jinkela_wire_4693;
    wire n_0702_;
    wire new_Jinkela_wire_8211;
    wire new_Jinkela_wire_8512;
    wire new_Jinkela_wire_2008;
    wire new_Jinkela_wire_7168;
    wire new_Jinkela_wire_548;
    wire n_0590_;
    wire new_Jinkela_wire_6567;
    wire new_Jinkela_wire_769;
    wire new_Jinkela_wire_1028;
    wire new_Jinkela_wire_6592;
    wire n_0251_;
    wire new_Jinkela_wire_8937;
    wire n_1365_;
    wire new_Jinkela_wire_4185;
    wire n_1092_;
    wire new_Jinkela_wire_991;
    wire new_Jinkela_wire_534;
    wire new_Jinkela_wire_4472;
    wire new_Jinkela_wire_9345;
    wire n_0162_;
    wire new_Jinkela_wire_411;
    wire new_Jinkela_wire_2872;
    wire new_Jinkela_wire_645;
    wire new_Jinkela_wire_8755;
    wire new_Jinkela_wire_4992;
    wire new_Jinkela_wire_6076;
    wire new_Jinkela_wire_6918;
    wire new_Jinkela_wire_8817;
    wire new_Jinkela_wire_8690;
    wire new_Jinkela_wire_1134;
    wire new_Jinkela_wire_247;
    wire new_Jinkela_wire_2675;
    wire new_Jinkela_wire_4601;
    wire new_Jinkela_wire_1924;
    wire new_Jinkela_wire_10332;
    wire new_Jinkela_wire_5566;
    wire new_Jinkela_wire_6479;
    wire n_0352_;
    wire new_Jinkela_wire_4877;
    wire new_Jinkela_wire_3655;
    wire new_Jinkela_wire_8223;
    wire new_Jinkela_wire_8642;
    wire new_Jinkela_wire_7569;
    wire new_Jinkela_wire_8424;
    wire new_Jinkela_wire_9362;
    wire new_Jinkela_wire_2834;
    wire new_Jinkela_wire_4874;
    wire new_Jinkela_wire_9140;
    wire new_Jinkela_wire_1877;
    wire new_Jinkela_wire_482;
    wire new_Jinkela_wire_8000;
    wire new_Jinkela_wire_7673;
    wire n_0526_;
    wire new_Jinkela_wire_4530;
    wire new_Jinkela_wire_9421;
    wire new_Jinkela_wire_6010;
    wire new_Jinkela_wire_1432;
    wire new_Jinkela_wire_9666;
    wire new_Jinkela_wire_10218;
    wire new_Jinkela_wire_5583;
    wire new_Jinkela_wire_7289;
    wire new_Jinkela_wire_1401;
    wire new_Jinkela_wire_8786;
    wire new_Jinkela_wire_2617;
    wire new_Jinkela_wire_9335;
    wire new_Jinkela_wire_93;
    wire new_Jinkela_wire_7749;
    wire new_Jinkela_wire_9984;
    wire new_Jinkela_wire_3938;
    wire new_Jinkela_wire_6778;
    wire n_0368_;
    wire new_Jinkela_wire_4418;
    wire new_Jinkela_wire_5778;
    wire new_Jinkela_wire_2636;
    wire new_Jinkela_wire_5496;
    wire new_Jinkela_wire_8084;
    wire new_Jinkela_wire_61;
    wire new_Jinkela_wire_3546;
    wire new_Jinkela_wire_5866;
    wire new_Jinkela_wire_9283;
    wire n_0774_;
    wire new_Jinkela_wire_1619;
    wire new_Jinkela_wire_4586;
    wire new_Jinkela_wire_2910;
    wire n_0539_;
    wire new_Jinkela_wire_5650;
    wire new_Jinkela_wire_9330;
    wire new_Jinkela_wire_8488;
    wire new_Jinkela_wire_6332;
    wire n_0176_;
    wire new_Jinkela_wire_7047;
    wire new_Jinkela_wire_9030;
    wire new_Jinkela_wire_8056;
    wire n_1363_;
    wire new_Jinkela_wire_1083;
    wire new_Jinkela_wire_5135;
    wire new_Jinkela_wire_5295;
    wire new_Jinkela_wire_6304;
    wire new_Jinkela_wire_5089;
    wire new_Jinkela_wire_6561;
    wire new_Jinkela_wire_8288;
    wire new_Jinkela_wire_10475;
    wire new_Jinkela_wire_4694;
    wire new_Jinkela_wire_4007;
    wire new_Jinkela_wire_8196;
    wire new_Jinkela_wire_4860;
    wire new_Jinkela_wire_5280;
    wire new_Jinkela_wire_3469;
    wire new_Jinkela_wire_3124;
    wire new_Jinkela_wire_1411;
    wire new_Jinkela_wire_7081;
    wire new_Jinkela_wire_9135;
    wire new_Jinkela_wire_8534;
    wire new_Jinkela_wire_9363;
    wire new_Jinkela_wire_6362;
    wire new_Jinkela_wire_5635;
    wire new_Jinkela_wire_7774;
    wire new_net_2489;
    wire new_Jinkela_wire_4498;
    wire new_Jinkela_wire_6571;
    wire new_Jinkela_wire_7764;
    wire n_0113_;
    wire new_Jinkela_wire_8438;
    wire new_Jinkela_wire_5992;
    wire new_Jinkela_wire_5117;
    wire new_Jinkela_wire_9312;
    wire n_0604_;
    wire new_Jinkela_wire_7062;
    wire new_Jinkela_wire_10123;
    wire new_Jinkela_wire_447;
    wire new_Jinkela_wire_7993;
    wire new_Jinkela_wire_3017;
    wire new_Jinkela_wire_3188;
    wire new_Jinkela_wire_6169;
    wire new_Jinkela_wire_9540;
    wire new_Jinkela_wire_9129;
    wire new_Jinkela_wire_7948;
    wire new_Jinkela_wire_2227;
    wire new_Jinkela_wire_514;
    wire n_1169_;
    wire new_Jinkela_wire_8893;
    wire new_Jinkela_wire_4217;
    wire new_Jinkela_wire_4974;
    wire new_Jinkela_wire_4690;
    wire new_Jinkela_wire_10448;
    wire n_0349_;
    wire n_0507_;
    wire new_Jinkela_wire_5712;
    wire new_Jinkela_wire_3309;
    wire new_Jinkela_wire_3444;
    wire new_Jinkela_wire_7723;
    wire new_Jinkela_wire_8585;
    wire new_Jinkela_wire_4105;
    wire new_Jinkela_wire_3102;
    wire new_Jinkela_wire_4335;
    wire new_Jinkela_wire_10251;
    wire new_Jinkela_wire_4954;
    wire new_Jinkela_wire_10005;
    wire new_Jinkela_wire_5562;
    wire new_Jinkela_wire_5062;
    wire new_Jinkela_wire_10051;
    wire new_Jinkela_wire_3256;
    wire new_Jinkela_wire_7244;
    wire new_Jinkela_wire_5093;
    wire n_0438_;
    wire new_Jinkela_wire_632;
    wire new_Jinkela_wire_799;
    wire new_Jinkela_wire_5158;
    wire new_Jinkela_wire_5308;
    wire new_Jinkela_wire_4943;
    wire new_Jinkela_wire_8563;
    wire new_Jinkela_wire_8399;
    wire new_Jinkela_wire_10554;
    wire new_Jinkela_wire_8449;
    wire new_Jinkela_wire_4422;
    wire new_Jinkela_wire_3088;
    wire new_Jinkela_wire_9539;
    wire new_Jinkela_wire_3729;
    wire new_Jinkela_wire_2657;
    wire new_Jinkela_wire_3847;
    wire n_0782_;
    wire new_Jinkela_wire_4594;
    wire new_Jinkela_wire_3743;
    wire new_Jinkela_wire_5313;
    wire new_Jinkela_wire_4427;
    wire new_Jinkela_wire_10194;
    wire new_Jinkela_wire_3245;
    wire new_Jinkela_wire_6284;
    wire new_Jinkela_wire_2859;
    wire n_0461_;
    wire new_Jinkela_wire_2210;
    wire new_Jinkela_wire_7361;
    wire n_1163_;
    wire new_Jinkela_wire_88;
    wire new_Jinkela_wire_6281;
    wire new_Jinkela_wire_1762;
    wire new_Jinkela_wire_4259;
    wire new_Jinkela_wire_4198;
    wire new_Jinkela_wire_5272;
    wire new_Jinkela_wire_6781;
    wire new_Jinkela_wire_7806;
    wire new_Jinkela_wire_6450;
    wire new_Jinkela_wire_8671;
    wire new_Jinkela_wire_9892;
    wire new_Jinkela_wire_10022;
    wire new_Jinkela_wire_9974;
    wire new_Jinkela_wire_10577;
    wire new_Jinkela_wire_1691;
    wire new_Jinkela_wire_8225;
    wire n_0418_;
    wire new_Jinkela_wire_7601;
    wire new_Jinkela_wire_426;
    wire new_Jinkela_wire_7460;
    wire new_Jinkela_wire_3522;
    wire n_1045_;
    wire new_Jinkela_wire_3874;
    wire new_Jinkela_wire_5180;
    wire new_Jinkela_wire_802;
    wire new_Jinkela_wire_3804;
    wire new_Jinkela_wire_3118;
    wire n_1276_;
    wire new_Jinkela_wire_8385;
    wire new_Jinkela_wire_795;
    wire new_Jinkela_wire_8865;
    wire n_1070_;
    wire new_Jinkela_wire_3566;
    wire new_Jinkela_wire_2109;
    wire new_Jinkela_wire_4214;
    wire new_Jinkela_wire_1304;
    wire n_0811_;
    wire new_Jinkela_wire_4745;
    wire new_Jinkela_wire_8452;
    wire new_Jinkela_wire_9099;
    wire new_Jinkela_wire_4448;
    wire new_Jinkela_wire_2029;
    wire new_Jinkela_wire_3952;
    wire new_Jinkela_wire_1493;
    wire n_0630_;
    wire new_Jinkela_wire_7308;
    wire new_Jinkela_wire_5056;
    wire new_Jinkela_wire_3222;
    wire n_0253_;
    wire new_Jinkela_wire_9007;
    wire new_Jinkela_wire_3234;
    wire new_Jinkela_wire_7476;
    wire new_Jinkela_wire_382;
    wire new_Jinkela_wire_1196;
    wire new_Jinkela_wire_8172;
    wire new_Jinkela_wire_3632;
    wire new_Jinkela_wire_4552;
    wire new_Jinkela_wire_7582;
    wire new_Jinkela_wire_5898;
    wire new_Jinkela_wire_1725;
    wire new_Jinkela_wire_9395;
    wire new_Jinkela_wire_8978;
    wire new_Jinkela_wire_3448;
    wire n_0935_;
    wire n_0785_;
    wire new_Jinkela_wire_7123;
    wire new_Jinkela_wire_6593;
    wire new_Jinkela_wire_10279;
    wire new_Jinkela_wire_7734;
    wire new_Jinkela_wire_955;
    wire new_Jinkela_wire_9956;
    wire new_Jinkela_wire_8430;
    wire new_Jinkela_wire_7358;
    wire new_Jinkela_wire_10518;
    wire new_Jinkela_wire_10082;
    wire new_Jinkela_wire_2298;
    wire new_Jinkela_wire_10096;
    wire new_Jinkela_wire_9981;
    wire new_Jinkela_wire_3106;
    wire new_Jinkela_wire_7352;
    wire n_1075_;
    wire new_Jinkela_wire_6686;
    wire new_Jinkela_wire_6461;
    wire new_Jinkela_wire_5136;
    wire n_1017_;
    wire new_Jinkela_wire_2460;
    wire new_Jinkela_wire_3564;
    wire new_Jinkela_wire_3567;
    wire new_Jinkela_wire_5257;
    wire new_Jinkela_wire_3399;
    wire new_Jinkela_wire_9826;
    wire new_Jinkela_wire_4580;
    wire n_0190_;
    wire new_Jinkela_wire_7743;
    wire new_Jinkela_wire_8998;
    wire new_Jinkela_wire_10292;
    wire new_Jinkela_wire_8985;
    wire new_Jinkela_wire_8233;
    wire new_Jinkela_wire_2864;
    wire new_Jinkela_wire_5184;
    wire new_Jinkela_wire_2273;
    wire new_Jinkela_wire_5861;
    wire new_Jinkela_wire_9555;
    wire new_Jinkela_wire_9789;
    wire new_Jinkela_wire_7686;
    wire new_Jinkela_wire_5950;
    wire new_Jinkela_wire_5323;
    wire new_Jinkela_wire_3236;
    wire new_Jinkela_wire_3293;
    wire new_Jinkela_wire_6617;
    wire new_Jinkela_wire_2079;
    wire new_Jinkela_wire_4324;
    wire new_Jinkela_wire_8795;
    wire new_Jinkela_wire_9156;
    wire new_Jinkela_wire_7637;
    wire new_Jinkela_wire_779;
    wire new_Jinkela_wire_5634;
    wire new_Jinkela_wire_8153;
    wire n_0044_;
    wire n_1345_;
    wire new_Jinkela_wire_353;
    wire new_Jinkela_wire_8628;
    wire new_Jinkela_wire_3963;
    wire new_Jinkela_wire_562;
    wire n_1131_;
    wire new_Jinkela_wire_8562;
    wire new_Jinkela_wire_1200;
    wire new_Jinkela_wire_1071;
    wire n_0971_;
    wire new_Jinkela_wire_9744;
    wire new_Jinkela_wire_2961;
    wire new_Jinkela_wire_5753;
    wire new_Jinkela_wire_527;
    wire new_Jinkela_wire_8232;
    wire new_Jinkela_wire_10118;
    wire new_Jinkela_wire_4450;
    wire new_Jinkela_wire_4220;
    wire new_Jinkela_wire_9662;
    wire new_Jinkela_wire_5570;
    wire new_Jinkela_wire_7822;
    wire new_Jinkela_wire_7931;
    wire new_Jinkela_wire_8299;
    wire new_Jinkela_wire_10309;
    wire new_Jinkela_wire_977;
    wire new_Jinkela_wire_2750;
    wire new_Jinkela_wire_3100;
    wire new_Jinkela_wire_10027;
    wire new_Jinkela_wire_9531;
    wire n_1090_;
    wire new_Jinkela_wire_8598;
    wire new_net_2562;
    wire new_Jinkela_wire_1532;
    wire new_Jinkela_wire_7902;
    wire new_Jinkela_wire_6848;
    wire new_Jinkela_wire_5118;
    wire new_Jinkela_wire_4692;
    wire new_Jinkela_wire_5503;
    wire new_Jinkela_wire_1379;
    wire new_Jinkela_wire_9434;
    wire new_Jinkela_wire_3555;
    wire new_Jinkela_wire_2409;
    wire new_Jinkela_wire_4505;
    wire n_0577_;
    wire new_Jinkela_wire_4983;
    wire new_Jinkela_wire_717;
    wire new_Jinkela_wire_10044;
    wire n_1053_;
    wire new_Jinkela_wire_7510;
    wire new_Jinkela_wire_1229;
    wire new_Jinkela_wire_5457;
    wire new_Jinkela_wire_2495;
    wire new_Jinkela_wire_163;
    wire new_Jinkela_wire_9820;
    wire new_Jinkela_wire_5219;
    wire new_Jinkela_wire_1181;
    wire new_Jinkela_wire_4546;
    wire new_Jinkela_wire_9305;
    wire new_Jinkela_wire_7155;
    wire new_Jinkela_wire_9043;
    wire new_Jinkela_wire_9016;
    wire new_Jinkela_wire_2707;
    wire new_Jinkela_wire_1265;
    wire new_Jinkela_wire_2278;
    wire new_Jinkela_wire_7514;
    wire n_0311_;
    wire new_Jinkela_wire_8168;
    wire new_Jinkela_wire_128;
    wire n_0930_;
    wire n_0841_;
    wire new_Jinkela_wire_8327;
    wire new_Jinkela_wire_4252;
    wire new_Jinkela_wire_10228;
    wire new_Jinkela_wire_3884;
    wire new_Jinkela_wire_7635;
    wire n_0344_;
    wire new_Jinkela_wire_9749;
    wire new_Jinkela_wire_9229;
    wire new_Jinkela_wire_188;
    wire new_Jinkela_wire_213;
    wire new_Jinkela_wire_6590;
    wire n_1321_;
    wire new_Jinkela_wire_6648;
    wire new_Jinkela_wire_593;
    wire new_Jinkela_wire_9556;
    wire new_Jinkela_wire_7935;
    wire new_Jinkela_wire_1110;
    wire n_1326_;
    wire new_Jinkela_wire_105;
    wire new_Jinkela_wire_3677;
    wire new_Jinkela_wire_5642;
    wire new_Jinkela_wire_7318;
    wire new_Jinkela_wire_10223;
    wire new_Jinkela_wire_3702;
    wire new_Jinkela_wire_2393;
    wire new_Jinkela_wire_3665;
    wire new_Jinkela_wire_5732;
    wire new_Jinkela_wire_7210;
    wire new_Jinkela_wire_792;
    wire new_Jinkela_wire_9387;
    wire new_Jinkela_wire_5111;
    wire new_Jinkela_wire_6156;
    wire n_0300_;
    wire new_Jinkela_wire_3330;
    wire new_Jinkela_wire_4072;
    wire new_Jinkela_wire_7056;
    wire new_Jinkela_wire_10103;
    wire n_1300_;
    wire new_Jinkela_wire_249;
    wire new_Jinkela_wire_8589;
    wire new_Jinkela_wire_10060;
    wire new_Jinkela_wire_9102;
    wire new_Jinkela_wire_766;
    wire new_Jinkela_wire_3605;
    wire new_Jinkela_wire_8271;
    wire new_Jinkela_wire_5129;
    wire new_Jinkela_wire_8560;
    wire new_Jinkela_wire_1674;
    wire new_Jinkela_wire_3800;
    wire new_Jinkela_wire_6352;
    wire new_Jinkela_wire_8565;
    wire new_Jinkela_wire_1316;
    wire new_Jinkela_wire_3760;
    wire new_Jinkela_wire_7516;
    wire new_Jinkela_wire_986;
    wire new_Jinkela_wire_10510;
    wire new_Jinkela_wire_2245;
    wire new_Jinkela_wire_1654;
    wire new_Jinkela_wire_1480;
    wire new_Jinkela_wire_7322;
    wire new_Jinkela_wire_5973;
    wire new_Jinkela_wire_911;
    wire new_Jinkela_wire_7779;
    wire new_Jinkela_wire_8129;
    wire new_Jinkela_wire_3383;
    wire new_Jinkela_wire_9439;
    wire new_Jinkela_wire_9190;
    wire new_Jinkela_wire_1331;
    wire new_Jinkela_wire_2181;
    wire new_Jinkela_wire_1946;
    wire new_Jinkela_wire_251;
    wire new_Jinkela_wire_10357;
    wire new_Jinkela_wire_7938;
    wire new_Jinkela_wire_6399;
    wire new_Jinkela_wire_8542;
    wire n_1034_;
    wire new_Jinkela_wire_111;
    wire new_Jinkela_wire_9076;
    wire new_Jinkela_wire_7803;
    wire new_Jinkela_wire_5188;
    wire new_Jinkela_wire_2202;
    wire new_Jinkela_wire_4306;
    wire new_Jinkela_wire_5115;
    wire new_Jinkela_wire_2861;
    wire new_Jinkela_wire_10160;
    wire new_Jinkela_wire_2644;
    wire new_Jinkela_wire_8235;
    wire new_Jinkela_wire_3719;
    wire new_Jinkela_wire_7526;
    wire new_Jinkela_wire_1896;
    wire n_0054_;
    wire new_Jinkela_wire_4506;
    wire new_Jinkela_wire_7649;
    wire new_Jinkela_wire_1519;
    wire new_Jinkela_wire_6695;
    wire new_Jinkela_wire_2163;
    wire new_Jinkela_wire_5065;
    wire new_Jinkela_wire_4241;
    wire new_Jinkela_wire_7477;
    wire new_Jinkela_wire_3278;
    wire new_Jinkela_wire_4013;
    wire n_1006_;
    wire new_Jinkela_wire_4761;
    wire new_Jinkela_wire_3185;
    wire new_Jinkela_wire_2544;
    wire new_Jinkela_wire_1491;
    wire new_Jinkela_wire_386;
    wire n_0821_;
    wire new_Jinkela_wire_3835;
    wire new_Jinkela_wire_4155;
    wire new_Jinkela_wire_886;
    wire n_0936_;
    wire n_0332_;
    wire new_Jinkela_wire_8049;
    wire new_Jinkela_wire_9864;
    wire new_Jinkela_wire_481;
    wire new_Jinkela_wire_7768;
    wire new_Jinkela_wire_2730;
    wire new_Jinkela_wire_2293;
    wire new_Jinkela_wire_9507;
    wire new_Jinkela_wire_9374;
    wire new_Jinkela_wire_1717;
    wire new_Jinkela_wire_7404;
    wire new_Jinkela_wire_9475;
    wire new_Jinkela_wire_2470;
    wire new_Jinkela_wire_987;
    wire n_0004_;
    wire new_Jinkela_wire_3507;
    wire new_Jinkela_wire_1657;
    wire new_Jinkela_wire_5436;
    wire new_Jinkela_wire_8536;
    wire new_Jinkela_wire_5435;
    wire new_Jinkela_wire_583;
    wire n_0896_;
    wire new_Jinkela_wire_10176;
    wire new_Jinkela_wire_2207;
    wire new_Jinkela_wire_3589;
    wire new_Jinkela_wire_1861;
    wire new_Jinkela_wire_8106;
    wire new_Jinkela_wire_2879;
    wire n_0191_;
    wire n_1102_;
    wire new_Jinkela_wire_1076;
    wire new_Jinkela_wire_9035;
    wire new_Jinkela_wire_7905;
    wire new_Jinkela_wire_1144;
    wire new_Jinkela_wire_2525;
    wire new_Jinkela_wire_5170;
    wire new_Jinkela_wire_3968;
    wire new_Jinkela_wire_302;
    wire new_Jinkela_wire_4070;
    wire new_Jinkela_wire_10618;
    wire new_Jinkela_wire_9094;
    wire new_Jinkela_wire_8764;
    wire new_Jinkela_wire_1193;
    wire new_Jinkela_wire_9388;
    wire new_Jinkela_wire_1143;
    wire new_Jinkela_wire_1603;
    wire new_Jinkela_wire_5953;
    wire new_Jinkela_wire_5400;
    wire new_Jinkela_wire_8195;
    wire new_Jinkela_wire_5333;
    wire new_Jinkela_wire_5472;
    wire new_Jinkela_wire_870;
    wire new_Jinkela_wire_2044;
    wire new_Jinkela_wire_8610;
    wire new_Jinkela_wire_337;
    wire new_Jinkela_wire_9909;
    wire new_Jinkela_wire_5437;
    wire new_Jinkela_wire_4267;
    wire new_Jinkela_wire_8916;
    wire new_Jinkela_wire_2822;
    wire n_0546_;
    wire new_Jinkela_wire_5041;
    wire new_Jinkela_wire_7913;
    wire new_Jinkela_wire_6556;
    wire new_Jinkela_wire_8070;
    wire new_Jinkela_wire_3676;
    wire new_Jinkela_wire_5971;
    wire new_net_2545;
    wire new_Jinkela_wire_6774;
    wire new_Jinkela_wire_2640;
    wire new_Jinkela_wire_1187;
    wire new_Jinkela_wire_10184;
    wire new_Jinkela_wire_6464;
    wire new_Jinkela_wire_9478;
    wire new_Jinkela_wire_6099;
    wire new_Jinkela_wire_7835;
    wire new_Jinkela_wire_3669;
    wire new_Jinkela_wire_8091;
    wire new_Jinkela_wire_4599;
    wire new_Jinkela_wire_1897;
    wire new_Jinkela_wire_7671;
    wire new_Jinkela_wire_2946;
    wire new_Jinkela_wire_3038;
    wire new_Jinkela_wire_5654;
    wire new_Jinkela_wire_6992;
    wire new_Jinkela_wire_9593;
    wire new_Jinkela_wire_178;
    wire new_Jinkela_wire_4300;
    wire new_Jinkela_wire_9901;
    wire new_Jinkela_wire_6970;
    wire new_Jinkela_wire_9936;
    wire new_Jinkela_wire_4197;
    wire new_Jinkela_wire_6127;
    wire new_Jinkela_wire_70;
    wire new_Jinkela_wire_10512;
    wire new_Jinkela_wire_8711;
    wire n_0211_;
    wire new_Jinkela_wire_6218;
    wire new_Jinkela_wire_945;
    wire new_Jinkela_wire_3808;
    wire new_Jinkela_wire_8097;
    wire new_Jinkela_wire_9069;
    wire new_Jinkela_wire_10219;
    wire new_Jinkela_wire_4000;
    wire new_Jinkela_wire_3460;
    wire new_Jinkela_wire_10541;
    wire new_Jinkela_wire_1464;
    wire new_Jinkela_wire_882;
    wire new_Jinkela_wire_4248;
    wire new_Jinkela_wire_4066;
    wire new_Jinkela_wire_6091;
    wire new_Jinkela_wire_10203;
    wire new_Jinkela_wire_4315;
    wire new_Jinkela_wire_969;
    wire new_Jinkela_wire_9146;
    wire new_Jinkela_wire_10312;
    wire new_Jinkela_wire_4044;
    wire new_Jinkela_wire_10180;
    wire new_Jinkela_wire_7339;
    wire n_0377_;
    wire new_Jinkela_wire_9049;
    wire new_Jinkela_wire_9154;
    wire new_Jinkela_wire_3557;
    wire n_1109_;
    wire new_Jinkela_wire_3796;
    wire new_Jinkela_wire_4177;
    wire new_Jinkela_wire_12;
    wire new_Jinkela_wire_4998;
    wire new_Jinkela_wire_4359;
    wire new_Jinkela_wire_7970;
    wire new_Jinkela_wire_6896;
    wire new_Jinkela_wire_6202;
    wire new_Jinkela_wire_5794;
    wire new_Jinkela_wire_5560;
    wire new_Jinkela_wire_9;
    wire new_Jinkela_wire_5038;
    wire new_Jinkela_wire_3225;
    wire new_Jinkela_wire_696;
    wire new_Jinkela_wire_7581;
    wire new_Jinkela_wire_7838;
    wire new_Jinkela_wire_6546;
    wire new_Jinkela_wire_8151;
    wire new_Jinkela_wire_7650;
    wire new_Jinkela_wire_1199;
    wire new_Jinkela_wire_2306;
    wire new_Jinkela_wire_8073;
    wire new_Jinkela_wire_10296;
    wire new_Jinkela_wire_8668;
    wire new_Jinkela_wire_7975;
    wire new_Jinkela_wire_5587;
    wire new_Jinkela_wire_6136;
    wire new_Jinkela_wire_3958;
    wire n_0371_;
    wire new_Jinkela_wire_9776;
    wire new_Jinkela_wire_7511;
    wire new_Jinkela_wire_3208;
    wire new_Jinkela_wire_2522;
    wire new_Jinkela_wire_4550;
    wire new_Jinkela_wire_5877;
    wire new_Jinkela_wire_2074;
    wire new_Jinkela_wire_3140;
    wire new_Jinkela_wire_6396;
    wire new_Jinkela_wire_851;
    wire new_Jinkela_wire_4528;
    wire new_Jinkela_wire_3003;
    wire new_Jinkela_wire_4905;
    wire new_Jinkela_wire_6488;
    wire new_Jinkela_wire_2600;
    wire new_Jinkela_wire_3005;
    wire new_Jinkela_wire_2201;
    wire new_Jinkela_wire_3966;
    wire n_0911_;
    wire new_Jinkela_wire_2885;
    wire n_0689_;
    wire new_Jinkela_wire_2669;
    wire new_Jinkela_wire_8274;
    wire new_Jinkela_wire_8099;
    wire new_Jinkela_wire_8324;
    wire new_Jinkela_wire_10481;
    wire new_Jinkela_wire_6024;
    wire new_Jinkela_wire_7230;
    wire new_Jinkela_wire_3539;
    wire new_Jinkela_wire_8079;
    wire new_Jinkela_wire_7912;
    wire n_0402_;
    wire n_1255_;
    wire new_Jinkela_wire_6550;
    wire new_Jinkela_wire_2305;
    wire new_Jinkela_wire_10392;
    wire new_Jinkela_wire_165;
    wire new_Jinkela_wire_4215;
    wire new_Jinkela_wire_1373;
    wire new_Jinkela_wire_1682;
    wire new_Jinkela_wire_7152;
    wire new_Jinkela_wire_4161;
    wire new_Jinkela_wire_3032;
    wire new_Jinkela_wire_4253;
    wire new_Jinkela_wire_3810;
    wire n_0803_;
    wire new_Jinkela_wire_5668;
    wire new_Jinkela_wire_8222;
    wire new_Jinkela_wire_6829;
    wire new_Jinkela_wire_496;
    wire new_Jinkela_wire_3890;
    wire new_Jinkela_wire_3623;
    wire new_Jinkela_wire_8722;
    wire new_Jinkela_wire_4034;
    wire n_1082_;
    wire new_Jinkela_wire_7568;
    wire new_Jinkela_wire_9863;
    wire new_Jinkela_wire_3312;
    wire new_Jinkela_wire_4795;
    wire new_Jinkela_wire_1769;
    wire new_Jinkela_wire_7324;
    wire new_Jinkela_wire_2212;
    wire new_Jinkela_wire_10388;
    wire new_Jinkela_wire_10625;
    wire new_Jinkela_wire_838;
    wire new_Jinkela_wire_9582;
    wire new_Jinkela_wire_6119;
    wire new_Jinkela_wire_4361;
    wire new_Jinkela_wire_891;
    wire new_Jinkela_wire_3371;
    wire n_1178_;
    wire n_0415_;
    wire n_0201_;
    wire new_Jinkela_wire_6473;
    wire n_1081_;
    wire n_1173_;
    wire new_Jinkela_wire_9647;
    wire new_Jinkela_wire_4481;
    wire new_Jinkela_wire_9411;
    wire new_Jinkela_wire_96;
    wire new_Jinkela_wire_7169;
    wire n_0238_;
    wire n_0033_;
    wire new_Jinkela_wire_7496;
    wire n_0403_;
    wire new_Jinkela_wire_5024;
    wire new_Jinkela_wire_9459;
    wire new_Jinkela_wire_3239;
    wire new_Jinkela_wire_2140;
    wire new_Jinkela_wire_10374;
    wire new_Jinkela_wire_3580;
    wire new_Jinkela_wire_5722;
    wire new_Jinkela_wire_4569;
    wire new_Jinkela_wire_4748;
    wire new_Jinkela_wire_6969;
    wire new_Jinkela_wire_3023;
    wire new_Jinkela_wire_9881;
    wire new_Jinkela_wire_1712;
    wire new_Jinkela_wire_6806;
    wire new_Jinkela_wire_102;
    wire new_Jinkela_wire_3286;
    wire new_Jinkela_wire_4322;
    wire new_Jinkela_wire_3910;
    wire new_Jinkela_wire_5935;
    wire new_Jinkela_wire_9836;
    wire new_Jinkela_wire_4287;
    wire new_Jinkela_wire_7237;
    wire new_Jinkela_wire_7831;
    wire new_Jinkela_wire_4937;
    wire new_Jinkela_wire_2732;
    wire new_Jinkela_wire_7515;
    wire new_Jinkela_wire_5999;
    wire new_Jinkela_wire_4334;
    wire new_Jinkela_wire_9915;
    wire new_Jinkela_wire_1632;
    wire new_Jinkela_wire_4288;
    wire new_Jinkela_wire_5905;
    wire new_Jinkela_wire_5196;
    wire new_Jinkela_wire_7453;
    wire new_Jinkela_wire_9553;
    wire new_Jinkela_wire_3636;
    wire new_Jinkela_wire_2748;
    wire new_Jinkela_wire_9645;
    wire n_0389_;
    wire new_Jinkela_wire_2012;
    wire new_Jinkela_wire_1796;
    wire new_Jinkela_wire_1738;
    wire new_Jinkela_wire_3748;
    wire new_Jinkela_wire_7483;
    wire new_Jinkela_wire_4810;
    wire new_Jinkela_wire_2482;
    wire new_Jinkela_wire_1056;
    wire new_Jinkela_wire_6943;
    wire new_Jinkela_wire_6363;
    wire new_Jinkela_wire_5961;
    wire new_Jinkela_wire_4707;
    wire new_Jinkela_wire_8410;
    wire n_1103_;
    wire new_Jinkela_wire_8516;
    wire new_Jinkela_wire_4320;
    wire new_Jinkela_wire_6035;
    wire new_Jinkela_wire_9306;
    wire new_Jinkela_wire_9390;
    wire new_Jinkela_wire_8958;
    wire new_Jinkela_wire_9218;
    wire new_Jinkela_wire_8524;
    wire n_0088_;
    wire new_Jinkela_wire_6074;
    wire new_Jinkela_wire_7594;
    wire new_Jinkela_wire_9686;
    wire new_Jinkela_wire_8489;
    wire n_0806_;
    wire new_Jinkela_wire_2499;
    wire new_Jinkela_wire_8346;
    wire new_Jinkela_wire_3109;
    wire new_Jinkela_wire_9649;
    wire new_Jinkela_wire_8453;
    wire new_Jinkela_wire_3903;
    wire new_Jinkela_wire_701;
    wire new_Jinkela_wire_3542;
    wire new_Jinkela_wire_8849;
    wire new_Jinkela_wire_18;
    wire new_Jinkela_wire_7708;
    wire new_Jinkela_wire_9840;
    wire new_Jinkela_wire_9500;
    wire new_Jinkela_wire_658;
    wire new_Jinkela_wire_2860;
    wire new_Jinkela_wire_3008;
    wire new_Jinkela_wire_9288;
    wire new_Jinkela_wire_6280;
    wire new_Jinkela_wire_4193;
    wire new_Jinkela_wire_1829;
    wire new_Jinkela_wire_8229;
    wire n_1124_;
    wire new_Jinkela_wire_4164;
    wire new_Jinkela_wire_3869;
    wire new_Jinkela_wire_5209;
    wire new_Jinkela_wire_1987;
    wire new_Jinkela_wire_2777;
    wire new_Jinkela_wire_5801;
    wire new_Jinkela_wire_2186;
    wire new_Jinkela_wire_3633;
    wire new_Jinkela_wire_5889;
    wire new_Jinkela_wire_5981;
    wire new_Jinkela_wire_3868;
    wire new_Jinkela_wire_9667;
    wire new_Jinkela_wire_5045;
    wire n_1339_;
    wire n_0701_;
    wire new_Jinkela_wire_4172;
    wire new_Jinkela_wire_10068;
    wire new_Jinkela_wire_3218;
    wire new_Jinkela_wire_9325;
    wire new_Jinkela_wire_5480;
    wire new_Jinkela_wire_11;
    wire new_Jinkela_wire_387;
    wire new_Jinkela_wire_8824;
    wire new_Jinkela_wire_6891;
    wire new_Jinkela_wire_8539;
    wire new_Jinkela_wire_2407;
    wire new_Jinkela_wire_3050;
    wire new_Jinkela_wire_6034;
    wire n_0790_;
    wire new_Jinkela_wire_4377;
    wire new_Jinkela_wire_5873;
    wire new_Jinkela_wire_6084;
    wire new_Jinkela_wire_2662;
    wire new_Jinkela_wire_1053;
    wire new_Jinkela_wire_2746;
    wire new_Jinkela_wire_3987;
    wire new_Jinkela_wire_117;
    wire new_Jinkela_wire_8901;
    wire new_Jinkela_wire_5361;
    wire new_Jinkela_wire_4246;
    wire new_Jinkela_wire_1707;
    wire new_Jinkela_wire_722;
    wire new_Jinkela_wire_9659;
    wire new_Jinkela_wire_3089;
    wire new_Jinkela_wire_5004;
    wire new_Jinkela_wire_1197;
    wire new_Jinkela_wire_4798;
    wire new_Jinkela_wire_4098;
    wire new_Jinkela_wire_529;
    wire new_Jinkela_wire_2498;
    wire new_Jinkela_wire_2601;
    wire new_Jinkela_wire_3661;
    wire new_Jinkela_wire_1687;
    wire new_Jinkela_wire_6439;
    wire new_Jinkela_wire_5325;
    wire new_Jinkela_wire_2412;
    wire new_Jinkela_wire_2106;
    wire new_Jinkela_wire_7104;
    wire new_Jinkela_wire_4134;
    wire new_Jinkela_wire_9223;
    wire new_Jinkela_wire_9286;
    wire n_1226_;
    wire new_Jinkela_wire_9106;
    wire new_Jinkela_wire_7276;
    wire new_Jinkela_wire_9177;
    wire new_Jinkela_wire_9160;
    wire new_Jinkela_wire_5002;
    wire new_Jinkela_wire_298;
    wire new_Jinkela_wire_6331;
    wire new_Jinkela_wire_5258;
    wire new_Jinkela_wire_4224;
    wire new_Jinkela_wire_7906;
    wire new_Jinkela_wire_724;
    wire new_Jinkela_wire_2570;
    wire n_1212_;
    wire new_Jinkela_wire_4783;
    wire new_Jinkela_wire_9797;
    wire n_0979_;
    wire new_Jinkela_wire_9179;
    wire new_Jinkela_wire_3431;
    wire new_Jinkela_wire_642;
    wire new_Jinkela_wire_4872;
    wire new_Jinkela_wire_4612;
    wire new_Jinkela_wire_9406;
    wire new_Jinkela_wire_2083;
    wire new_Jinkela_wire_9481;
    wire new_Jinkela_wire_5863;
    wire new_Jinkela_wire_2045;
    wire new_Jinkela_wire_9416;
    wire new_Jinkela_wire_4060;
    wire new_Jinkela_wire_5179;
    wire new_Jinkela_wire_2343;
    wire n_0018_;
    wire new_Jinkela_wire_4358;
    wire n_0052_;
    wire new_Jinkela_wire_4873;
    wire new_Jinkela_wire_9427;
    wire new_Jinkela_wire_8060;
    wire new_Jinkela_wire_5506;
    wire new_Jinkela_wire_8381;
    wire new_Jinkela_wire_7984;
    wire new_Jinkela_wire_7934;
    wire new_Jinkela_wire_57;
    wire new_Jinkela_wire_10410;
    wire new_Jinkela_wire_404;
    wire new_Jinkela_wire_2414;
    wire n_0733_;
    wire new_Jinkela_wire_3613;
    wire new_Jinkela_wire_2553;
    wire n_1060_;
    wire new_Jinkela_wire_7059;
    wire new_Jinkela_wire_1757;
    wire new_Jinkela_wire_9346;
    wire new_Jinkela_wire_349;
    wire new_Jinkela_wire_8181;
    wire n_0568_;
    wire new_Jinkela_wire_4616;
    wire new_Jinkela_wire_3558;
    wire n_1251_;
    wire new_Jinkela_wire_5839;
    wire new_Jinkela_wire_64;
    wire new_Jinkela_wire_1521;
    wire new_Jinkela_wire_10268;
    wire new_Jinkela_wire_30;
    wire new_Jinkela_wire_9871;
    wire new_Jinkela_wire_4938;
    wire new_Jinkela_wire_1786;
    wire new_Jinkela_wire_7603;
    wire n_0696_;
    wire new_Jinkela_wire_4026;
    wire new_Jinkela_wire_8640;
    wire new_Jinkela_wire_1754;
    wire new_Jinkela_wire_8395;
    wire new_Jinkela_wire_9521;
    wire n_1049_;
    wire new_Jinkela_wire_3067;
    wire n_0797_;
    wire new_Jinkela_wire_9151;
    wire new_Jinkela_wire_9355;
    wire new_Jinkela_wire_3338;
    wire new_Jinkela_wire_8822;
    wire new_Jinkela_wire_4115;
    wire new_Jinkela_wire_10007;
    wire new_Jinkela_wire_7402;
    wire new_Jinkela_wire_4511;
    wire n_0565_;
    wire new_Jinkela_wire_1348;
    wire n_0189_;
    wire new_Jinkela_wire_19;
    wire new_Jinkela_wire_8061;
    wire new_Jinkela_wire_6543;
    wire n_0770_;
    wire n_0892_;
    wire n_0257_;
    wire new_Jinkela_wire_6126;
    wire new_Jinkela_wire_2962;
    wire n_0261_;
    wire new_Jinkela_wire_7338;
    wire new_Jinkela_wire_483;
    wire new_Jinkela_wire_394;
    wire new_Jinkela_wire_1752;
    wire new_Jinkela_wire_7579;
    wire new_Jinkela_wire_4503;
    wire new_Jinkela_wire_1015;
    wire new_Jinkela_wire_9814;
    wire new_Jinkela_wire_873;
    wire n_0682_;
    wire new_Jinkela_wire_4336;
    wire new_Jinkela_wire_10517;
    wire new_Jinkela_wire_2167;
    wire new_Jinkela_wire_173;
    wire new_Jinkela_wire_5028;
    wire new_Jinkela_wire_1981;
    wire new_Jinkela_wire_7563;
    wire new_Jinkela_wire_1785;
    wire new_Jinkela_wire_8616;
    wire new_Jinkela_wire_8712;
    wire new_Jinkela_wire_5653;
    wire new_Jinkela_wire_6142;
    wire new_Jinkela_wire_3055;
    wire new_Jinkela_wire_2865;
    wire new_Jinkela_wire_7071;
    wire new_Jinkela_wire_3250;
    wire new_Jinkela_wire_3162;
    wire n_1342_;
    wire n_1104_;
    wire n_1183_;
    wire new_Jinkela_wire_9858;
    wire new_Jinkela_wire_5202;
    wire new_Jinkela_wire_10032;
    wire new_Jinkela_wire_3603;
    wire new_Jinkela_wire_4604;
    wire new_Jinkela_wire_2379;
    wire new_Jinkela_wire_6565;
    wire new_Jinkela_wire_1011;
    wire new_Jinkela_wire_2779;
    wire new_Jinkela_wire_2968;
    wire new_Jinkela_wire_1873;
    wire new_Jinkela_wire_3415;
    wire new_Jinkela_wire_6147;
    wire new_Jinkela_wire_3895;
    wire new_Jinkela_wire_3472;
    wire new_Jinkela_wire_1225;
    wire new_Jinkela_wire_3687;
    wire new_Jinkela_wire_7093;
    wire new_Jinkela_wire_6110;
    wire new_Jinkela_wire_3896;
    wire new_Jinkela_wire_1323;
    wire new_Jinkela_wire_112;
    wire new_Jinkela_wire_6536;
    wire new_Jinkela_wire_4471;
    wire new_Jinkela_wire_7103;
    wire new_Jinkela_wire_511;
    wire new_Jinkela_wire_7258;
    wire new_Jinkela_wire_7574;
    wire new_Jinkela_wire_3336;
    wire n_0397_;
    wire new_Jinkela_wire_7233;
    wire new_Jinkela_wire_9377;
    wire new_Jinkela_wire_9898;
    wire new_Jinkela_wire_8048;
    wire new_Jinkela_wire_2033;
    wire new_Jinkela_wire_4277;
    wire new_Jinkela_wire_10584;
    wire new_Jinkela_wire_5256;
    wire new_Jinkela_wire_8888;
    wire new_Jinkela_wire_8020;
    wire new_Jinkela_wire_3325;
    wire new_Jinkela_wire_6349;
    wire new_Jinkela_wire_1402;
    wire new_Jinkela_wire_5620;
    wire new_Jinkela_wire_7366;
    wire new_Jinkela_wire_9234;
    wire new_Jinkela_wire_10244;
    wire new_Jinkela_wire_4768;
    wire new_Jinkela_wire_3198;
    wire new_Jinkela_wire_9126;
    wire new_Jinkela_wire_5157;
    wire new_Jinkela_wire_2035;
    wire new_Jinkela_wire_10187;
    wire n_0574_;
    wire new_Jinkela_wire_2040;
    wire new_Jinkela_wire_4456;
    wire new_Jinkela_wire_2890;
    wire new_Jinkela_wire_2195;
    wire new_Jinkela_wire_8403;
    wire new_Jinkela_wire_4709;
    wire new_Jinkela_wire_3935;
    wire n_0552_;
    wire new_Jinkela_wire_2492;
    wire n_0903_;
    wire new_Jinkela_wire_4328;
    wire new_Jinkela_wire_9246;
    wire new_Jinkela_wire_2144;
    wire new_Jinkela_wire_8780;
    wire new_Jinkela_wire_10033;
    wire new_Jinkela_wire_237;
    wire new_Jinkela_wire_7879;
    wire new_Jinkela_wire_10181;
    wire new_Jinkela_wire_3159;
    wire new_Jinkela_wire_3892;
    wire new_Jinkela_wire_1433;
    wire new_Jinkela_wire_8187;
    wire new_Jinkela_wire_8094;
    wire n_0439_;
    wire new_Jinkela_wire_821;
    wire new_Jinkela_wire_2471;
    wire new_Jinkela_wire_8032;
    wire new_Jinkela_wire_10303;
    wire new_Jinkela_wire_3267;
    wire n_0157_;
    wire new_Jinkela_wire_2183;
    wire n_0312_;
    wire n_0441_;
    wire new_Jinkela_wire_10100;
    wire new_Jinkela_wire_1058;
    wire n_0611_;
    wire new_Jinkela_wire_6748;
    wire new_Jinkela_wire_1618;
    wire new_Jinkela_wire_2232;
    wire new_Jinkela_wire_3900;
    wire new_Jinkela_wire_1442;
    wire new_Jinkela_wire_4533;
    wire n_0816_;
    wire new_Jinkela_wire_37;
    wire new_Jinkela_wire_4232;
    wire new_Jinkela_wire_8696;
    wire new_Jinkela_wire_10591;
    wire new_Jinkela_wire_9221;
    wire new_Jinkela_wire_6334;
    wire new_Jinkela_wire_8784;
    wire new_Jinkela_wire_4663;
    wire new_Jinkela_wire_6557;
    wire new_Jinkela_wire_7892;
    wire new_Jinkela_wire_9273;
    wire new_Jinkela_wire_7775;
    wire new_Jinkela_wire_6227;
    wire n_0093_;
    wire new_Jinkela_wire_2102;
    wire new_Jinkela_wire_7147;
    wire new_Jinkela_wire_9144;
    wire new_Jinkela_wire_2401;
    wire n_0681_;
    wire n_1256_;
    wire n_0222_;
    wire n_0608_;
    wire new_Jinkela_wire_9955;
    wire new_Jinkela_wire_7667;
    wire new_Jinkela_wire_6197;
    wire new_Jinkela_wire_7010;
    wire new_Jinkela_wire_5048;
    wire new_Jinkela_wire_1695;
    wire new_Jinkela_wire_9281;
    wire new_Jinkela_wire_4740;
    wire n_0042_;
    wire new_Jinkela_wire_6299;
    wire new_Jinkela_wire_4190;
    wire new_Jinkela_wire_7242;
    wire new_Jinkela_wire_1065;
    wire new_Jinkela_wire_7294;
    wire new_Jinkela_wire_2920;
    wire new_Jinkela_wire_7088;
    wire n_0520_;
    wire n_0092_;
    wire n_0062_;
    wire new_Jinkela_wire_3883;
    wire new_Jinkela_wire_6851;
    wire new_Jinkela_wire_2583;
    wire new_Jinkela_wire_940;
    wire new_Jinkela_wire_190;
    wire new_Jinkela_wire_5505;
    wire new_Jinkela_wire_2480;
    wire new_Jinkela_wire_1625;
    wire n_0679_;
    wire n_0746_;
    wire new_Jinkela_wire_4063;
    wire n_0657_;
    wire new_Jinkela_wire_3969;
    wire new_Jinkela_wire_5315;
    wire new_Jinkela_wire_1262;
    wire new_Jinkela_wire_8254;
    wire new_Jinkela_wire_6342;
    wire new_Jinkela_wire_7830;
    wire n_0065_;
    wire n_0085_;
    wire new_Jinkela_wire_10169;
    wire new_Jinkela_wire_2574;
    wire new_Jinkela_wire_9938;
    wire n_0836_;
    wire new_Jinkela_wire_6547;
    wire new_Jinkela_wire_3604;
    wire new_Jinkela_wire_103;
    wire n_0999_;
    wire n_0964_;
    wire new_Jinkela_wire_4593;
    wire new_Jinkela_wire_9829;
    wire new_Jinkela_wire_10064;
    wire new_Jinkela_wire_4845;
    wire n_1294_;
    wire new_Jinkela_wire_4199;
    wire new_Jinkela_wire_7;
    wire new_Jinkela_wire_9842;
    wire new_Jinkela_wire_10182;
    wire n_0223_;
    wire new_Jinkela_wire_1954;
    wire new_Jinkela_wire_4352;
    wire new_Jinkela_wire_10198;
    wire new_Jinkela_wire_2782;
    wire new_Jinkela_wire_5453;
    wire new_Jinkela_wire_4135;
    wire new_Jinkela_wire_3433;
    wire new_Jinkela_wire_964;
    wire n_0230_;
    wire new_Jinkela_wire_622;
    wire new_Jinkela_wire_1112;
    wire new_Jinkela_wire_2439;
    wire n_0457_;
    wire new_Jinkela_wire_1194;
    wire new_Jinkela_wire_6101;
    wire new_Jinkela_wire_5684;
    wire new_Jinkela_wire_2751;
    wire new_Jinkela_wire_9800;
    wire new_Jinkela_wire_6874;
    wire n_1236_;
    wire new_Jinkela_wire_4089;
    wire new_Jinkela_wire_5374;
    wire new_Jinkela_wire_557;
    wire new_Jinkela_wire_9143;
    wire new_Jinkela_wire_7766;
    wire new_Jinkela_wire_4654;
    wire new_Jinkela_wire_6060;
    wire new_Jinkela_wire_8839;
    wire n_0372_;
    wire new_Jinkela_wire_8240;
    wire new_Jinkela_wire_7571;
    wire new_Jinkela_wire_9260;
    wire new_Jinkela_wire_3999;
    wire new_Jinkela_wire_7107;
    wire new_Jinkela_wire_1788;
    wire new_Jinkela_wire_2847;
    wire new_Jinkela_wire_6572;
    wire new_Jinkela_wire_3887;
    wire new_Jinkela_wire_2760;
    wire new_Jinkela_wire_2091;
    wire new_Jinkela_wire_7908;
    wire new_Jinkela_wire_10241;
    wire new_Jinkela_wire_8697;
    wire new_Jinkela_wire_5499;
    wire n_0760_;
    wire new_Jinkela_wire_1716;
    wire new_Jinkela_wire_7026;
    wire new_Jinkela_wire_9527;
    wire new_Jinkela_wire_5144;
    wire new_Jinkela_wire_3281;
    wire new_Jinkela_wire_10310;
    wire new_Jinkela_wire_4163;
    wire new_Jinkela_wire_6433;
    wire n_0305_;
    wire new_Jinkela_wire_7493;
    wire new_Jinkela_wire_6701;
    wire new_Jinkela_wire_9861;
    wire n_0731_;
    wire new_Jinkela_wire_6846;
    wire new_Jinkela_wire_5796;
    wire new_Jinkela_wire_3786;
    wire new_Jinkela_wire_5536;
    wire new_Jinkela_wire_5539;
    wire new_Jinkela_wire_1624;
    wire new_Jinkela_wire_1100;
    wire new_Jinkela_wire_1090;
    wire new_Jinkela_wire_6621;
    wire n_0155_;
    wire new_Jinkela_wire_3916;
    wire new_Jinkela_wire_3404;
    wire new_Jinkela_wire_10119;
    wire new_Jinkela_wire_6822;
    wire new_Jinkela_wire_4691;
    wire new_Jinkela_wire_5602;
    wire n_0114_;
    wire new_Jinkela_wire_9609;
    wire new_Jinkela_wire_3543;
    wire new_net_10;
    wire new_Jinkela_wire_7498;
    wire new_Jinkela_wire_1329;
    wire n_0853_;
    wire new_Jinkela_wire_7701;
    wire new_Jinkela_wire_2594;
    wire new_Jinkela_wire_1633;
    wire new_Jinkela_wire_1037;
    wire n_1299_;
    wire new_Jinkela_wire_7821;
    wire new_Jinkela_wire_780;
    wire new_Jinkela_wire_3858;
    wire new_Jinkela_wire_8867;
    wire new_Jinkela_wire_7869;
    wire new_Jinkela_wire_10457;
    wire n_0179_;
    wire new_Jinkela_wire_3647;
    wire new_Jinkela_wire_8638;
    wire new_Jinkela_wire_8607;
    wire n_0890_;
    wire new_Jinkela_wire_1660;
    wire new_Jinkela_wire_4362;
    wire new_Jinkela_wire_7545;
    wire new_Jinkela_wire_9954;
    wire new_Jinkela_wire_4793;
    wire new_Jinkela_wire_9711;
    wire new_Jinkela_wire_2398;
    wire new_Jinkela_wire_3855;
    wire n_0086_;
    wire new_Jinkela_wire_2050;
    wire new_Jinkela_wire_6790;
    wire n_0234_;
    wire new_Jinkela_wire_385;
    wire n_0217_;
    wire new_Jinkela_wire_8707;
    wire new_Jinkela_wire_1743;
    wire new_Jinkela_wire_1423;
    wire new_Jinkela_wire_7140;
    wire new_Jinkela_wire_8727;
    wire new_Jinkela_wire_7629;
    wire n_0146_;
    wire new_Jinkela_wire_6367;
    wire new_Jinkela_wire_1237;
    wire new_Jinkela_wire_1368;
    wire new_Jinkela_wire_1587;
    wire new_Jinkela_wire_10423;
    wire new_Jinkela_wire_2378;
    wire new_Jinkela_wire_10021;
    wire new_Jinkela_wire_7360;
    wire new_Jinkela_wire_8535;
    wire new_Jinkela_wire_8180;
    wire new_Jinkela_wire_6070;
    wire new_Jinkela_wire_2626;
    wire new_Jinkela_wire_8515;
    wire n_0477_;
    wire new_Jinkela_wire_2591;
    wire new_Jinkela_wire_637;
    wire n_0729_;
    wire new_Jinkela_wire_3535;
    wire new_Jinkela_wire_7017;
    wire n_1318_;
    wire new_Jinkela_wire_1959;
    wire new_Jinkela_wire_9202;
    wire new_Jinkela_wire_1806;
    wire new_Jinkela_wire_4116;
    wire new_Jinkela_wire_4106;
    wire new_Jinkela_wire_10555;
    wire new_Jinkela_wire_9183;
    wire new_Jinkela_wire_79;
    wire new_Jinkela_wire_5439;
    wire new_Jinkela_wire_7199;
    wire new_Jinkela_wire_7438;
    wire n_0512_;
    wire new_Jinkela_wire_1935;
    wire new_Jinkela_wire_7997;
    wire new_Jinkela_wire_5148;
    wire new_Jinkela_wire_6746;
    wire new_Jinkela_wire_8406;
    wire new_Jinkela_wire_6914;
    wire new_Jinkela_wire_1780;
    wire new_Jinkela_wire_3096;
    wire new_Jinkela_wire_8606;
    wire new_Jinkela_wire_3571;
    wire new_Jinkela_wire_4137;
    wire new_Jinkela_wire_5917;
    wire new_Jinkela_wire_4465;
    wire new_Jinkela_wire_1489;
    wire new_Jinkela_wire_804;
    wire new_Jinkela_wire_4997;
    wire new_Jinkela_wire_2639;
    wire new_Jinkela_wire_8725;
    wire new_Jinkela_wire_8155;
    wire new_Jinkela_wire_3801;
    wire new_Jinkela_wire_6647;
    wire new_Jinkela_wire_2824;
    wire new_Jinkela_wire_5127;
    wire n_1332_;
    wire new_Jinkela_wire_3820;
    wire new_Jinkela_wire_9690;
    wire new_Jinkela_wire_2196;
    wire new_Jinkela_wire_6602;
    wire new_Jinkela_wire_6146;
    wire new_Jinkela_wire_10487;
    wire new_Jinkela_wire_54;
    wire new_Jinkela_wire_563;
    wire new_Jinkela_wire_3943;
    wire new_Jinkela_wire_3285;
    wire new_Jinkela_wire_7314;
    wire new_Jinkela_wire_4925;
    wire new_Jinkela_wire_4426;
    wire new_Jinkela_wire_2037;
    wire new_Jinkela_wire_4111;
    wire new_Jinkela_wire_2922;
    wire new_Jinkela_wire_6864;
    wire new_Jinkela_wire_2870;
    wire new_Jinkela_wire_9041;
    wire new_Jinkela_wire_914;
    wire new_Jinkela_wire_1938;
    wire new_Jinkela_wire_9900;
    wire n_0514_;
    wire new_Jinkela_wire_4496;
    wire new_Jinkela_wire_6684;
    wire new_Jinkela_wire_6002;
    wire new_Jinkela_wire_9490;
    wire new_Jinkela_wire_7407;
    wire n_0459_;
    wire new_Jinkela_wire_6678;
    wire new_Jinkela_wire_3120;
    wire n_0437_;
    wire new_Jinkela_wire_4059;
    wire new_Jinkela_wire_953;
    wire new_Jinkela_wire_2318;
    wire new_Jinkela_wire_9082;
    wire new_Jinkela_wire_798;
    wire new_Jinkela_wire_9774;
    wire new_Jinkela_wire_8508;
    wire new_Jinkela_wire_10578;
    wire new_Jinkela_wire_8881;
    wire new_Jinkela_wire_4144;
    wire new_Jinkela_wire_9872;
    wire new_Jinkela_wire_6628;
    wire n_0588_;
    wire new_Jinkela_wire_10598;
    wire n_1134_;
    wire n_1089_;
    wire new_Jinkela_wire_4229;
    wire new_Jinkela_wire_8735;
    wire new_Jinkela_wire_921;
    wire new_Jinkela_wire_3840;
    wire new_Jinkela_wire_3176;
    wire new_Jinkela_wire_2871;
    wire new_Jinkela_wire_2313;
    wire new_Jinkela_wire_7557;
    wire new_Jinkela_wire_1590;
    wire n_0920_;
    wire new_Jinkela_wire_9215;
    wire new_Jinkela_wire_1490;
    wire new_Jinkela_wire_1773;
    wire new_Jinkela_wire_5573;
    wire new_Jinkela_wire_10189;
    wire new_Jinkela_wire_7178;
    wire new_Jinkela_wire_9561;
    wire new_Jinkela_wire_4366;
    wire new_Jinkela_wire_1951;
    wire n_0691_;
    wire new_Jinkela_wire_7888;
    wire new_Jinkela_wire_8860;
    wire n_0676_;
    wire new_Jinkela_wire_271;
    wire new_Jinkela_wire_6372;
    wire new_Jinkela_wire_8415;
    wire new_Jinkela_wire_9620;
    wire new_Jinkela_wire_5451;
    wire new_Jinkela_wire_10263;
    wire new_Jinkela_wire_7040;
    wire new_Jinkela_wire_9293;
    wire new_Jinkela_wire_1943;
    wire new_Jinkela_wire_9732;
    wire new_Jinkela_wire_3475;
    wire new_Jinkela_wire_868;
    wire new_Jinkela_wire_9983;
    wire new_Jinkela_wire_924;
    wire new_Jinkela_wire_7328;
    wire new_Jinkela_wire_7256;
    wire new_Jinkela_wire_3599;
    wire new_Jinkela_wire_8338;
    wire new_Jinkela_wire_84;
    wire new_Jinkela_wire_520;
    wire new_Jinkela_wire_3781;
    wire new_Jinkela_wire_7828;
    wire new_Jinkela_wire_6872;
    wire new_Jinkela_wire_5649;
    wire new_Jinkela_wire_6665;
    wire new_Jinkela_wire_6624;
    wire new_Jinkela_wire_5926;
    wire new_Jinkela_wire_3833;
    wire new_Jinkela_wire_5703;
    wire new_Jinkela_wire_9093;
    wire new_Jinkela_wire_6098;
    wire new_Jinkela_wire_5416;
    wire new_Jinkela_wire_9299;
    wire new_Jinkela_wire_9515;
    wire new_Jinkela_wire_9604;
    wire new_Jinkela_wire_5671;
    wire new_Jinkela_wire_3947;
    wire new_Jinkela_wire_4666;
    wire n_0029_;
    wire n_0055_;
    wire new_Jinkela_wire_129;
    wire n_1243_;
    wire new_Jinkela_wire_8608;
    wire new_Jinkela_wire_7694;
    wire new_Jinkela_wire_1029;
    wire new_Jinkela_wire_777;
    wire new_Jinkela_wire_3622;
    wire new_Jinkela_wire_3367;
    wire new_Jinkela_wire_5168;
    wire new_Jinkela_wire_10115;
    wire new_Jinkela_wire_7373;
    wire new_Jinkela_wire_4275;
    wire n_1026_;
    wire new_Jinkela_wire_9825;
    wire new_Jinkela_wire_5645;
    wire new_Jinkela_wire_9996;
    wire new_Jinkela_wire_9337;
    wire n_0451_;
    wire new_Jinkela_wire_10486;
    wire new_Jinkela_wire_4728;
    wire new_Jinkela_wire_6693;
    wire new_Jinkela_wire_6492;
    wire new_Jinkela_wire_6152;
    wire new_Jinkela_wire_3340;
    wire n_1249_;
    wire new_Jinkela_wire_7634;
    wire n_1340_;
    wire new_Jinkela_wire_8053;
    wire new_Jinkela_wire_10595;
    wire new_Jinkela_wire_8658;
    wire new_Jinkela_wire_8122;
    wire new_Jinkela_wire_4075;
    wire new_Jinkela_wire_9480;
    wire new_Jinkela_wire_5765;
    wire new_Jinkela_wire_9723;
    wire new_Jinkela_wire_974;
    wire new_Jinkela_wire_8794;
    wire new_Jinkela_wire_5716;
    wire new_Jinkela_wire_3400;
    wire new_Jinkela_wire_6257;
    wire new_Jinkela_wire_564;
    wire new_Jinkela_wire_9925;
    wire new_Jinkela_wire_10409;
    wire new_Jinkela_wire_628;
    wire new_Jinkela_wire_9075;
    wire new_Jinkela_wire_4609;
    wire new_Jinkela_wire_5015;
    wire new_Jinkela_wire_5098;
    wire n_1143_;
    wire new_Jinkela_wire_9425;
    wire new_Jinkela_wire_5467;
    wire new_Jinkela_wire_6675;
    wire new_Jinkela_wire_7712;
    wire new_Jinkela_wire_2282;
    wire n_0939_;
    wire new_Jinkela_wire_1651;
    wire new_Jinkela_wire_8917;
    wire n_1064_;
    wire new_Jinkela_wire_29;
    wire new_Jinkela_wire_9172;
    wire new_Jinkela_wire_10036;
    wire new_Jinkela_wire_9170;
    wire new_Jinkela_wire_80;
    wire new_Jinkela_wire_3782;
    wire new_Jinkela_wire_6522;
    wire new_Jinkela_wire_3637;
    wire new_Jinkela_wire_4611;
    wire new_Jinkela_wire_2345;
    wire new_Jinkela_wire_8643;
    wire new_Jinkela_wire_1481;
    wire n_1156_;
    wire new_Jinkela_wire_5991;
    wire new_Jinkela_wire_3456;
    wire n_0324_;
    wire new_Jinkela_wire_6427;
    wire new_Jinkela_wire_1303;
    wire new_Jinkela_wire_3036;
    wire new_Jinkela_wire_794;
    wire n_0109_;
    wire new_Jinkela_wire_7158;
    wire new_Jinkela_wire_9926;
    wire new_Jinkela_wire_809;
    wire new_Jinkela_wire_2921;
    wire new_Jinkela_wire_1522;
    wire new_Jinkela_wire_3981;
    wire new_Jinkela_wire_3664;
    wire new_Jinkela_wire_8191;
    wire n_0281_;
    wire new_Jinkela_wire_2642;
    wire new_Jinkela_wire_8030;
    wire new_Jinkela_wire_7112;
    wire new_Jinkela_wire_6072;
    wire new_Jinkela_wire_2204;
    wire new_Jinkela_wire_3686;
    wire n_1327_;
    wire n_0095_;
    wire new_Jinkela_wire_9848;
    wire new_Jinkela_wire_2440;
    wire new_Jinkela_wire_4897;
    wire n_0929_;
    wire new_Jinkela_wire_5550;
    wire new_Jinkela_wire_3184;
    wire new_Jinkela_wire_913;
    wire new_Jinkela_wire_330;
    wire new_Jinkela_wire_6535;
    wire new_Jinkela_wire_2571;
    wire new_Jinkela_wire_4108;
    wire new_Jinkela_wire_796;
    wire new_Jinkela_wire_8409;
    wire new_Jinkela_wire_5909;
    wire new_Jinkela_wire_5647;
    wire n_0973_;
    wire new_Jinkela_wire_7901;
    wire n_0840_;
    wire new_Jinkela_wire_9603;
    wire n_1220_;
    wire new_Jinkela_wire_25;
    wire new_Jinkela_wire_6720;
    wire new_Jinkela_wire_1358;
    wire new_Jinkela_wire_709;
    wire new_Jinkela_wire_7769;
    wire new_Jinkela_wire_5770;
    wire new_Jinkela_wire_8087;
    wire new_Jinkela_wire_3629;
    wire new_Jinkela_wire_7343;
    wire new_Jinkela_wire_7085;
    wire new_Jinkela_wire_7741;
    wire new_Jinkela_wire_5389;
    wire new_Jinkela_wire_3856;
    wire new_Jinkela_wire_1397;
    wire new_Jinkela_wire_2316;
    wire new_Jinkela_wire_6106;
    wire new_Jinkela_wire_36;
    wire new_Jinkela_wire_4118;
    wire n_1137_;
    wire new_Jinkela_wire_9912;
    wire new_Jinkela_wire_9054;
    wire new_Jinkela_wire_9945;
    wire n_0563_;
    wire new_Jinkela_wire_9688;
    wire n_0282_;
    wire new_Jinkela_wire_5232;
    wire new_Jinkela_wire_4758;
    wire n_0688_;
    wire new_Jinkela_wire_6986;
    wire new_Jinkela_wire_107;
    wire n_0265_;
    wire new_Jinkela_wire_3712;
    wire new_Jinkela_wire_6884;
    wire new_Jinkela_wire_3095;
    wire new_net_12;
    wire new_Jinkela_wire_5037;
    wire new_Jinkela_wire_2324;
    wire new_Jinkela_wire_3165;
    wire new_Jinkela_wire_9700;
    wire new_Jinkela_wire_2336;
    wire new_Jinkela_wire_6293;
    wire new_Jinkela_wire_4058;
    wire new_Jinkela_wire_2301;
    wire new_Jinkela_wire_2148;
    wire new_Jinkela_wire_5509;
    wire new_Jinkela_wire_2014;
    wire new_Jinkela_wire_6460;
    wire new_Jinkela_wire_449;
    wire new_Jinkela_wire_9630;
    wire new_Jinkela_wire_9573;
    wire new_Jinkela_wire_9200;
    wire new_Jinkela_wire_2548;
    wire new_Jinkela_wire_3187;
    wire new_Jinkela_wire_8702;
    wire new_Jinkela_wire_7976;
    wire new_Jinkela_wire_1544;
    wire new_Jinkela_wire_4841;
    wire new_Jinkela_wire_6852;
    wire new_Jinkela_wire_6315;
    wire new_Jinkela_wire_4787;
    wire n_0615_;
    wire new_Jinkela_wire_10190;
    wire new_Jinkela_wire_8841;
    wire new_Jinkela_wire_538;
    wire new_Jinkela_wire_3446;
    wire new_Jinkela_wire_4669;
    wire new_Jinkela_wire_1336;
    wire n_0406_;
    wire new_Jinkela_wire_6839;
    wire new_Jinkela_wire_3251;
    wire n_0193_;
    wire new_Jinkela_wire_6615;
    wire new_Jinkela_wire_8873;
    wire new_Jinkela_wire_5286;
    wire new_Jinkela_wire_7737;
    wire new_Jinkela_wire_8396;
    wire n_0268_;
    wire new_Jinkela_wire_242;
    wire new_Jinkela_wire_607;
    wire new_Jinkela_wire_7977;
    wire new_Jinkela_wire_2775;
    wire new_Jinkela_wire_3213;
    wire new_Jinkela_wire_4468;
    wire new_Jinkela_wire_8176;
    wire new_Jinkela_wire_7143;
    wire new_Jinkela_wire_6071;
    wire new_Jinkela_wire_9935;
    wire new_Jinkela_wire_7321;
    wire new_Jinkela_wire_2543;
    wire new_Jinkela_wire_3298;
    wire new_Jinkela_wire_8599;
    wire new_Jinkela_wire_2634;
    wire new_Jinkela_wire_4827;
    wire n_0889_;
    wire new_Jinkela_wire_7711;
    wire new_Jinkela_wire_7320;
    wire new_Jinkela_wire_7151;
    wire new_Jinkela_wire_7465;
    wire new_Jinkela_wire_7388;
    wire new_Jinkela_wire_10375;
    wire new_Jinkela_wire_7507;
    wire new_Jinkela_wire_6900;
    wire new_Jinkela_wire_5640;
    wire new_Jinkela_wire_7018;
    wire new_Jinkela_wire_6537;
    wire new_Jinkela_wire_6030;
    wire new_Jinkela_wire_3445;
    wire new_Jinkela_wire_3652;
    wire new_Jinkela_wire_2939;
    wire new_Jinkela_wire_4138;
    wire new_Jinkela_wire_1250;
    wire new_Jinkela_wire_6455;
    wire new_Jinkela_wire_1511;
    wire n_0667_;
    wire new_Jinkela_wire_3476;
    wire new_Jinkela_wire_10138;
    wire new_Jinkela_wire_710;
    wire new_Jinkela_wire_7790;
    wire new_Jinkela_wire_5632;
    wire new_Jinkela_wire_1081;
    wire new_Jinkela_wire_4904;
    wire new_Jinkela_wire_8838;
    wire new_Jinkela_wire_3596;
    wire new_Jinkela_wire_6447;
    wire new_Jinkela_wire_8931;
    wire n_0925_;
    wire new_Jinkela_wire_6394;
    wire n_0762_;
    wire new_Jinkela_wire_8869;
    wire new_Jinkela_wire_5691;
    wire new_Jinkela_wire_5428;
    wire new_Jinkela_wire_7609;
    wire new_Jinkela_wire_10452;
    wire new_Jinkela_wire_3551;
    wire new_Jinkela_wire_4879;
    wire new_Jinkela_wire_6511;
    wire new_Jinkela_wire_8464;
    wire new_Jinkela_wire_1876;
    wire new_Jinkela_wire_6261;
    wire new_Jinkela_wire_9125;
    wire new_Jinkela_wire_2965;
    wire new_Jinkela_wire_4242;
    wire new_Jinkela_wire_3287;
    wire n_0798_;
    wire new_Jinkela_wire_9483;
    wire new_Jinkela_wire_1821;
    wire new_Jinkela_wire_659;
    wire new_Jinkela_wire_888;
    wire new_Jinkela_wire_4623;
    wire new_Jinkela_wire_10401;
    wire new_Jinkela_wire_7670;
    wire new_Jinkela_wire_373;
    wire new_Jinkela_wire_1410;
    wire new_Jinkela_wire_174;
    wire new_Jinkela_wire_10428;
    wire n_1150_;
    wire new_Jinkela_wire_3531;
    wire new_Jinkela_wire_5067;
    wire new_Jinkela_wire_315;
    wire new_Jinkela_wire_9932;
    wire new_Jinkela_wire_7279;
    wire new_Jinkela_wire_2152;
    wire new_Jinkela_wire_3953;
    wire new_Jinkela_wire_9253;
    wire new_Jinkela_wire_5101;
    wire new_Jinkela_wire_7724;
    wire new_Jinkela_wire_9694;
    wire new_Jinkela_wire_4042;
    wire new_Jinkela_wire_5275;
    wire new_Jinkela_wire_1703;
    wire new_Jinkela_wire_3770;
    wire new_Jinkela_wire_3495;
    wire new_Jinkela_wire_49;
    wire new_Jinkela_wire_1732;
    wire new_Jinkela_wire_7291;
    wire new_Jinkela_wire_775;
    wire new_Jinkela_wire_6670;
    wire new_Jinkela_wire_1457;
    wire new_Jinkela_wire_1666;
    wire new_Jinkela_wire_6145;
    wire new_Jinkela_wire_5975;
    wire new_Jinkela_wire_9095;
    wire new_Jinkela_wire_7280;
    wire new_Jinkela_wire_2290;
    wire new_Jinkela_wire_10234;
    wire n_0724_;
    wire new_Jinkela_wire_1530;
    wire n_0022_;
    wire new_net_2491;
    wire new_Jinkela_wire_1141;
    wire n_0057_;
    wire new_Jinkela_wire_7420;
    wire new_Jinkela_wire_6217;
    wire new_Jinkela_wire_3326;
    wire new_Jinkela_wire_5617;
    wire new_Jinkela_wire_5091;
    wire new_Jinkela_wire_7381;
    wire new_Jinkela_wire_7518;
    wire n_1084_;
    wire n_0118_;
    wire new_Jinkela_wire_3891;
    wire new_Jinkela_wire_8777;
    wire new_Jinkela_wire_9854;
    wire new_Jinkela_wire_8704;
    wire new_Jinkela_wire_10098;
    wire n_0694_;
    wire new_Jinkela_wire_2963;
    wire new_Jinkela_wire_5217;
    wire new_Jinkela_wire_3660;
    wire n_1208_;
    wire new_Jinkela_wire_9529;
    wire new_Jinkela_wire_5183;
    wire new_Jinkela_wire_2327;
    wire new_Jinkela_wire_4618;
    wire new_Jinkela_wire_867;
    wire new_Jinkela_wire_9965;
    wire new_Jinkela_wire_1929;
    wire new_Jinkela_wire_10532;
    wire new_Jinkela_wire_2919;
    wire new_Jinkela_wire_3545;
    wire new_Jinkela_wire_7226;
    wire new_Jinkela_wire_3806;
    wire new_Jinkela_wire_9083;
    wire new_Jinkela_wire_4129;
    wire new_Jinkela_wire_4216;
    wire n_0835_;
    wire new_Jinkela_wire_3588;
    wire new_Jinkela_wire_8332;
    wire new_Jinkela_wire_3621;
    wire new_Jinkela_wire_365;
    wire new_Jinkela_wire_9982;
    wire new_Jinkela_wire_2115;
    wire n_0158_;
    wire new_Jinkela_wire_5293;
    wire new_Jinkela_wire_47;
    wire new_Jinkela_wire_2763;
    wire new_Jinkela_wire_5047;
    wire new_Jinkela_wire_7866;
    wire new_Jinkela_wire_5079;
    wire new_Jinkela_wire_3737;
    wire new_Jinkela_wire_5161;
    wire n_0904_;
    wire new_Jinkela_wire_8482;
    wire new_Jinkela_wire_7799;
    wire new_Jinkela_wire_5911;
    wire new_Jinkela_wire_1435;
    wire new_Jinkela_wire_3403;
    wire new_Jinkela_wire_10092;
    wire new_Jinkela_wire_1018;
    wire new_Jinkela_wire_10546;
    wire new_Jinkela_wire_6558;
    wire new_Jinkela_wire_3988;
    wire new_Jinkela_wire_2726;
    wire new_Jinkela_wire_6577;
    wire new_Jinkela_wire_2771;
    wire new_Jinkela_wire_3923;
    wire new_Jinkela_wire_5903;
    wire n_0433_;
    wire new_Jinkela_wire_6584;
    wire n_1247_;
    wire new_Jinkela_wire_3011;
    wire new_Jinkela_wire_10574;
    wire new_Jinkela_wire_7728;
    wire new_Jinkela_wire_1151;
    wire n_1352_;
    wire n_1012_;
    wire new_Jinkela_wire_5087;
    wire new_Jinkela_wire_1296;
    wire new_Jinkela_wire_1300;
    wire new_Jinkela_wire_8443;
    wire new_Jinkela_wire_308;
    wire new_Jinkela_wire_9990;
    wire new_Jinkela_wire_8213;
    wire n_1297_;
    wire new_Jinkela_wire_2817;
    wire new_Jinkela_wire_7685;
    wire new_Jinkela_wire_1523;
    wire new_Jinkela_wire_9468;
    wire n_0379_;
    wire new_Jinkela_wire_7092;
    wire new_Jinkela_wire_5545;
    wire new_Jinkela_wire_9598;
    wire new_Jinkela_wire_5687;
    wire new_Jinkela_wire_2884;
    wire new_Jinkela_wire_4529;
    wire n_1222_;
    wire new_Jinkela_wire_1184;
    wire new_Jinkela_wire_9997;
    wire new_Jinkela_wire_10610;
    wire new_Jinkela_wire_8926;
    wire new_Jinkela_wire_8386;
    wire new_Jinkela_wire_383;
    wire new_Jinkela_wire_3452;
    wire new_Jinkela_wire_2118;
    wire n_0017_;
    wire new_Jinkela_wire_3216;
    wire new_Jinkela_wire_7560;
    wire new_Jinkela_wire_10542;
    wire new_Jinkela_wire_4700;
    wire new_Jinkela_wire_4653;
    wire new_Jinkela_wire_10492;
    wire n_1039_;
    wire new_Jinkela_wire_4176;
    wire new_Jinkela_wire_5580;
    wire new_Jinkela_wire_2515;
    wire new_Jinkela_wire_9471;
    wire new_Jinkela_wire_6696;
    wire new_Jinkela_wire_9476;
    wire new_Jinkela_wire_3879;
    wire new_Jinkela_wire_1676;
    wire new_Jinkela_wire_4067;
    wire new_Jinkela_wire_4547;
    wire new_Jinkela_wire_2468;
    wire new_Jinkela_wire_1770;
    wire new_Jinkela_wire_7425;
    wire new_Jinkela_wire_4811;
    wire new_Jinkela_wire_5417;
    wire new_Jinkela_wire_10220;
    wire new_Jinkela_wire_8051;
    wire new_Jinkela_wire_1208;
    wire n_0954_;
    wire new_Jinkela_wire_2179;
    wire new_Jinkela_wire_4014;
    wire new_Jinkela_wire_6965;
    wire new_Jinkela_wire_8428;
    wire new_Jinkela_wire_4870;
    wire new_Jinkela_wire_1962;
    wire new_Jinkela_wire_4615;
    wire new_Jinkela_wire_1842;
    wire new_Jinkela_wire_10087;
    wire new_Jinkela_wire_7726;
    wire new_Jinkela_wire_4437;
    wire new_Jinkela_wire_6911;
    wire new_Jinkela_wire_1950;
    wire new_Jinkela_wire_8470;
    wire new_Jinkela_wire_1979;
    wire n_1344_;
    wire n_0206_;
    wire new_Jinkela_wire_3172;
    wire n_0424_;
    wire new_Jinkela_wire_402;
    wire new_Jinkela_wire_6129;
    wire new_Jinkela_wire_10089;
    wire new_Jinkela_wire_7305;
    wire new_Jinkela_wire_2155;
    wire new_Jinkela_wire_8737;
    wire new_Jinkela_wire_5508;
    wire new_Jinkela_wire_4796;
    wire new_Jinkela_wire_3122;
    wire new_Jinkela_wire_7378;
    wire new_Jinkela_wire_8772;
    wire new_Jinkela_wire_2567;
    wire new_Jinkela_wire_1764;
    wire new_Jinkela_wire_4951;
    wire new_Jinkela_wire_7038;
    wire new_Jinkela_wire_3692;
    wire new_Jinkela_wire_2138;
    wire new_Jinkela_wire_9296;
    wire new_Jinkela_wire_5165;
    wire n_0553_;
    wire new_Jinkela_wire_4699;
    wire new_Jinkela_wire_6503;
    wire new_Jinkela_wire_1393;
    wire new_Jinkela_wire_2359;
    wire n_0783_;
    wire n_1278_;
    wire new_Jinkela_wire_1241;
    wire new_Jinkela_wire_749;
    wire new_Jinkela_wire_9242;
    wire new_Jinkela_wire_6714;
    wire n_0219_;
    wire new_Jinkela_wire_9386;
    wire new_Jinkela_wire_87;
    wire new_Jinkela_wire_5736;
    wire new_Jinkela_wire_6858;
    wire new_Jinkela_wire_7296;
    wire new_Jinkela_wire_10111;
    wire new_Jinkela_wire_1879;
    wire new_Jinkela_wire_8268;
    wire new_Jinkela_wire_6175;
    wire new_Jinkela_wire_7856;
    wire new_Jinkela_wire_2766;
    wire n_1218_;
    wire new_Jinkela_wire_6666;
    wire new_Jinkela_wire_9648;
    wire new_Jinkela_wire_6813;
    wire new_Jinkela_wire_9883;
    wire new_Jinkela_wire_9340;
    wire new_Jinkela_wire_1694;
    wire new_Jinkela_wire_8946;
    wire new_Jinkela_wire_1074;
    wire n_1356_;
    wire n_0292_;
    wire new_Jinkela_wire_2648;
    wire new_Jinkela_wire_5887;
    wire new_Jinkela_wire_3742;
    wire new_Jinkela_wire_2778;
    wire new_Jinkela_wire_6941;
    wire new_Jinkela_wire_2299;
    wire new_Jinkela_wire_7819;
    wire new_Jinkela_wire_1113;
    wire new_Jinkela_wire_3149;
    wire new_Jinkela_wire_8152;
    wire n_0167_;
    wire n_1008_;
    wire new_Jinkela_wire_8670;
    wire new_Jinkela_wire_8649;
    wire n_0895_;
    wire n_0245_;
    wire n_1000_;
    wire new_Jinkela_wire_257;
    wire new_Jinkela_wire_1649;
    wire new_Jinkela_wire_3572;
    wire new_Jinkela_wire_9794;
    wire new_Jinkela_wire_1211;
    wire n_0370_;
    wire new_Jinkela_wire_7550;
    wire new_Jinkela_wire_4689;
    wire new_Jinkela_wire_9279;
    wire new_Jinkela_wire_4952;
    wire new_Jinkela_wire_7431;
    wire new_Jinkela_wire_4773;
    wire new_Jinkela_wire_6792;
    wire new_Jinkela_wire_6917;
    wire new_Jinkela_wire_1445;
    wire new_Jinkela_wire_6416;
    wire new_Jinkela_wire_5319;
    wire new_Jinkela_wire_681;
    wire new_Jinkela_wire_4871;
    wire new_Jinkela_wire_661;
    wire new_Jinkela_wire_2365;
    wire n_0538_;
    wire new_Jinkela_wire_4548;
    wire new_Jinkela_wire_9721;
    wire n_0204_;
    wire new_Jinkela_wire_265;
    wire new_Jinkela_wire_773;
    wire new_Jinkela_wire_1656;
    wire new_Jinkela_wire_742;
    wire new_Jinkela_wire_292;
    wire new_Jinkela_wire_9002;
    wire new_Jinkela_wire_6528;
    wire new_Jinkela_wire_4863;
    wire new_Jinkela_wire_2643;
    wire new_Jinkela_wire_1932;
    wire new_Jinkela_wire_4276;
    wire new_Jinkela_wire_8752;
    wire new_Jinkela_wire_4837;
    wire new_Jinkela_wire_1927;
    wire new_Jinkela_wire_5979;
    wire new_Jinkela_wire_9338;
    wire new_Jinkela_wire_10355;
    wire new_Jinkela_wire_972;
    wire new_Jinkela_wire_6229;
    wire new_Jinkela_wire_10283;
    wire new_Jinkela_wire_5110;
    wire new_Jinkela_wire_1509;
    wire new_Jinkela_wire_8042;
    wire new_Jinkela_wire_8703;
    wire new_Jinkela_wire_4685;
    wire n_0743_;
    wire new_Jinkela_wire_3875;
    wire new_Jinkela_wire_9763;
    wire new_Jinkela_wire_4739;
    wire n_0350_;
    wire new_Jinkela_wire_5413;
    wire new_Jinkela_wire_3612;
    wire new_Jinkela_wire_790;
    wire new_Jinkela_wire_16;
    wire new_Jinkela_wire_1487;
    wire new_Jinkela_wire_425;
    wire n_1042_;
    wire new_Jinkela_wire_3385;
    wire new_Jinkela_wire_10478;
    wire new_Jinkela_wire_8002;
    wire new_Jinkela_wire_4613;
    wire new_Jinkela_wire_4391;
    wire new_Jinkela_wire_5818;
    wire new_Jinkela_wire_285;
    wire new_Jinkela_wire_2461;
    wire new_Jinkela_wire_4266;
    wire new_Jinkela_wire_9695;
    wire new_Jinkela_wire_1180;
    wire new_Jinkela_wire_7777;
    wire n_0135_;
    wire new_Jinkela_wire_3680;
    wire new_Jinkela_wire_4973;
    wire n_0697_;
    wire new_Jinkela_wire_7148;
    wire new_Jinkela_wire_5799;
    wire n_0423_;
    wire new_Jinkela_wire_3544;
    wire new_Jinkela_wire_3954;
    wire new_Jinkela_wire_1599;
    wire new_Jinkela_wire_2702;
    wire new_Jinkela_wire_10255;
    wire n_0883_;
    wire new_Jinkela_wire_9403;
    wire new_Jinkela_wire_3119;
    wire new_Jinkela_wire_234;
    wire new_Jinkela_wire_4393;
    wire new_Jinkela_wire_6703;
    wire new_Jinkela_wire_2930;
    wire new_Jinkela_wire_629;
    wire new_Jinkela_wire_6993;
    wire new_Jinkela_wire_2566;
    wire new_Jinkela_wire_8962;
    wire new_Jinkela_wire_2309;
    wire new_Jinkela_wire_7580;
    wire new_Jinkela_wire_2645;
    wire new_Jinkela_wire_4843;
    wire new_Jinkela_wire_9972;
    wire new_Jinkela_wire_524;
    wire new_Jinkela_wire_3881;
    wire n_0495_;
    wire new_Jinkela_wire_9761;
    wire new_Jinkela_wire_6983;
    wire new_Jinkela_wire_1042;
    wire new_Jinkela_wire_9241;
    wire n_0787_;
    wire new_Jinkela_wire_7457;
    wire n_0602_;
    wire new_Jinkela_wire_1930;
    wire new_Jinkela_wire_2993;
    wire new_Jinkela_wire_2103;
    wire new_Jinkela_wire_10265;
    wire new_Jinkela_wire_854;
    wire new_Jinkela_wire_5872;
    wire new_Jinkela_wire_1043;
    wire new_Jinkela_wire_7046;
    wire new_Jinkela_wire_5705;
    wire new_Jinkela_wire_7082;
    wire new_Jinkela_wire_6220;
    wire n_0100_;
    wire new_Jinkela_wire_1578;
    wire new_Jinkela_wire_7089;
    wire new_Jinkela_wire_4168;
    wire new_Jinkela_wire_3401;
    wire new_Jinkela_wire_5823;
    wire n_1197_;
    wire new_Jinkela_wire_4460;
    wire new_Jinkela_wire_10596;
    wire new_Jinkela_wire_6816;
    wire new_Jinkela_wire_2705;
    wire new_Jinkela_wire_182;
    wire new_Jinkela_wire_519;
    wire new_Jinkela_wire_7523;
    wire new_Jinkela_wire_445;
    wire new_Jinkela_wire_5951;
    wire new_Jinkela_wire_2426;
    wire new_Jinkela_wire_7865;
    wire new_Jinkela_wire_7078;
    wire new_Jinkela_wire_9110;
    wire n_1152_;
    wire new_Jinkela_wire_2123;
    wire new_Jinkela_wire_2311;
    wire new_Jinkela_wire_5063;
    wire new_Jinkela_wire_2927;
    wire n_0916_;
    wire new_Jinkela_wire_3971;
    wire n_1147_;
    wire new_Jinkela_wire_9236;
    wire n_0623_;
    wire new_Jinkela_wire_2717;
    wire new_Jinkela_wire_9019;
    wire new_Jinkela_wire_6380;
    wire new_Jinkela_wire_916;
    wire new_Jinkela_wire_6113;
    wire n_1272_;
    wire new_Jinkela_wire_6140;
    wire new_Jinkela_wire_10509;
    wire new_Jinkela_wire_10301;
    wire n_0717_;
    wire new_Jinkela_wire_171;
    wire new_Jinkela_wire_768;
    wire new_Jinkela_wire_1510;
    wire new_Jinkela_wire_912;
    wire new_Jinkela_wire_1176;
    wire new_Jinkela_wire_5018;
    wire n_1364_;
    wire new_Jinkela_wire_2804;
    wire new_Jinkela_wire_2402;
    wire new_Jinkela_wire_278;
    wire new_Jinkela_wire_122;
    wire new_Jinkela_wire_2628;
    wire new_Jinkela_wire_10579;
    wire new_Jinkela_wire_6343;
    wire new_Jinkela_wire_4149;
    wire new_Jinkela_wire_4289;
    wire new_Jinkela_wire_175;
    wire new_Jinkela_wire_1582;
    wire new_Jinkela_wire_1146;
    wire new_Jinkela_wire_4646;
    wire new_Jinkela_wire_3478;
    wire new_Jinkela_wire_5254;
    wire new_Jinkela_wire_7600;
    wire n_0498_;
    wire new_Jinkela_wire_10568;
    wire new_Jinkela_wire_6540;
    wire n_1180_;
    wire new_Jinkela_wire_1309;
    wire n_1028_;
    wire new_Jinkela_wire_3759;
    wire new_Jinkela_wire_4807;
    wire new_Jinkela_wire_4139;
    wire n_0541_;
    wire new_Jinkela_wire_7480;
    wire new_Jinkela_wire_2489;
    wire new_Jinkela_wire_6938;
    wire new_Jinkela_wire_5549;
    wire new_Jinkela_wire_2658;
    wire new_Jinkela_wire_787;
    wire new_Jinkela_wire_3600;
    wire new_Jinkela_wire_7332;
    wire new_Jinkela_wire_1016;
    wire new_Jinkela_wire_8765;
    wire new_Jinkela_wire_4309;
    wire new_Jinkela_wire_2610;
    wire new_Jinkela_wire_8922;
    wire new_Jinkela_wire_3948;
    wire new_Jinkela_wire_2051;
    wire new_Jinkela_wire_920;
    wire new_Jinkela_wire_10069;
    wire new_Jinkela_wire_3837;
    wire new_Jinkela_wire_4894;
    wire new_Jinkela_wire_951;
    wire new_Jinkela_wire_1038;
    wire new_Jinkela_wire_10353;
    wire new_Jinkela_wire_4891;
    wire new_Jinkela_wire_3424;
    wire new_Jinkela_wire_10070;
    wire n_0839_;
    wire new_Jinkela_wire_2631;
    wire new_Jinkela_wire_1854;
    wire new_Jinkela_wire_9404;
    wire n_0987_;
    wire new_Jinkela_wire_694;
    wire new_Jinkela_wire_5334;
    wire new_Jinkela_wire_7682;
    wire new_Jinkela_wire_6582;
    wire n_0266_;
    wire new_Jinkela_wire_889;
    wire new_Jinkela_wire_3275;
    wire new_Jinkela_wire_10553;
    wire new_Jinkela_wire_3691;
    wire new_Jinkela_wire_4239;
    wire new_Jinkela_wire_714;
    wire n_1113_;
    wire new_Jinkela_wire_9510;
    wire new_Jinkela_wire_7098;
    wire new_Jinkela_wire_9508;
    wire new_Jinkela_wire_2793;
    wire new_Jinkela_wire_1060;
    wire new_Jinkela_wire_4744;
    wire new_Jinkela_wire_2158;
    wire new_Jinkela_wire_4127;
    wire new_Jinkela_wire_7072;
    wire new_Jinkela_wire_1345;
    wire new_Jinkela_wire_509;
    wire new_Jinkela_wire_9360;
    wire new_Jinkela_wire_7529;
    wire new_Jinkela_wire_4893;
    wire new_Jinkela_wire_323;
    wire new_Jinkela_wire_7596;
    wire new_Jinkela_wire_325;
    wire new_Jinkela_wire_7870;
    wire new_Jinkela_wire_3315;
    wire new_Jinkela_wire_8969;
    wire new_Jinkela_wire_6763;
    wire new_Jinkela_wire_7883;
    wire new_net_1;
    wire new_Jinkela_wire_10304;
    wire n_0103_;
    wire new_Jinkela_wire_621;
    wire new_Jinkela_wire_7099;
    wire new_Jinkela_wire_10154;
    wire new_Jinkela_wire_8771;
    wire new_Jinkela_wire_34;
    wire n_1009_;
    wire new_Jinkela_wire_231;
    wire new_Jinkela_wire_6853;
    wire new_Jinkela_wire_7252;
    wire new_Jinkela_wire_957;
    wire n_0871_;
    wire new_Jinkela_wire_6601;
    wire new_Jinkela_wire_3083;
    wire new_Jinkela_wire_8810;
    wire new_Jinkela_wire_4235;
    wire new_Jinkela_wire_2759;
    wire new_Jinkela_wire_5492;
    wire new_Jinkela_wire_6269;
    wire new_Jinkela_wire_10134;
    wire new_Jinkela_wire_1834;
    wire new_Jinkela_wire_5588;
    wire new_Jinkela_wire_9724;
    wire new_Jinkela_wire_1559;
    wire new_Jinkela_wire_266;
    wire new_Jinkela_wire_5675;
    wire new_Jinkela_wire_9699;
    wire n_0693_;
    wire new_Jinkela_wire_8533;
    wire n_0748_;
    wire new_Jinkela_wire_6468;
    wire new_Jinkela_wire_660;
    wire new_Jinkela_wire_4537;
    wire new_Jinkela_wire_3920;
    wire new_Jinkela_wire_10141;
    wire new_Jinkela_wire_2428;
    wire new_Jinkela_wire_5003;
    wire new_Jinkela_wire_859;
    wire new_Jinkela_wire_6267;
    wire new_Jinkela_wire_3441;
    wire new_Jinkela_wire_2340;
    wire new_Jinkela_wire_10427;
    wire new_Jinkela_wire_194;
    wire new_Jinkela_wire_3280;
    wire new_Jinkela_wire_5274;
    wire new_Jinkela_wire_428;
    wire new_Jinkela_wire_9470;
    wire new_Jinkela_wire_8469;
    wire new_Jinkela_wire_21;
    wire new_Jinkela_wire_7045;
    wire new_Jinkela_wire_9092;
    wire new_Jinkela_wire_3196;
    wire new_Jinkela_wire_8983;
    wire new_Jinkela_wire_3915;
    wire new_Jinkela_wire_1367;
    wire new_Jinkela_wire_3047;
    wire new_Jinkela_wire_6871;
    wire new_Jinkela_wire_3496;
    wire new_Jinkela_wire_6040;
    wire new_Jinkela_wire_8745;
    wire new_Jinkela_wire_4051;
    wire new_Jinkela_wire_6393;
    wire new_Jinkela_wire_8047;
    wire new_Jinkela_wire_5918;
    wire new_Jinkela_wire_7277;
    wire new_Jinkela_wire_7687;
    wire new_Jinkela_wire_3328;
    wire new_Jinkela_wire_650;
    wire new_Jinkela_wire_7615;
    wire new_Jinkela_wire_1538;
    wire new_Jinkela_wire_8335;
    wire new_Jinkela_wire_3536;
    wire new_Jinkela_wire_4238;
    wire new_Jinkela_wire_4682;
    wire new_Jinkela_wire_9856;
    wire new_Jinkela_wire_4457;
    wire new_Jinkela_wire_6700;
    wire n_0387_;
    wire new_Jinkela_wire_5267;
    wire new_Jinkela_wire_8719;
    wire new_Jinkela_wire_7456;
    wire new_Jinkela_wire_7891;
    wire new_Jinkela_wire_7481;
    wire new_Jinkela_wire_7699;
    wire new_Jinkela_wire_3624;
    wire new_Jinkela_wire_8660;
    wire new_Jinkela_wire_9586;
    wire new_Jinkela_wire_5159;
    wire new_Jinkela_wire_8126;
    wire new_Jinkela_wire_2984;
    wire new_Jinkela_wire_4735;
    wire new_Jinkela_wire_6171;
    wire new_Jinkela_wire_4417;
    wire new_Jinkela_wire_6962;
    wire new_Jinkela_wire_7073;
    wire n_1191_;
    wire new_Jinkela_wire_5553;
    wire new_Jinkela_wire_1976;
    wire new_Jinkela_wire_8372;
    wire new_Jinkela_wire_6516;
    wire new_Jinkela_wire_6604;
    wire new_Jinkela_wire_9052;
    wire new_Jinkela_wire_2279;
    wire new_Jinkela_wire_6600;
    wire n_0083_;
    wire new_Jinkela_wire_10589;
    wire new_Jinkela_wire_81;
    wire new_Jinkela_wire_355;
    wire new_Jinkela_wire_5581;
    wire new_Jinkela_wire_2221;
    wire new_Jinkela_wire_9934;
    wire new_Jinkela_wire_1073;
    wire n_0828_;
    wire new_Jinkela_wire_7121;
    wire new_Jinkela_wire_3230;
    wire new_Jinkela_wire_3949;
    wire new_Jinkela_wire_5350;
    wire new_Jinkela_wire_9727;
    wire new_Jinkela_wire_4915;
    wire n_0974_;
    wire new_Jinkela_wire_929;
    wire new_Jinkela_wire_6599;
    wire new_Jinkela_wire_679;
    wire new_Jinkela_wire_7064;
    wire new_Jinkela_wire_10302;
    wire new_Jinkela_wire_7188;
    wire new_Jinkela_wire_9764;
    wire new_Jinkela_wire_5042;
    wire n_0990_;
    wire new_Jinkela_wire_10028;
    wire new_Jinkela_wire_8105;
    wire new_Jinkela_wire_5090;
    wire new_Jinkela_wire_4523;
    wire n_1273_;
    wire new_Jinkela_wire_5128;
    wire new_Jinkela_wire_4605;
    wire new_Jinkela_wire_5698;
    wire new_Jinkela_wire_1246;
    wire new_Jinkela_wire_10373;
    wire new_Jinkela_wire_4936;
    wire new_Jinkela_wire_7412;
    wire new_Jinkela_wire_10011;
    wire new_Jinkela_wire_9462;
    wire new_Jinkela_wire_10369;
    wire new_Jinkela_wire_6832;
    wire new_Jinkela_wire_2078;
    wire new_Jinkela_wire_2246;
    wire new_Jinkela_wire_2369;
    wire n_0986_;
    wire new_Jinkela_wire_8577;
    wire new_Jinkela_wire_7656;
    wire new_Jinkela_wire_4512;
    wire new_Jinkela_wire_4054;
    wire new_Jinkela_wire_6612;
    wire new_Jinkela_wire_5265;
    wire new_Jinkela_wire_6247;
    wire new_Jinkela_wire_9777;
    wire new_Jinkela_wire_5594;
    wire new_Jinkela_wire_3662;
    wire new_Jinkela_wire_2154;
    wire new_Jinkela_wire_8855;
    wire new_Jinkela_wire_8604;
    wire new_Jinkela_wire_5768;
    wire new_Jinkela_wire_7307;
    wire new_Jinkela_wire_6877;
    wire new_Jinkela_wire_6723;
    wire new_Jinkela_wire_908;
    wire new_Jinkela_wire_9670;
    wire new_Jinkela_wire_3365;
    wire new_Jinkela_wire_8098;
    wire new_Jinkela_wire_10631;
    wire new_Jinkela_wire_4406;
    wire new_Jinkela_wire_361;
    wire new_Jinkela_wire_3186;
    wire new_Jinkela_wire_8914;
    wire new_Jinkela_wire_7809;
    wire new_Jinkela_wire_4454;
    wire new_Jinkela_wire_1344;
    wire new_Jinkela_wire_7618;
    wire new_Jinkela_wire_9452;
    wire new_Jinkela_wire_835;
    wire new_Jinkela_wire_1420;
    wire n_0209_;
    wire new_Jinkela_wire_6474;
    wire n_0777_;
    wire new_Jinkela_wire_6400;
    wire new_Jinkela_wire_6410;
    wire n_1002_;
    wire new_Jinkela_wire_1107;
    wire new_Jinkela_wire_6219;
    wire new_Jinkela_wire_1812;
    wire new_Jinkela_wire_2441;
    wire new_Jinkela_wire_6282;
    wire n_1101_;
    wire new_Jinkela_wire_1820;
    wire new_Jinkela_wire_8834;
    wire new_Jinkela_wire_5230;
    wire new_Jinkela_wire_1543;
    wire new_Jinkela_wire_10396;
    wire new_Jinkela_wire_7117;
    wire new_Jinkela_wire_1850;
    wire new_Jinkela_wire_10321;
    wire new_Jinkela_wire_2676;
    wire new_Jinkela_wire_4003;
    wire new_Jinkela_wire_9008;
    wire new_Jinkela_wire_6953;
    wire new_Jinkela_wire_1476;
    wire new_Jinkela_wire_9702;
    wire new_Jinkela_wire_204;
    wire new_Jinkela_wire_6589;
    wire new_Jinkela_wire_10150;
    wire new_Jinkela_wire_510;
    wire new_Jinkela_wire_5137;
    wire new_Jinkela_wire_9017;
    wire new_Jinkela_wire_7684;
    wire n_0226_;
    wire new_Jinkela_wire_4886;
    wire new_Jinkela_wire_934;
    wire new_Jinkela_wire_4809;
    wire new_Jinkela_wire_4764;
    wire new_Jinkela_wire_1385;
    wire new_Jinkela_wire_9157;
    wire new_Jinkela_wire_4146;
    wire new_Jinkela_wire_5829;
    wire new_Jinkela_wire_6767;
    wire new_Jinkela_wire_9845;
    wire new_Jinkela_wire_3414;
    wire n_0978_;
    wire new_Jinkela_wire_1969;
    wire n_0050_;
    wire n_0535_;
    wire new_Jinkela_wire_7924;
    wire new_Jinkela_wire_933;
    wire new_Jinkela_wire_1597;
    wire new_Jinkela_wire_1424;
    wire new_Jinkela_wire_4719;
    wire new_Jinkela_wire_6651;
    wire new_Jinkela_wire_4491;
    wire new_Jinkela_wire_3402;
    wire n_0567_;
    wire new_Jinkela_wire_2850;
    wire new_Jinkela_wire_4544;
    wire new_Jinkela_wire_5621;
    wire new_Jinkela_wire_7096;
    wire new_Jinkela_wire_1558;
    wire new_Jinkela_wire_5140;
    wire new_Jinkela_wire_7270;
    wire new_Jinkela_wire_5487;
    wire new_Jinkela_wire_4132;
    wire new_Jinkela_wire_10533;
    wire new_Jinkela_wire_6886;
    wire new_Jinkela_wire_9832;
    wire new_Jinkela_wire_5372;
    wire new_Jinkela_wire_9866;
    wire n_1096_;
    wire new_Jinkela_wire_5378;
    wire new_Jinkela_wire_1968;
    wire new_Jinkela_wire_55;
    wire new_Jinkela_wire_3197;
    wire new_Jinkela_wire_7290;
    wire new_Jinkela_wire_1324;
    wire new_Jinkela_wire_5419;
    wire new_Jinkela_wire_9276;
    wire new_Jinkela_wire_7941;
    wire new_Jinkela_wire_6697;
    wire new_Jinkela_wire_574;
    wire new_Jinkela_wire_10451;
    wire n_0330_;
    wire new_Jinkela_wire_4423;
    wire new_Jinkela_wire_4557;
    wire new_Jinkela_wire_1245;
    wire n_1271_;
    wire new_Jinkela_wire_2015;
    wire new_Jinkela_wire_3265;
    wire new_Jinkela_wire_1415;
    wire new_Jinkela_wire_5307;
    wire new_Jinkela_wire_2116;
    wire new_Jinkela_wire_8930;
    wire new_Jinkela_wire_5463;
    wire new_Jinkela_wire_1268;
    wire new_Jinkela_wire_9341;
    wire new_Jinkela_wire_8879;
    wire new_Jinkela_wire_2773;
    wire new_Jinkela_wire_7079;
    wire new_Jinkela_wire_570;
    wire new_Jinkela_wire_5743;
    wire new_Jinkela_wire_3144;
    wire new_Jinkela_wire_7127;
    wire new_Jinkela_wire_2133;
    wire new_Jinkela_wire_3178;
    wire new_Jinkela_wire_4924;
    wire new_Jinkela_wire_4175;
    wire new_Jinkela_wire_6552;
    wire new_Jinkela_wire_7124;
    wire new_Jinkela_wire_8024;
    wire new_Jinkela_wire_10620;
    wire new_Jinkela_wire_6003;
    wire new_Jinkela_wire_4434;
    wire new_Jinkela_wire_6637;
    wire new_Jinkela_wire_523;
    wire new_Jinkela_wire_6231;
    wire new_Jinkela_wire_5083;
    wire new_Jinkela_wire_3301;
    wire n_0923_;
    wire new_Jinkela_wire_5625;
    wire new_Jinkela_wire_4416;
    wire new_Jinkela_wire_685;
    wire new_Jinkela_wire_5466;
    wire new_Jinkela_wire_609;
    wire n_0967_;
    wire new_Jinkela_wire_3131;
    wire new_Jinkela_wire_8954;
    wire n_0902_;
    wire new_Jinkela_wire_10145;
    wire new_Jinkela_wire_5270;
    wire new_Jinkela_wire_1228;
    wire n_0874_;
    wire new_Jinkela_wire_7989;
    wire new_Jinkela_wire_5830;
    wire n_1148_;
    wire new_Jinkela_wire_9795;
    wire new_Jinkela_wire_5046;
    wire new_Jinkela_wire_3513;
    wire new_Jinkela_wire_5816;
    wire new_Jinkela_wire_10431;
    wire new_Jinkela_wire_6726;
    wire new_Jinkela_wire_8579;
    wire new_Jinkela_wire_10019;
    wire new_Jinkela_wire_1178;
    wire new_Jinkela_wire_847;
    wire new_Jinkela_wire_711;
    wire new_Jinkela_wire_2709;
    wire n_0523_;
    wire new_Jinkela_wire_3269;
    wire new_Jinkela_wire_2338;
    wire new_Jinkela_wire_8340;
    wire new_Jinkela_wire_2891;
    wire new_Jinkela_wire_6346;
    wire new_Jinkela_wire_2478;
    wire new_Jinkela_wire_1441;
    wire new_Jinkela_wire_1882;
    wire n_0515_;
    wire new_Jinkela_wire_8999;
    wire new_Jinkela_wire_4990;
    wire new_Jinkela_wire_1277;
    wire new_Jinkela_wire_975;
    wire n_0505_;
    wire n_0859_;
    wire new_Jinkela_wire_9629;
    wire new_Jinkela_wire_5760;
    wire n_0390_;
    wire new_Jinkela_wire_1103;
    wire new_Jinkela_wire_1555;
    wire new_Jinkela_wire_8957;
    wire new_Jinkela_wire_2995;
    wire new_Jinkela_wire_71;
    wire new_Jinkela_wire_4910;
    wire new_Jinkela_wire_4145;
    wire new_Jinkela_wire_4380;
    wire new_Jinkela_wire_243;
    wire new_Jinkela_wire_4436;
    wire new_Jinkela_wire_3253;
    wire new_Jinkela_wire_4500;
    wire new_Jinkela_wire_4817;
    wire n_0077_;
    wire new_Jinkela_wire_7356;
    wire new_Jinkela_wire_5967;
    wire new_Jinkela_wire_140;
    wire new_Jinkela_wire_9719;
    wire new_Jinkela_wire_8190;
    wire new_Jinkela_wire_8435;
    wire new_Jinkela_wire_2698;
    wire new_Jinkela_wire_310;
    wire new_Jinkela_wire_10565;
    wire new_Jinkela_wire_5283;
    wire new_Jinkela_wire_1569;
    wire new_Jinkela_wire_5066;
    wire n_0240_;
    wire new_Jinkela_wire_17;
    wire n_0662_;
    wire new_Jinkela_wire_3792;
    wire n_0737_;
    wire n_0961_;
    wire new_Jinkela_wire_7855;
    wire new_Jinkela_wire_10615;
    wire new_Jinkela_wire_1760;
    wire new_Jinkela_wire_5355;
    wire new_Jinkela_wire_7495;
    wire n_0429_;
    wire n_0327_;
    wire new_Jinkela_wire_4455;
    wire new_Jinkela_wire_7608;
    wire new_Jinkela_wire_979;
    wire new_Jinkela_wire_9142;
    wire new_Jinkela_wire_1068;
    wire new_Jinkela_wire_2944;
    wire new_Jinkela_wire_5181;
    wire new_Jinkela_wire_783;
    wire new_Jinkela_wire_535;
    wire new_Jinkela_wire_3229;
    wire new_Jinkela_wire_7595;
    wire n_0631_;
    wire new_Jinkela_wire_1653;
    wire new_Jinkela_wire_3921;
    wire new_Jinkela_wire_3397;
    wire new_Jinkela_wire_2606;
    wire new_Jinkela_wire_8016;
    wire new_Jinkela_wire_7754;
    wire n_0421_;
    wire new_Jinkela_wire_2991;
    wire new_Jinkela_wire_738;
    wire new_Jinkela_wire_1997;
    wire new_Jinkela_wire_3751;
    wire new_Jinkela_wire_10012;
    wire new_Jinkela_wire_3259;
    wire n_0019_;
    wire new_Jinkela_wire_4679;
    wire new_Jinkela_wire_6555;
    wire n_0876_;
    wire new_Jinkela_wire_4651;
    wire new_Jinkela_wire_1224;
    wire new_Jinkela_wire_4822;
    wire new_Jinkela_wire_9554;
    wire new_Jinkela_wire_4039;
    wire new_Jinkela_wire_5342;
    wire n_0554_;
    wire new_Jinkela_wire_896;
    wire new_Jinkela_wire_6291;
    wire new_Jinkela_wire_9372;
    wire n_1244_;
    wire new_Jinkela_wire_9098;
    wire new_Jinkela_wire_7354;
    wire new_Jinkela_wire_7421;
    wire new_Jinkela_wire_7666;
    wire new_Jinkela_wire_2484;
    wire new_Jinkela_wire_377;
    wire n_0646_;
    wire new_Jinkela_wire_8297;
    wire new_Jinkela_wire_8528;
    wire new_Jinkela_wire_1448;
    wire n_0307_;
    wire new_Jinkela_wire_9835;
    wire new_Jinkela_wire_4151;
    wire new_Jinkela_wire_3827;
    wire new_Jinkela_wire_5941;
    wire new_Jinkela_wire_8131;
    wire new_Jinkela_wire_342;
    wire new_Jinkela_wire_2886;
    wire new_Jinkela_wire_6270;
    wire new_Jinkela_wire_1202;
    wire new_Jinkela_wire_5266;
    wire new_Jinkela_wire_8333;
    wire n_0241_;
    wire new_Jinkela_wire_491;
    wire new_Jinkela_wire_6542;
    wire new_Jinkela_wire_8390;
    wire new_Jinkela_wire_4179;
    wire n_0870_;
    wire n_0453_;
    wire n_1175_;
    wire new_Jinkela_wire_8647;
    wire new_Jinkela_wire_9010;
    wire new_Jinkela_wire_9410;
    wire new_Jinkela_wire_3907;
    wire new_Jinkela_wire_10333;
    wire new_Jinkela_wire_1075;
    wire new_Jinkela_wire_3635;
    wire new_Jinkela_wire_1039;
    wire new_Jinkela_wire_936;
    wire new_Jinkela_wire_8902;
    wire new_Jinkela_wire_1647;
    wire n_0313_;
    wire new_Jinkela_wire_1002;
    wire new_Jinkela_wire_438;
    wire new_Jinkela_wire_4632;
    wire new_Jinkela_wire_4596;
    wire new_Jinkela_wire_6348;
    wire n_1105_;
    wire new_Jinkela_wire_9927;
    wire new_Jinkela_wire_8611;
    wire new_Jinkela_wire_10599;
    wire new_Jinkela_wire_9536;
    wire new_Jinkela_wire_1174;
    wire new_Jinkela_wire_7530;
    wire new_Jinkela_wire_6920;
    wire n_0605_;
    wire new_Jinkela_wire_10269;
    wire new_Jinkela_wire_7802;
    wire n_0398_;
    wire new_Jinkela_wire_3135;
    wire new_Jinkela_wire_9678;
    wire new_Jinkela_wire_4670;
    wire new_Jinkela_wire_1248;
    wire new_Jinkela_wire_3945;
    wire new_Jinkela_wire_1777;
    wire n_0584_;
    wire new_Jinkela_wire_8416;
    wire new_Jinkela_wire_9802;
    wire new_Jinkela_wire_550;
    wire new_Jinkela_wire_4562;
    wire new_Jinkela_wire_10053;
    wire new_Jinkela_wire_1525;
    wire new_Jinkela_wire_857;
    wire new_Jinkela_wire_7342;
    wire new_Jinkela_wire_9931;
    wire new_Jinkela_wire_3429;
    wire new_Jinkela_wire_319;
    wire new_Jinkela_wire_5711;
    wire new_Jinkela_wire_8591;
    wire new_Jinkela_wire_1013;
    wire new_Jinkela_wire_784;
    wire new_Jinkela_wire_4825;
    wire new_Jinkela_wire_10587;
    wire new_Jinkela_wire_332;
    wire new_Jinkela_wire_5299;
    wire new_Jinkela_wire_3439;
    wire new_Jinkela_wire_10564;
    wire n_0420_;
    wire n_0180_;
    wire new_Jinkela_wire_7632;
    wire new_Jinkela_wire_9492;
    wire new_Jinkela_wire_10253;
    wire new_Jinkela_wire_6755;
    wire new_Jinkela_wire_740;
    wire new_Jinkela_wire_7019;
    wire new_Jinkela_wire_358;
    wire n_0125_;
    wire n_0711_;
    wire new_Jinkela_wire_10202;
    wire new_Jinkela_wire_8846;
    wire n_1221_;
    wire new_Jinkela_wire_5614;
    wire new_Jinkela_wire_9986;
    wire new_Jinkela_wire_8455;
    wire new_Jinkela_wire_8109;
    wire new_Jinkela_wire_7472;
    wire new_Jinkela_wire_5310;
    wire new_Jinkela_wire_5318;
    wire new_Jinkela_wire_573;
    wire new_Jinkela_wire_6539;
    wire new_Jinkela_wire_2466;
    wire new_Jinkela_wire_5058;
    wire new_Jinkela_wire_8874;
    wire new_Jinkela_wire_2559;
    wire new_Jinkela_wire_4370;
    wire new_Jinkela_wire_633;
    wire new_Jinkela_wire_3818;
    wire new_Jinkela_wire_9918;
    wire new_Jinkela_wire_5646;
    wire new_Jinkela_wire_67;
    wire new_Jinkela_wire_2331;
    wire new_Jinkela_wire_1091;
    wire new_Jinkela_wire_8006;
    wire new_Jinkela_wire_7177;
    wire new_Jinkela_wire_5053;
    wire new_Jinkela_wire_7325;
    wire new_Jinkela_wire_6125;
    wire new_Jinkela_wire_6623;
    wire new_Jinkela_wire_10108;
    wire new_Jinkela_wire_1809;
    wire n_0229_;
    wire n_1043_;
    wire new_Jinkela_wire_7384;
    wire new_Jinkela_wire_1589;
    wire new_Jinkela_wire_1201;
    wire new_Jinkela_wire_3029;
    wire new_Jinkela_wire_1453;
    wire new_Jinkela_wire_8974;
    wire new_Jinkela_wire_2561;
    wire new_Jinkela_wire_7007;
    wire new_Jinkela_wire_3395;
    wire new_Jinkela_wire_5568;
    wire new_Jinkela_wire_9708;
    wire new_Jinkela_wire_10278;
    wire new_Jinkela_wire_1321;
    wire new_Jinkela_wire_3880;
    wire new_Jinkela_wire_8708;
    wire new_Jinkela_wire_6235;
    wire n_0346_;
    wire n_1159_;
    wire new_Jinkela_wire_4133;
    wire new_Jinkela_wire_8744;
    wire new_Jinkela_wire_7833;
    wire n_0409_;
    wire new_Jinkela_wire_3069;
    wire new_Jinkela_wire_10132;
    wire new_Jinkela_wire_6475;
    wire new_Jinkela_wire_9243;
    wire n_0160_;
    wire new_Jinkela_wire_5860;
    wire new_Jinkela_wire_4207;
    wire n_0273_;
    wire new_Jinkela_wire_9197;
    wire new_Jinkela_wire_2972;
    wire n_1186_;
    wire new_Jinkela_wire_8592;
    wire new_Jinkela_wire_9893;
    wire new_Jinkela_wire_5812;
    wire new_Jinkela_wire_4461;
    wire new_Jinkela_wire_6027;
    wire new_Jinkela_wire_6252;
    wire new_Jinkela_wire_2367;
    wire new_Jinkela_wire_10317;
    wire new_Jinkela_wire_5022;
    wire new_Jinkela_wire_8754;
    wire new_Jinkela_wire_2738;
    wire new_Jinkela_wire_3684;
    wire new_Jinkela_wire_10543;
    wire n_0508_;
    wire new_Jinkela_wire_6873;
    wire new_Jinkela_wire_3132;
    wire new_Jinkela_wire_1638;
    wire new_Jinkela_wire_6397;
    wire new_Jinkela_wire_2171;
    wire new_Jinkela_wire_2225;
    wire new_Jinkela_wire_7653;
    wire new_Jinkela_wire_9105;
    wire new_Jinkela_wire_6611;
    wire new_Jinkela_wire_5348;
    wire new_Jinkela_wire_2875;
    wire new_Jinkela_wire_9705;
    wire new_Jinkela_wire_3291;
    wire new_Jinkela_wire_7907;
    wire new_Jinkela_wire_6486;
    wire n_0444_;
    wire new_Jinkela_wire_5896;
    wire new_net_2509;
    wire n_1265_;
    wire new_Jinkela_wire_4399;
    wire new_Jinkela_wire_10079;
    wire n_0120_;
    wire new_Jinkela_wire_1856;
    wire new_Jinkela_wire_368;
    wire new_Jinkela_wire_100;
    wire n_0540_;
    wire new_Jinkela_wire_6150;
    wire new_Jinkela_wire_4953;
    wire new_Jinkela_wire_7413;
    wire new_Jinkela_wire_2629;
    wire new_Jinkela_wire_1890;
    wire new_Jinkela_wire_10390;
    wire new_Jinkela_wire_6149;
    wire new_Jinkela_wire_6775;
    wire new_Jinkela_wire_2072;
    wire new_Jinkela_wire_8384;
    wire new_Jinkela_wire_2646;
    wire new_Jinkela_wire_567;
    wire new_Jinkela_wire_6815;
    wire new_Jinkela_wire_6999;
    wire new_Jinkela_wire_3228;
    wire new_Jinkela_wire_739;
    wire new_Jinkela_wire_5399;
    wire new_Jinkela_wire_1996;
    wire new_Jinkela_wire_5672;
    wire new_Jinkela_wire_5152;
    wire new_Jinkela_wire_2632;
    wire new_Jinkela_wire_4570;
    wire n_1237_;
    wire new_Jinkela_wire_2816;
    wire new_Jinkela_wire_8046;
    wire new_Jinkela_wire_2151;
    wire new_Jinkela_wire_8241;
    wire new_Jinkela_wire_6154;
    wire n_1025_;
    wire new_Jinkela_wire_2326;
    wire n_0059_;
    wire n_0705_;
    wire new_Jinkela_wire_5155;
    wire new_Jinkela_wire_5094;
    wire new_Jinkela_wire_8779;
    wire new_Jinkela_wire_5811;
    wire new_Jinkela_wire_5248;
    wire new_Jinkela_wire_6925;
    wire new_Jinkela_wire_1734;
    wire new_Jinkela_wire_9588;
    wire new_Jinkela_wire_7452;
    wire new_Jinkela_wire_2989;
    wire new_Jinkela_wire_5449;
    wire new_Jinkela_wire_8078;
    wire new_Jinkela_wire_7521;
    wire new_Jinkela_wire_3484;
    wire new_Jinkela_wire_7022;
    wire n_0598_;
    wire new_Jinkela_wire_3577;
    wire n_0006_;
    wire new_Jinkela_wire_2932;
    wire new_Jinkela_wire_2415;
    wire new_Jinkela_wire_1724;
    wire new_Jinkela_wire_5424;
    wire new_Jinkela_wire_5540;
    wire n_1353_;
    wire n_0483_;
    wire new_Jinkela_wire_4065;
    wire new_Jinkela_wire_5962;
    wire new_Jinkela_wire_9730;
    wire new_Jinkela_wire_1059;
    wire new_Jinkela_wire_4524;
    wire n_0196_;
    wire new_Jinkela_wire_5051;
    wire new_Jinkela_wire_7895;
    wire new_Jinkela_wire_4438;
    wire new_Jinkela_wire_8130;
    wire new_Jinkela_wire_6446;
    wire new_Jinkela_wire_6338;
    wire new_Jinkela_wire_1036;
    wire n_0448_;
    wire new_Jinkela_wire_2346;
    wire new_Jinkela_wire_4319;
    wire new_Jinkela_wire_5578;
    wire n_0035_;
    wire new_Jinkela_wire_10607;
    wire new_Jinkela_wire_6055;
    wire new_Jinkela_wire_356;
    wire n_0236_;
    wire new_Jinkela_wire_6123;
    wire n_0376_;
    wire new_Jinkela_wire_3631;
    wire new_Jinkela_wire_6922;
    wire new_Jinkela_wire_3882;
    wire new_Jinkela_wire_9838;
    wire new_Jinkela_wire_5326;
    wire new_Jinkela_wire_7534;
    wire new_Jinkela_wire_7031;
    wire new_Jinkela_wire_4916;
    wire new_Jinkela_wire_2089;
    wire new_Jinkela_wire_462;
    wire new_Jinkela_wire_1825;
    wire new_Jinkela_wire_4836;
    wire new_Jinkela_wire_9580;
    wire new_Jinkela_wire_2464;
    wire new_Jinkela_wire_9442;
    wire new_Jinkela_wire_1325;
    wire new_Jinkela_wire_8984;
    wire new_Jinkela_wire_5717;
    wire n_0873_;
    wire new_Jinkela_wire_895;
    wire new_Jinkela_wire_8242;
    wire n_0845_;
    wire new_Jinkela_wire_3112;
    wire new_Jinkela_wire_2933;
    wire n_0314_;
    wire new_Jinkela_wire_10157;
    wire new_Jinkela_wire_1266;
    wire new_Jinkela_wire_1849;
    wire new_Jinkela_wire_3793;
    wire new_Jinkela_wire_3517;
    wire new_Jinkela_wire_631;
    wire n_0958_;
    wire new_Jinkela_wire_9808;
    wire new_Jinkela_wire_4440;
    wire new_Jinkela_wire_6326;
    wire new_Jinkela_wire_10556;
    wire n_0638_;
    wire new_Jinkela_wire_3667;
    wire new_Jinkela_wire_5694;
    wire n_1115_;
    wire new_Jinkela_wire_10408;
    wire new_Jinkela_wire_7374;
    wire new_Jinkela_wire_9167;
    wire new_Jinkela_wire_6232;
    wire new_Jinkela_wire_2534;
    wire new_Jinkela_wire_8280;
    wire new_Jinkela_wire_6139;
    wire n_1121_;
    wire new_Jinkela_wire_3466;
    wire new_Jinkela_wire_4021;
    wire new_Jinkela_wire_5026;
    wire new_Jinkela_wire_9317;
    wire new_Jinkela_wire_2893;
    wire new_Jinkela_wire_7074;
    wire n_0575_;
    wire new_Jinkela_wire_6716;
    wire n_1282_;
    wire new_Jinkela_wire_6417;
    wire new_Jinkela_wire_3418;
    wire new_Jinkela_wire_1920;
    wire new_Jinkela_wire_7590;
    wire new_Jinkela_wire_4071;
    wire new_Jinkela_wire_4025;
    wire new_Jinkela_wire_1295;
    wire new_Jinkela_wire_2772;
    wire new_Jinkela_wire_2192;
    wire new_Jinkela_wire_8161;
    wire new_Jinkela_wire_6344;
    wire new_Jinkela_wire_8593;
    wire new_Jinkela_wire_8851;
    wire new_Jinkela_wire_5517;
    wire new_Jinkela_wire_1803;
    wire new_Jinkela_wire_10163;
    wire new_Jinkela_wire_8612;
    wire new_net_5;
    wire n_1330_;
    wire new_Jinkela_wire_958;
    wire new_Jinkela_wire_6679;
    wire new_Jinkela_wire_2862;
    wire new_Jinkela_wire_10371;
    wire new_Jinkela_wire_4702;
    wire n_1086_;
    wire new_Jinkela_wire_3423;
    wire new_Jinkela_wire_9614;
    wire new_Jinkela_wire_398;
    wire new_Jinkela_wire_10117;
    wire new_Jinkela_wire_8413;
    wire new_Jinkela_wire_4093;
    wire new_Jinkela_wire_10360;
    wire new_Jinkela_wire_6856;
    wire new_Jinkela_wire_6253;
    wire new_Jinkela_wire_10515;
    wire new_Jinkela_wire_126;
    wire new_Jinkela_wire_6148;
    wire new_Jinkela_wire_5469;
    wire new_Jinkela_wire_947;
    wire new_Jinkela_wire_9517;
    wire n_0447_;
    wire new_Jinkela_wire_901;
    wire new_Jinkela_wire_5216;
    wire new_Jinkela_wire_9907;
    wire new_Jinkela_wire_1084;
    wire new_Jinkela_wire_1390;
    wire new_Jinkela_wire_1024;
    wire n_0504_;
    wire new_Jinkela_wire_217;
    wire new_Jinkela_wire_8363;
    wire new_Jinkela_wire_9530;
    wire new_Jinkela_wire_8501;
    wire new_Jinkela_wire_433;
    wire new_Jinkela_wire_24;
    wire new_Jinkela_wire_943;
    wire new_Jinkela_wire_4637;
    wire n_1307_;
    wire new_Jinkela_wire_3242;
    wire new_Jinkela_wire_2650;
    wire new_Jinkela_wire_10161;
    wire new_Jinkela_wire_723;
    wire new_Jinkela_wire_1495;
    wire new_Jinkela_wire_4165;
    wire new_Jinkela_wire_5251;
    wire new_Jinkela_wire_172;
    wire new_Jinkela_wire_9928;
    wire new_Jinkela_wire_3146;
    wire new_Jinkela_wire_5040;
    wire new_Jinkela_wire_5194;
    wire new_Jinkela_wire_6840;
    wire new_Jinkela_wire_9158;
    wire new_Jinkela_wire_5278;
    wire new_Jinkela_wire_9114;
    wire new_Jinkela_wire_8812;
    wire new_Jinkela_wire_9585;
    wire n_0210_;
    wire new_Jinkela_wire_7899;
    wire new_Jinkela_wire_7396;
    wire new_Jinkela_wire_4262;
    wire new_Jinkela_wire_3344;
    wire new_Jinkela_wire_5138;
    wire n_1347_;
    wire new_Jinkela_wire_5780;
    wire new_Jinkela_wire_9350;
    wire new_Jinkela_wire_9367;
    wire new_Jinkela_wire_6713;
    wire new_Jinkela_wire_4097;
    wire new_Jinkela_wire_7474;
    wire n_1296_;
    wire new_Jinkela_wire_6538;
    wire new_Jinkela_wire_4510;
    wire n_1293_;
    wire new_Jinkela_wire_4104;
    wire new_Jinkela_wire_1721;
    wire new_Jinkela_wire_5360;
    wire new_Jinkela_wire_9611;
    wire new_Jinkela_wire_3774;
    wire new_Jinkela_wire_10613;
    wire new_Jinkela_wire_10008;
    wire new_Jinkela_wire_1771;
    wire new_Jinkela_wire_9118;
    wire new_Jinkela_wire_6862;
    wire new_Jinkela_wire_5412;
    wire new_Jinkela_wire_6365;
    wire new_Jinkela_wire_7719;
    wire new_Jinkela_wire_10114;
    wire new_Jinkela_wire_3359;
    wire new_Jinkela_wire_670;
    wire new_Jinkela_wire_10345;
    wire new_Jinkela_wire_706;
    wire new_Jinkela_wire_7543;
    wire n_0243_;
    wire new_Jinkela_wire_5121;
    wire new_Jinkela_wire_9491;
    wire new_Jinkela_wire_4084;
    wire new_Jinkela_wire_9720;
    wire new_Jinkela_wire_6302;
    wire new_Jinkela_wire_5142;
    wire n_1309_;
    wire new_Jinkela_wire_2692;
    wire new_Jinkela_wire_2164;
    wire new_Jinkela_wire_3753;
    wire new_Jinkela_wire_8466;
    wire new_Jinkela_wire_5741;
    wire new_Jinkela_wire_3382;
    wire new_Jinkela_wire_5965;
    wire new_Jinkela_wire_983;
    wire new_Jinkela_wire_379;
    wire new_Jinkela_wire_6643;
    wire new_Jinkela_wire_397;
    wire new_Jinkela_wire_1824;
    wire new_Jinkela_wire_8412;
    wire new_Jinkela_wire_7499;
    wire new_Jinkela_wire_7329;
    wire n_0263_;
    wire new_Jinkela_wire_3803;
    wire new_Jinkela_wire_2071;
    wire new_Jinkela_wire_7827;
    wire n_1072_;
    wire new_Jinkela_wire_5904;
    wire new_Jinkela_wire_10274;
    wire n_0880_;
    wire new_Jinkela_wire_393;
    wire new_Jinkela_wire_9617;
    wire new_Jinkela_wire_1496;
    wire new_Jinkela_wire_9036;
    wire new_Jinkela_wire_1307;
    wire new_net_2523;
    wire new_Jinkela_wire_7182;
    wire new_Jinkela_wire_3597;
    wire new_Jinkela_wire_1195;
    wire new_Jinkela_wire_10378;
    wire new_Jinkela_wire_8278;
    wire new_Jinkela_wire_10212;
    wire new_Jinkela_wire_2802;
    wire n_1050_;
    wire new_Jinkela_wire_556;
    wire new_Jinkela_wire_10342;
    wire new_Jinkela_wire_7519;
    wire new_Jinkela_wire_10386;
    wire new_Jinkela_wire_1356;
    wire new_Jinkela_wire_5990;
    wire new_Jinkela_wire_452;
    wire n_0618_;
    wire new_Jinkela_wire_5352;
    wire new_Jinkela_wire_9713;
    wire new_Jinkela_wire_9661;
    wire new_Jinkela_wire_2010;
    wire new_Jinkela_wire_3177;
    wire new_Jinkela_wire_8010;
    wire n_1069_;
    wire new_Jinkela_wire_3494;
    wire new_Jinkela_wire_2182;
    wire new_Jinkela_wire_3167;
    wire new_Jinkela_wire_7095;
    wire new_Jinkela_wire_2174;
    wire new_Jinkela_wire_8816;
    wire new_Jinkela_wire_8279;
    wire new_Jinkela_wire_7979;
    wire new_Jinkela_wire_6991;
    wire new_Jinkela_wire_9074;
    wire new_Jinkela_wire_4305;
    wire new_Jinkela_wire_5797;
    wire new_Jinkela_wire_5836;
    wire new_Jinkela_wire_5537;
    wire new_Jinkela_wire_5846;
    wire new_Jinkela_wire_9911;
    wire new_Jinkela_wire_7399;
    wire new_Jinkela_wire_2949;
    wire new_Jinkela_wire_3738;
    wire new_Jinkela_wire_427;
    wire new_Jinkela_wire_5408;
    wire n_0879_;
    wire new_Jinkela_wire_6249;
    wire new_Jinkela_wire_3756;
    wire new_Jinkela_wire_9939;
    wire new_Jinkela_wire_2162;
    wire new_Jinkela_wire_4956;
    wire new_Jinkela_wire_6421;
    wire new_Jinkela_wire_6271;
    wire new_Jinkela_wire_3788;
    wire new_Jinkela_wire_2455;
    wire new_Jinkela_wire_7302;
    wire n_0192_;
    wire n_0968_;
    wire new_Jinkela_wire_949;
    wire new_Jinkela_wire_9115;
    wire new_Jinkela_wire_6437;
    wire new_Jinkela_wire_915;
    wire new_Jinkela_wire_9297;
    wire n_0358_;
    wire new_Jinkela_wire_7841;
    wire new_Jinkela_wire_10364;
    wire n_0685_;
    wire new_Jinkela_wire_10403;
    wire new_Jinkela_wire_8373;
    wire n_0284_;
    wire new_Jinkela_wire_9081;
    wire new_Jinkela_wire_454;
    wire new_Jinkela_wire_8037;
    wire new_Jinkela_wire_4494;
    wire new_Jinkela_wire_4941;
    wire new_Jinkela_wire_2203;
    wire new_Jinkela_wire_976;
    wire n_0428_;
    wire new_Jinkela_wire_4064;
    wire new_Jinkela_wire_1867;
    wire n_0562_;
    wire new_Jinkela_wire_9233;
    wire new_Jinkela_wire_10047;
    wire new_Jinkela_wire_5618;
    wire new_Jinkela_wire_4602;
    wire new_Jinkela_wire_1914;
    wire new_Jinkela_wire_2258;
    wire new_Jinkela_wire_8588;
    wire new_Jinkela_wire_4701;
    wire new_Jinkela_wire_2514;
    wire new_Jinkela_wire_8890;
    wire new_Jinkela_wire_1249;
    wire new_Jinkela_wire_7295;
    wire new_Jinkela_wire_3526;
    wire new_Jinkela_wire_1468;
    wire new_Jinkela_wire_1371;
    wire new_Jinkela_wire_6133;
    wire new_Jinkela_wire_3904;
    wire new_Jinkela_wire_1702;
    wire new_Jinkela_wire_4236;
    wire new_Jinkela_wire_6329;
    wire new_Jinkela_wire_1838;
    wire new_Jinkela_wire_4142;
    wire new_Jinkela_wire_10606;
    wire new_Jinkela_wire_5928;
    wire new_Jinkela_wire_7660;
    wire new_Jinkela_wire_2602;
    wire new_Jinkela_wire_7800;
    wire new_Jinkela_wire_5160;
    wire new_Jinkela_wire_7862;
    wire new_Jinkela_wire_5593;
    wire new_Jinkela_wire_2664;
    wire new_Jinkela_wire_469;
    wire new_Jinkela_wire_9148;
    wire new_Jinkela_wire_1549;
    wire n_0991_;
    wire new_Jinkela_wire_6312;
    wire new_Jinkela_wire_4559;
    wire n_1325_;
    wire n_0197_;
    wire new_Jinkela_wire_2956;
    wire new_Jinkela_wire_2349;
    wire new_Jinkela_wire_2704;
    wire new_Jinkela_wire_9327;
    wire new_Jinkela_wire_985;
    wire new_Jinkela_wire_2381;
    wire new_Jinkela_wire_1463;
    wire new_Jinkela_wire_316;
    wire new_Jinkela_wire_3214;
    wire new_Jinkela_wire_1035;
    wire new_Jinkela_wire_10523;
    wire new_Jinkela_wire_5876;
    wire new_Jinkela_wire_6544;
    wire new_Jinkela_wire_8496;
    wire new_Jinkela_wire_8366;
    wire new_Jinkela_wire_1212;
    wire new_Jinkela_wire_624;
    wire new_Jinkela_wire_9494;
    wire new_Jinkela_wire_10624;
    wire new_Jinkela_wire_8644;
    wire n_0909_;
    wire new_Jinkela_wire_5807;
    wire new_Jinkela_wire_8688;
    wire new_Jinkela_wire_9779;
    wire new_Jinkela_wire_853;
    wire new_Jinkela_wire_2977;
    wire new_Jinkela_wire_3357;
    wire n_0026_;
    wire n_0481_;
    wire new_Jinkela_wire_2364;
    wire new_Jinkela_wire_932;
    wire new_Jinkela_wire_7241;
    wire new_Jinkela_wire_7555;
    wire new_Jinkela_wire_9111;
    wire new_Jinkela_wire_3506;
    wire new_Jinkela_wire_484;
    wire n_0686_;
    wire n_0801_;
    wire new_Jinkela_wire_874;
    wire n_0846_;
    wire new_Jinkela_wire_9056;
    wire new_Jinkela_wire_8;
    wire new_Jinkela_wire_1965;
    wire new_Jinkela_wire_9141;
    wire new_Jinkela_wire_5832;
    wire new_Jinkela_wire_9922;
    wire n_0894_;
    wire new_Jinkela_wire_9673;
    wire new_Jinkela_wire_4409;
    wire new_Jinkela_wire_5321;
    wire new_Jinkela_wire_5526;
    wire new_Jinkela_wire_245;
    wire new_Jinkela_wire_147;
    wire new_Jinkela_wire_10277;
    wire new_Jinkela_wire_8115;
    wire new_Jinkela_wire_8507;
    wire new_Jinkela_wire_5193;
    wire new_Jinkela_wire_444;
    wire n_1057_;
    wire n_0384_;
    wire new_Jinkela_wire_4385;
    wire new_Jinkela_wire_7029;
    wire new_Jinkela_wire_1339;
    wire new_Jinkela_wire_4447;
    wire new_Jinkela_wire_839;
    wire new_Jinkela_wire_3668;
    wire new_Jinkela_wire_8394;
    wire new_Jinkela_wire_2595;
    wire new_Jinkela_wire_8226;
    wire new_Jinkela_wire_6259;
    wire new_Jinkela_wire_8769;
    wire new_Jinkela_wire_5842;
    wire new_Jinkela_wire_6808;
    wire new_Jinkela_wire_5344;
    wire n_0919_;
    wire n_1245_;
    wire new_Jinkela_wire_9960;
    wire new_Jinkela_wire_858;
    wire new_Jinkela_wire_8316;
    wire new_Jinkela_wire_824;
    wire new_Jinkela_wire_10491;
    wire new_Jinkela_wire_8019;
    wire n_0068_;
    wire new_Jinkela_wire_8419;
    wire new_Jinkela_wire_3575;
    wire new_Jinkela_wire_5072;
    wire new_Jinkela_wire_6225;
    wire new_Jinkela_wire_8523;
    wire new_Jinkela_wire_8561;
    wire new_Jinkela_wire_2806;
    wire new_Jinkela_wire_6711;
    wire new_Jinkela_wire_5686;
    wire new_Jinkela_wire_3432;
    wire new_Jinkela_wire_9852;
    wire new_Jinkela_wire_4804;
    wire new_Jinkela_wire_10192;
    wire new_Jinkela_wire_3951;
    wire n_0353_;
    wire new_Jinkela_wire_2903;
    wire n_0997_;
    wire new_Jinkela_wire_6041;
    wire new_Jinkela_wire_4128;
    wire new_Jinkela_wire_1019;
    wire new_Jinkela_wire_1273;
    wire new_Jinkela_wire_2043;
    wire new_Jinkela_wire_9455;
    wire new_Jinkela_wire_7576;
    wire new_Jinkela_wire_8540;
    wire new_Jinkela_wire_432;
    wire new_Jinkela_wire_8558;
    wire new_Jinkela_wire_5798;
    wire new_Jinkela_wire_5680;
    wire new_Jinkela_wire_6936;
    wire n_0287_;
    wire new_Jinkela_wire_577;
    wire new_Jinkela_wire_10349;
    wire new_Jinkela_wire_8124;
    wire new_Jinkela_wire_9408;
    wire new_Jinkela_wire_10488;
    wire new_Jinkela_wire_3849;
    wire new_Jinkela_wire_7403;
    wire n_1171_;
    wire new_Jinkela_wire_7136;
    wire new_Jinkela_wire_4086;
    wire new_Jinkela_wire_5263;
    wire n_0087_;
    wire new_Jinkela_wire_2473;
    wire n_1349_;
    wire new_Jinkela_wire_6940;
    wire new_Jinkela_wire_1097;
    wire new_Jinkela_wire_9905;
    wire new_Jinkela_wire_9636;
    wire new_Jinkela_wire_8308;
    wire new_Jinkela_wire_2935;
    wire new_Jinkela_wire_9418;
    wire new_Jinkela_wire_1008;
    wire new_Jinkela_wire_8736;
    wire n_0597_;
    wire new_Jinkela_wire_9904;
    wire new_Jinkela_wire_1862;
    wire n_0214_;
    wire new_Jinkela_wire_752;
    wire new_Jinkela_wire_1198;
    wire new_Jinkela_wire_8567;
    wire new_Jinkela_wire_8654;
    wire n_1126_;
    wire new_Jinkela_wire_9238;
    wire new_Jinkela_wire_6124;
    wire n_1292_;
    wire new_Jinkela_wire_7208;
    wire n_0302_;
    wire new_Jinkela_wire_1380;
    wire n_0529_;
    wire new_Jinkela_wire_2699;
    wire n_1129_;
    wire new_Jinkela_wire_7910;
    wire new_Jinkela_wire_3027;
    wire new_Jinkela_wire_7504;
    wire n_0148_;
    wire new_Jinkela_wire_6062;
    wire new_Jinkela_wire_9226;
    wire new_Jinkela_wire_7273;
    wire n_1239_;
    wire new_Jinkela_wire_2342;
    wire new_Jinkela_wire_2421;
    wire new_Jinkela_wire_3009;
    wire new_Jinkela_wire_2105;
    wire new_Jinkela_wire_1340;
    wire new_Jinkela_wire_7607;
    wire new_Jinkela_wire_5468;
    wire new_Jinkela_wire_3690;
    wire new_Jinkela_wire_10442;
    wire new_Jinkela_wire_2524;
    wire n_0388_;
    wire new_Jinkela_wire_205;
    wire new_Jinkela_wire_4073;
    wire new_Jinkela_wire_6756;
    wire new_Jinkela_wire_4094;
    wire new_Jinkela_wire_5030;
    wire new_Jinkela_wire_4731;
    wire new_Jinkela_wire_3757;
    wire n_0751_;
    wire new_Jinkela_wire_6386;
    wire new_Jinkela_wire_4712;
    wire n_1161_;
    wire new_Jinkela_wire_9198;
    wire new_Jinkela_wire_2280;
    wire new_Jinkela_wire_999;
    wire new_Jinkela_wire_4608;
    wire new_Jinkela_wire_3529;
    wire new_Jinkela_wire_6093;
    wire new_Jinkela_wire_2596;
    wire new_Jinkela_wire_2673;
    wire new_Jinkela_wire_6933;
    wire new_Jinkela_wire_384;
    wire new_Jinkela_wire_7350;
    wire new_Jinkela_wire_8178;
    wire new_Jinkela_wire_9432;
    wire n_1305_;
    wire new_Jinkela_wire_680;
    wire new_Jinkela_wire_9793;
    wire new_Jinkela_wire_7008;
    wire new_Jinkela_wire_5773;
    wire new_Jinkela_wire_2774;
    wire new_Jinkela_wire_2523;
    wire new_Jinkela_wire_7228;
    wire new_Jinkela_wire_9138;
    wire new_Jinkela_wire_2654;
    wire new_Jinkela_wire_5187;
    wire new_Jinkela_wire_2129;
    wire new_Jinkela_wire_6588;
    wire new_Jinkela_wire_9877;
    wire new_Jinkela_wire_5309;
    wire new_Jinkela_wire_4439;
    wire n_1232_;
    wire new_Jinkela_wire_3841;
    wire new_Jinkela_wire_1787;
    wire new_Jinkela_wire_8499;
    wire new_Jinkela_wire_1845;
    wire new_Jinkela_wire_2562;
    wire new_Jinkela_wire_6398;
    wire new_Jinkela_wire_2462;
    wire new_Jinkela_wire_7864;
    wire new_Jinkela_wire_115;
    wire new_Jinkela_wire_10144;
    wire new_Jinkela_wire_6050;
    wire new_Jinkela_wire_4838;
    wire new_Jinkela_wire_3075;
    wire new_Jinkela_wire_6498;
    wire new_Jinkela_wire_2312;
    wire new_Jinkela_wire_359;
    wire n_0994_;
    wire new_Jinkela_wire_7454;
    wire new_Jinkela_wire_6842;
    wire new_Jinkela_wire_8310;
    wire new_Jinkela_wire_9755;
    wire new_Jinkela_wire_5387;
    wire new_Jinkela_wire_5936;
    wire new_Jinkela_wire_6642;
    wire new_Jinkela_wire_8837;
    wire new_Jinkela_wire_5447;
    wire n_0564_;
    wire new_Jinkela_wire_2436;
    wire new_Jinkela_wire_8884;
    wire new_Jinkela_wire_4204;
    wire new_Jinkela_wire_9295;
    wire new_Jinkela_wire_2789;
    wire new_Jinkela_wire_9463;
    wire new_Jinkela_wire_1515;
    wire new_Jinkela_wire_9339;
    wire new_Jinkela_wire_6092;
    wire new_Jinkela_wire_4543;
    wire new_Jinkela_wire_9602;
    wire new_Jinkela_wire_99;
    wire new_Jinkela_wire_2874;
    wire new_Jinkela_wire_8698;
    wire new_Jinkela_wire_4365;
    wire new_Jinkela_wire_2592;
    wire new_Jinkela_wire_1063;
    wire n_1146_;
    wire new_Jinkela_wire_5055;
    wire new_Jinkela_wire_4122;
    wire new_Jinkela_wire_312;
    wire new_Jinkela_wire_7758;
    wire n_1037_;
    wire new_Jinkela_wire_4079;
    wire new_Jinkela_wire_9323;
    wire new_Jinkela_wire_528;
    wire new_Jinkela_wire_4432;
    wire new_Jinkela_wire_518;
    wire new_Jinkela_wire_2791;
    wire n_0917_;
    wire new_Jinkela_wire_2653;
    wire n_0585_;
    wire new_Jinkela_wire_1527;
    wire new_Jinkela_wire_7106;
    wire new_Jinkela_wire_8408;
    wire new_Jinkela_wire_9600;
    wire new_Jinkela_wire_5592;
    wire new_Jinkela_wire_9322;
    wire new_Jinkela_wire_10603;
    wire new_Jinkela_wire_467;
    wire new_Jinkela_wire_6905;
    wire new_Jinkela_wire_1159;
    wire new_Jinkela_wire_10295;
    wire new_Jinkela_wire_5255;
    wire new_Jinkela_wire_6607;
    wire new_Jinkela_wire_9897;
    wire new_Jinkela_wire_4657;
    wire new_Jinkela_wire_401;
    wire n_1268_;
    wire new_Jinkela_wire_5759;
    wire new_Jinkela_wire_65;
    wire new_Jinkela_wire_8687;
    wire new_Jinkela_wire_7662;
    wire new_Jinkela_wire_6183;
    wire new_Jinkela_wire_4617;
    wire new_Jinkela_wire_9353;
    wire new_Jinkela_wire_8551;
    wire new_Jinkela_wire_9311;
    wire new_Jinkela_wire_8108;
    wire new_Jinkela_wire_1528;
    wire new_Jinkela_wire_5125;
    wire new_Jinkela_wire_104;
    wire new_Jinkela_wire_6575;
    wire new_Jinkela_wire_6449;
    wire new_Jinkela_wire_5561;
    wire new_Jinkela_wire_8570;
    wire new_Jinkela_wire_8085;
    wire new_Jinkela_wire_5252;
    wire new_Jinkela_wire_594;
    wire new_Jinkela_wire_4103;
    wire new_Jinkela_wire_3861;
    wire new_Jinkela_wire_3021;
    wire new_Jinkela_wire_10367;
    wire n_0557_;
    wire n_1080_;
    wire new_Jinkela_wire_7048;
    wire new_Jinkela_wire_2122;
    wire new_Jinkela_wire_89;
    wire new_Jinkela_wire_2329;
    wire new_Jinkela_wire_3829;
    wire new_Jinkela_wire_9265;
    wire new_Jinkela_wire_3846;
    wire new_Jinkela_wire_8483;
    wire new_Jinkela_wire_5751;
    wire new_Jinkela_wire_1292;
    wire new_Jinkela_wire_3898;
    wire new_Jinkela_wire_4018;
    wire n_0579_;
    wire new_Jinkela_wire_707;
    wire new_Jinkela_wire_9520;
    wire new_Jinkela_wire_8045;
    wire new_Jinkela_wire_6286;
    wire new_Jinkela_wire_9437;
    wire new_Jinkela_wire_2272;
    wire new_Jinkela_wire_8284;
    wire new_Jinkela_wire_4074;
    wire new_Jinkela_wire_4770;
    wire new_Jinkela_wire_764;
    wire new_Jinkela_wire_8177;
    wire new_Jinkela_wire_5481;
    wire new_Jinkela_wire_2701;
    wire new_Jinkela_wire_8209;
    wire new_Jinkela_wire_9398;
    wire new_Jinkela_wire_6742;
    wire new_Jinkela_wire_7876;
    wire new_Jinkela_wire_184;
    wire new_Jinkela_wire_6641;
    wire new_Jinkela_wire_5696;
    wire new_Jinkela_wire_6541;
    wire new_Jinkela_wire_1346;
    wire new_Jinkela_wire_8613;
    wire new_Jinkela_wire_2481;
    wire new_Jinkela_wire_8746;
    wire new_Jinkela_wire_7002;
    wire new_Jinkela_wire_2912;
    wire new_Jinkela_wire_2936;
    wire new_Jinkela_wire_2094;
    wire new_Jinkela_wire_2283;
    wire new_Jinkela_wire_4421;
    wire new_Jinkela_wire_4061;
    wire new_Jinkela_wire_1972;
    wire new_Jinkela_wire_708;
    wire new_Jinkela_wire_6950;
    wire new_Jinkela_wire_2193;
    wire new_Jinkela_wire_8997;
    wire new_net_2543;
    wire n_0297_;
    wire new_Jinkela_wire_10320;
    wire new_Jinkela_wire_8376;
    wire n_0410_;
    wire n_0144_;
    wire new_Jinkela_wire_8088;
    wire new_Jinkela_wire_4157;
    wire new_Jinkela_wire_5623;
    wire new_Jinkela_wire_9917;
    wire new_Jinkela_wire_5008;
    wire n_0640_;
    wire new_Jinkela_wire_5576;
    wire new_Jinkela_wire_4444;
    wire new_Jinkela_wire_9080;
    wire new_Jinkela_wire_4349;
    wire new_Jinkela_wire_8063;
    wire new_Jinkela_wire_5461;
    wire new_Jinkela_wire_170;
    wire new_Jinkela_wire_8843;
    wire new_Jinkela_wire_3554;
    wire n_0531_;
    wire new_Jinkela_wire_5613;
    wire new_Jinkela_wire_584;
    wire new_Jinkela_wire_3137;
    wire new_Jinkela_wire_6520;
    wire new_Jinkela_wire_5516;
    wire new_Jinkela_wire_9370;
    wire new_Jinkela_wire_4908;
    wire new_Jinkela_wire_6046;
    wire new_Jinkela_wire_2794;
    wire new_Jinkela_wire_7248;
    wire new_Jinkela_wire_6203;
    wire new_Jinkela_wire_8979;
    wire new_Jinkela_wire_7861;
    wire new_Jinkela_wire_10482;
    wire new_Jinkela_wire_9570;
    wire new_Jinkela_wire_2350;
    wire new_Jinkela_wire_248;
    wire new_Jinkela_wire_3138;
    wire new_Jinkela_wire_1351;
    wire new_Jinkela_wire_1282;
    wire new_Jinkela_wire_2488;
    wire new_Jinkela_wire_992;
    wire new_Jinkela_wire_6211;
    wire new_Jinkela_wire_9592;
    wire new_Jinkela_wire_472;
    wire new_Jinkela_wire_6850;
    wire new_Jinkela_wire_5241;
    wire new_Jinkela_wire_866;
    wire new_Jinkela_wire_791;
    wire new_Jinkela_wire_1588;
    wire new_Jinkela_wire_3341;
    wire n_0572_;
    wire new_Jinkela_wire_284;
    wire new_Jinkela_wire_2039;
    wire new_Jinkela_wire_9137;
    wire n_0981_;
    wire new_Jinkela_wire_7971;
    wire new_Jinkela_wire_9278;
    wire new_Jinkela_wire_4800;
    wire new_Jinkela_wire_5113;
    wire new_Jinkela_wire_944;
    wire new_Jinkela_wire_9001;
    wire new_Jinkela_wire_3763;
    wire new_Jinkela_wire_6463;
    wire new_Jinkela_wire_7940;
    wire new_Jinkela_wire_6690;
    wire new_Jinkela_wire_7823;
    wire new_Jinkela_wire_10083;
    wire new_Jinkela_wire_6631;
    wire new_Jinkela_wire_7771;
    wire n_1035_;
    wire new_Jinkela_wire_9650;
    wire n_0794_;
    wire new_Jinkela_wire_9583;
    wire new_Jinkela_wire_1102;
    wire new_Jinkela_wire_9754;
    wire new_Jinkela_wire_2240;
    wire new_Jinkela_wire_1557;
    wire new_Jinkela_wire_4926;
    wire new_Jinkela_wire_2184;
    wire new_Jinkela_wire_8716;
    wire new_Jinkela_wire_2696;
    wire new_Jinkela_wire_8621;
    wire new_Jinkela_wire_10057;
    wire new_Jinkela_wire_9924;
    wire new_Jinkela_wire_2665;
    wire new_Jinkela_wire_2046;
    wire new_Jinkela_wire_601;
    wire new_Jinkela_wire_1804;
    wire new_Jinkela_wire_9514;
    wire n_0669_;
    wire new_Jinkela_wire_3787;
    wire new_Jinkela_wire_1858;
    wire new_Jinkela_wire_162;
    wire new_Jinkela_wire_8538;
    wire new_Jinkela_wire_9753;
    wire new_Jinkela_wire_9809;
    wire new_Jinkela_wire_5277;
    wire new_Jinkela_wire_10201;
    wire new_Jinkela_wire_6995;
    wire new_Jinkela_wire_2095;
    wire new_Jinkela_wire_4091;
    wire new_Jinkela_wire_6496;
    wire new_Jinkela_wire_6658;
    wire new_Jinkela_wire_8641;
    wire new_Jinkela_wire_2220;
    wire n_0071_;
    wire n_1063_;
    wire n_0698_;
    wire new_Jinkela_wire_2057;
    wire new_Jinkela_wire_8426;
    wire new_Jinkela_wire_160;
    wire new_Jinkela_wire_8331;
    wire new_Jinkela_wire_8141;
    wire new_Jinkela_wire_7674;
    wire new_Jinkela_wire_6058;
    wire new_Jinkela_wire_1210;
    wire new_Jinkela_wire_3142;
    wire new_Jinkela_wire_6956;
    wire new_Jinkela_wire_6760;
    wire new_Jinkela_wire_143;
    wire new_Jinkela_wire_2913;
    wire n_0419_;
    wire new_Jinkela_wire_4382;
    wire new_Jinkela_wire_6341;
    wire new_Jinkela_wire_8545;
    wire new_Jinkela_wire_675;
    wire new_Jinkela_wire_6517;
    wire new_Jinkela_wire_10361;
    wire n_0127_;
    wire n_1174_;
    wire new_Jinkela_wire_2689;
    wire new_Jinkela_wire_7796;
    wire n_0692_;
    wire new_Jinkela_wire_9214;
    wire new_Jinkela_wire_2641;
    wire new_Jinkela_wire_10560;
    wire new_Jinkela_wire_6801;
    wire new_Jinkela_wire_695;
    wire new_Jinkela_wire_3190;
    wire new_Jinkela_wire_8672;
    wire new_Jinkela_wire_1239;
    wire new_Jinkela_wire_5291;
    wire new_Jinkela_wire_3223;
    wire new_Jinkela_wire_4208;
    wire new_Jinkela_wire_6963;
    wire new_Jinkela_wire_2295;
    wire new_Jinkela_wire_2400;
    wire new_Jinkela_wire_10152;
    wire new_Jinkela_wire_3747;
    wire new_Jinkela_wire_7161;
    wire new_Jinkela_wire_8239;
    wire new_Jinkela_wire_1462;
    wire new_Jinkela_wire_4765;
    wire new_Jinkela_wire_2356;
    wire new_Jinkela_wire_8692;
    wire new_Jinkela_wire_9681;
    wire new_Jinkela_wire_6570;
    wire new_Jinkela_wire_2128;
    wire n_0516_;
    wire new_Jinkela_wire_4270;
    wire new_Jinkela_wire_666;
    wire new_Jinkela_wire_9261;
    wire new_Jinkela_wire_2120;
    wire new_Jinkela_wire_8170;
    wire new_Jinkela_wire_1149;
    wire new_Jinkela_wire_3713;
    wire new_Jinkela_wire_9364;
    wire new_Jinkela_wire_5020;
    wire new_Jinkela_wire_9853;
    wire n_0152_;
    wire new_Jinkela_wire_558;
    wire new_Jinkela_wire_2429;
    wire new_Jinkela_wire_485;
    wire new_Jinkela_wire_918;
    wire new_Jinkela_wire_6054;
    wire new_Jinkela_wire_9682;
    wire n_0499_;
    wire n_1224_;
    wire new_Jinkela_wire_9072;
    wire new_Jinkela_wire_5156;
    wire new_Jinkela_wire_8511;
    wire new_Jinkela_wire_6831;
    wire new_Jinkela_wire_5075;
    wire new_Jinkela_wire_10402;
    wire new_Jinkela_wire_378;
    wire new_Jinkela_wire_7344;
    wire new_Jinkela_wire_3183;
    wire new_Jinkela_wire_9298;
    wire new_Jinkela_wire_8257;
    wire new_Jinkela_wire_9457;
    wire new_Jinkela_wire_7184;
    wire new_Jinkela_wire_2253;
    wire new_Jinkela_wire_10209;
    wire new_Jinkela_wire_6128;
    wire new_Jinkela_wire_10535;
    wire new_Jinkela_wire_5661;
    wire new_Jinkela_wire_9665;
    wire new_Jinkela_wire_5938;
    wire n_0011_;
    wire new_Jinkela_wire_5852;
    wire new_Jinkela_wire_6803;
    wire new_Jinkela_wire_7315;
    wire new_Jinkela_wire_1534;
    wire new_Jinkela_wire_2388;
    wire new_net_2511;
    wire new_Jinkela_wire_7494;
    wire new_Jinkela_wire_1188;
    wire new_Jinkela_wire_10446;
    wire new_Jinkela_wire_8328;
    wire new_Jinkela_wire_3616;
    wire new_Jinkela_wire_8096;
    wire new_Jinkela_wire_4502;
    wire n_0427_;
    wire new_Jinkela_wire_4964;
    wire new_Jinkela_wire_1403;
    wire new_Jinkela_wire_1563;
    wire new_Jinkela_wire_8353;
    wire new_Jinkela_wire_4561;
    wire new_Jinkela_wire_6239;
    wire new_Jinkela_wire_2652;
    wire new_Jinkela_wire_687;
    wire new_Jinkela_wire_7755;
    wire new_Jinkela_wire_3116;
    wire new_Jinkela_wire_5359;
    wire n_0422_;
    wire new_Jinkela_wire_4917;
    wire new_Jinkela_wire_8057;
    wire new_Jinkela_wire_6708;
    wire new_Jinkela_wire_2715;
    wire new_Jinkela_wire_9087;
    wire new_Jinkela_wire_152;
    wire new_Jinkela_wire_10511;
    wire new_Jinkela_wire_9920;
    wire new_Jinkela_wire_5606;
    wire new_Jinkela_wire_579;
    wire new_Jinkela_wire_9065;
    wire new_Jinkela_wire_8609;
    wire n_0254_;
    wire new_Jinkela_wire_5388;
    wire new_Jinkela_wire_3899;
    wire new_Jinkela_wire_1814;
    wire new_Jinkela_wire_6431;
    wire new_Jinkela_wire_5102;
    wire new_Jinkela_wire_309;
    wire new_Jinkela_wire_4630;
    wire new_Jinkela_wire_4459;
    wire new_Jinkela_wire_3300;
    wire new_Jinkela_wire_830;
    wire new_Jinkela_wire_1404;
    wire new_Jinkela_wire_8184;
    wire new_Jinkela_wire_3215;
    wire new_Jinkela_wire_8862;
    wire new_Jinkela_wire_3744;
    wire new_Jinkela_wire_746;
    wire new_Jinkela_wire_8544;
    wire new_Jinkela_wire_948;
    wire new_Jinkela_wire_10323;
    wire new_Jinkela_wire_8756;
    wire new_Jinkela_wire_571;
    wire n_1360_;
    wire new_Jinkela_wire_10443;
    wire n_0842_;
    wire n_0847_;
    wire new_Jinkela_wire_6934;
    wire new_Jinkela_wire_8058;
    wire new_Jinkela_wire_4367;
    wire new_Jinkela_wire_4853;
    wire new_Jinkela_wire_2755;
    wire new_Jinkela_wire_4009;
    wire new_Jinkela_wire_3972;
    wire new_Jinkela_wire_2951;
    wire new_Jinkela_wire_7584;
    wire new_Jinkela_wire_9692;
    wire new_Jinkela_wire_8891;
    wire new_Jinkela_wire_10129;
    wire new_Jinkela_wire_8882;
    wire new_Jinkela_wire_6223;
    wire new_Jinkela_wire_8351;
    wire new_Jinkela_wire_5097;
    wire n_0644_;
    wire new_Jinkela_wire_541;
    wire new_Jinkela_wire_9559;
    wire new_Jinkela_wire_5531;
    wire new_Jinkela_wire_5855;
    wire new_Jinkela_wire_2289;
    wire new_Jinkela_wire_10472;
    wire new_Jinkela_wire_4283;
    wire n_1266_;
    wire new_Jinkela_wire_9292;
    wire new_Jinkela_wire_8103;
    wire new_Jinkela_wire_7286;
    wire new_Jinkela_wire_4130;
    wire new_Jinkela_wire_3329;
    wire new_Jinkela_wire_1318;
    wire new_Jinkela_wire_5754;
    wire n_0414_;
    wire new_Jinkela_wire_1500;
    wire new_Jinkela_wire_7792;
    wire new_Jinkela_wire_208;
    wire new_Jinkela_wire_6406;
    wire new_Jinkela_wire_4839;
    wire new_Jinkela_wire_38;
    wire new_Jinkela_wire_1261;
    wire new_net_2519;
    wire new_Jinkela_wire_8494;
    wire new_Jinkela_wire_5697;
    wire n_1151_;
    wire new_Jinkela_wire_9780;
    wire new_Jinkela_wire_2960;
    wire new_Jinkela_wire_4479;
    wire new_Jinkela_wire_1881;
    wire new_Jinkela_wire_6151;
    wire new_Jinkela_wire_8407;
    wire new_Jinkela_wire_2952;
    wire new_Jinkela_wire_6744;
    wire new_Jinkela_wire_3192;
    wire new_Jinkela_wire_4045;
    wire new_Jinkela_wire_9823;
    wire n_1005_;
    wire n_1231_;
    wire new_Jinkela_wire_9512;
    wire new_Jinkela_wire_7736;
    wire new_Jinkela_wire_665;
    wire new_Jinkela_wire_6306;
    wire new_Jinkela_wire_3416;
    wire new_Jinkela_wire_9643;
    wire n_1241_;
    wire new_Jinkela_wire_3437;
    wire new_Jinkela_wire_2234;
    wire n_0570_;
    wire new_Jinkela_wire_9736;
    wire n_0863_;
    wire new_Jinkela_wire_1904;
    wire n_0804_;
    wire n_0555_;
    wire new_Jinkela_wire_10626;
    wire new_Jinkela_wire_1096;
    wire new_Jinkela_wire_4833;
    wire new_Jinkela_wire_965;
    wire new_Jinkela_wire_3912;
    wire new_Jinkela_wire_10513;
    wire new_Jinkela_wire_4024;
    wire new_Jinkela_wire_750;
    wire n_0683_;
    wire new_Jinkela_wire_10336;
    wire new_Jinkela_wire_7988;
    wire new_Jinkela_wire_10444;
    wire new_Jinkela_wire_10050;
    wire new_Jinkela_wire_8952;
    wire new_Jinkela_wire_7628;
    wire new_Jinkela_wire_9696;
    wire new_Jinkela_wire_1152;
    wire new_Jinkela_wire_3064;
    wire new_Jinkela_wire_3182;
    wire new_Jinkela_wire_2736;
    wire new_Jinkela_wire_7323;
    wire new_Jinkela_wire_2700;
    wire new_Jinkela_wire_435;
    wire new_Jinkela_wire_8525;
    wire new_Jinkela_wire_885;
    wire new_Jinkela_wire_6545;
    wire new_Jinkela_wire_7027;
    wire new_Jinkela_wire_504;
    wire new_Jinkela_wire_9876;
    wire new_Jinkela_wire_7804;
    wire new_Jinkela_wire_5166;
    wire new_Jinkela_wire_7447;
    wire new_Jinkela_wire_3305;
    wire new_Jinkela_wire_4152;
    wire new_Jinkela_wire_1156;
    wire new_Jinkela_wire_3169;
    wire n_1358_;
    wire new_Jinkela_wire_9048;
    wire new_Jinkela_wire_9161;
    wire new_Jinkela_wire_1439;
    wire new_Jinkela_wire_8796;
    wire n_0355_;
    wire new_Jinkela_wire_7642;
    wire new_Jinkela_wire_5988;
    wire new_Jinkela_wire_1105;
    wire new_Jinkela_wire_3741;
    wire new_Jinkela_wire_8929;
    wire new_Jinkela_wire_7430;
    wire n_0559_;
    wire new_Jinkela_wire_3644;
    wire new_Jinkela_wire_6233;
    wire new_Jinkela_wire_8726;
    wire new_Jinkela_wire_4445;
    wire new_Jinkela_wire_6037;
    wire n_0111_;
    wire new_Jinkela_wire_4493;
    wire new_Jinkela_wire_4140;
    wire new_Jinkela_wire_1621;
    wire new_Jinkela_wire_6313;
    wire new_Jinkela_wire_677;
    wire new_Jinkela_wire_1601;
    wire new_Jinkela_wire_10539;
    wire new_Jinkela_wire_8522;
    wire new_Jinkela_wire_280;
    wire new_Jinkela_wire_6841;
    wire new_Jinkela_wire_6052;
    wire new_Jinkela_wire_6610;
    wire new_Jinkela_wire_5954;
    wire new_Jinkela_wire_5430;
    wire new_Jinkela_wire_1580;
    wire new_Jinkela_wire_5191;
    wire new_Jinkela_wire_1147;
    wire new_Jinkela_wire_8101;
    wire new_Jinkela_wire_5786;
    wire new_Jinkela_wire_9401;
    wire new_Jinkela_wire_4143;
    wire new_Jinkela_wire_10605;
    wire new_Jinkela_wire_5061;
    wire new_Jinkela_wire_3508;
    wire new_Jinkela_wire_10522;
    wire new_Jinkela_wire_3349;
    wire new_Jinkela_wire_4732;
    wire new_Jinkela_wire_3758;
    wire new_Jinkela_wire_4518;
    wire new_Jinkela_wire_8526;
    wire new_Jinkela_wire_3927;
    wire new_Jinkela_wire_7150;
    wire new_Jinkela_wire_673;
    wire new_Jinkela_wire_3946;
    wire new_Jinkela_wire_5822;
    wire n_1114_;
    wire new_Jinkela_wire_1023;
    wire new_Jinkela_wire_8748;
    wire new_Jinkela_wire_8944;
    wire new_Jinkela_wire_2729;
    wire new_Jinkela_wire_341;
    wire new_Jinkela_wire_788;
    wire new_Jinkela_wire_6704;
    wire new_Jinkela_wire_2725;
    wire n_0249_;
    wire new_Jinkela_wire_9993;
    wire new_Jinkela_wire_6320;
    wire new_net_2495;
    wire new_Jinkela_wire_4970;
    wire new_Jinkela_wire_10102;
    wire n_1287_;
    wire n_0063_;
    wire new_Jinkela_wire_5201;
    wire n_1288_;
    wire new_Jinkela_wire_8823;
    wire new_Jinkela_wire_5226;
    wire new_Jinkela_wire_2007;
    wire new_Jinkela_wire_4521;
    wire new_Jinkela_wire_10524;
    wire new_Jinkela_wire_10151;
    wire new_Jinkela_wire_825;
    wire n_1370_;
    wire new_Jinkela_wire_4706;
    wire new_Jinkela_wire_1575;
    wire new_Jinkela_wire_9714;
    wire new_Jinkela_wire_8807;
    wire new_Jinkela_wire_2720;
    wire new_Jinkela_wire_1372;
    wire new_Jinkela_wire_2776;
    wire new_Jinkela_wire_4572;
    wire new_Jinkela_wire_1209;
    wire new_Jinkela_wire_6807;
    wire new_Jinkela_wire_1922;
    wire new_Jinkela_wire_2621;
    wire new_Jinkela_wire_5404;
    wire new_Jinkela_wire_8491;
    wire new_Jinkela_wire_10438;
    wire new_Jinkela_wire_48;
    wire new_Jinkela_wire_7376;
    wire n_0614_;
    wire new_Jinkela_wire_4944;
    wire new_Jinkela_wire_890;
    wire new_Jinkela_wire_3270;
    wire new_Jinkela_wire_5186;
    wire new_Jinkela_wire_6797;
    wire new_Jinkela_wire_3022;
    wire n_0765_;
    wire n_0469_;
    wire new_Jinkela_wire_1715;
    wire new_Jinkela_wire_7060;
    wire new_Jinkela_wire_3645;
    wire new_Jinkela_wire_5838;
    wire new_Jinkela_wire_9890;
    wire new_Jinkela_wire_6456;
    wire new_Jinkela_wire_1885;
    wire new_Jinkela_wire_9772;
    wire new_Jinkela_wire_10308;
    wire n_0177_;
    wire new_Jinkela_wire_4720;
    wire new_Jinkela_wire_7648;
    wire new_Jinkela_wire_871;
    wire new_Jinkela_wire_10469;
    wire new_Jinkela_wire_9572;
    wire new_Jinkela_wire_1652;
    wire new_Jinkela_wire_8293;
    wire new_Jinkela_wire_4329;
    wire new_Jinkela_wire_8514;
    wire new_Jinkela_wire_9691;
    wire new_Jinkela_wire_8162;
    wire new_Jinkela_wire_6645;
    wire new_Jinkela_wire_2218;
    wire new_Jinkela_wire_5100;
    wire new_Jinkela_wire_3471;
    wire n_1085_;
    wire new_Jinkela_wire_9219;
    wire new_Jinkela_wire_10593;
    wire new_Jinkela_wire_8791;
    wire n_0482_;
    wire n_0105_;
    wire new_Jinkela_wire_4219;
    wire new_Jinkela_wire_4428;
    wire new_Jinkela_wire_7015;
    wire new_Jinkela_wire_2264;
    wire new_net_9;
    wire new_Jinkela_wire_10171;
    wire new_Jinkela_wire_6020;
    wire new_Jinkela_wire_1363;
    wire new_Jinkela_wire_6438;
    wire new_Jinkela_wire_2710;
    wire new_Jinkela_wire_755;
    wire new_Jinkela_wire_6859;
    wire new_Jinkela_wire_8694;
    wire new_Jinkela_wire_1369;
    wire new_Jinkela_wire_745;
    wire new_Jinkela_wire_3525;
    wire new_Jinkela_wire_966;
    wire new_Jinkela_wire_6653;
    wire new_Jinkela_wire_5708;
    wire new_Jinkela_wire_4687;
    wire new_Jinkela_wire_8217;
    wire new_Jinkela_wire_2260;
    wire new_Jinkela_wire_6031;
    wire new_Jinkela_wire_8011;
    wire new_Jinkela_wire_2618;
    wire new_Jinkela_wire_9440;
    wire new_Jinkela_wire_1628;
    wire new_Jinkela_wire_3726;
    wire new_Jinkela_wire_9274;
    wire new_Jinkela_wire_4935;
    wire new_Jinkela_wire_6924;
    wire new_Jinkela_wire_2113;
    wire new_Jinkela_wire_1131;
    wire new_Jinkela_wire_4069;
    wire new_Jinkela_wire_8509;
    wire new_Jinkela_wire_2422;
    wire new_Jinkela_wire_1533;
    wire new_Jinkela_wire_6205;
    wire new_Jinkela_wire_2753;
    wire new_Jinkela_wire_10354;
    wire new_Jinkela_wire_3873;
    wire new_Jinkela_wire_6014;
    wire new_Jinkela_wire_950;
    wire new_Jinkela_wire_5638;
    wire new_Jinkela_wire_840;
    wire new_Jinkela_wire_3630;
    wire new_Jinkela_wire_2670;
    wire new_Jinkela_wire_5139;
    wire new_Jinkela_wire_8970;
    wire new_Jinkela_wire_3844;
    wire new_Jinkela_wire_9199;
    wire new_Jinkela_wire_1354;
    wire new_Jinkela_wire_2724;
    wire new_Jinkela_wire_1939;
    wire new_Jinkela_wire_4052;
    wire new_Jinkela_wire_1706;
    wire new_Jinkela_wire_1843;
    wire new_Jinkela_wire_3205;
    wire n_1106_;
    wire new_Jinkela_wire_1746;
    wire n_1094_;
    wire new_Jinkela_wire_2907;
    wire new_Jinkela_wire_5454;
    wire new_Jinkela_wire_6026;
    wire n_0455_;
    wire new_Jinkela_wire_1998;
    wire new_Jinkela_wire_6667;
    wire new_Jinkela_wire_7689;
    wire new_Jinkela_wire_9574;
    wire new_Jinkela_wire_7820;
    wire new_Jinkela_wire_6370;
    wire new_Jinkela_wire_169;
    wire new_Jinkela_wire_2510;
    wire n_0195_;
    wire new_Jinkela_wire_2286;
    wire new_Jinkela_wire_6513;
    wire new_Jinkela_wire_7030;
    wire new_Jinkela_wire_5405;
    wire n_0334_;
    wire n_0918_;
    wire new_Jinkela_wire_3851;
    wire new_Jinkela_wire_8797;
    wire new_Jinkela_wire_3767;
    wire new_Jinkela_wire_4011;
    wire new_Jinkela_wire_7372;
    wire new_Jinkela_wire_6117;
    wire new_Jinkela_wire_2391;
    wire n_0124_;
    wire new_Jinkela_wire_5595;
    wire new_Jinkela_wire_5978;
    wire new_Jinkela_wire_811;
    wire new_Jinkela_wire_5585;
    wire n_0322_;
    wire new_Jinkela_wire_5890;
    wire new_Jinkela_wire_4410;
    wire new_Jinkela_wire_1478;
    wire new_Jinkela_wire_1802;
    wire new_Jinkela_wire_254;
    wire new_Jinkela_wire_7756;
    wire new_Jinkela_wire_5699;
    wire new_Jinkela_wire_7554;
    wire n_0037_;
    wire new_Jinkela_wire_7700;
    wire new_Jinkela_wire_3405;
    wire n_0025_;
    wire new_Jinkela_wire_6395;
    wire new_Jinkela_wire_6096;
    wire new_Jinkela_wire_1907;
    wire new_Jinkela_wire_8270;
    wire new_Jinkela_wire_3463;
    wire new_Jinkela_wire_9414;
    wire new_Jinkela_wire_6462;
    wire new_Jinkela_wire_9504;
    wire new_Jinkela_wire_6945;
    wire new_Jinkela_wire_733;
    wire n_0472_;
    wire new_Jinkela_wire_6029;
    wire new_Jinkela_wire_1233;
    wire new_Jinkela_wire_4102;
    wire new_Jinkela_wire_3979;
    wire new_Jinkela_wire_9165;
    wire new_Jinkela_wire_474;
    wire n_0824_;
    wire new_Jinkela_wire_1961;
    wire new_Jinkela_wire_2533;
    wire new_Jinkela_wire_10466;
    wire new_Jinkela_wire_470;
    wire new_Jinkela_wire_590;
    wire new_Jinkela_wire_6676;
    wire new_Jinkela_wire_9289;
    wire new_Jinkela_wire_7231;
    wire new_Jinkela_wire_3768;
    wire new_Jinkela_wire_1836;
    wire new_Jinkela_wire_9987;
    wire new_Jinkela_wire_6255;
    wire new_Jinkela_wire_6618;
    wire n_0675_;
    wire new_Jinkela_wire_6901;
    wire new_Jinkela_wire_212;
    wire new_Jinkela_wire_2805;
    wire new_Jinkela_wire_1072;
    wire new_Jinkela_wire_10612;
    wire n_0061_;
    wire new_Jinkela_wire_8971;
    wire new_Jinkela_wire_191;
    wire new_Jinkela_wire_9867;
    wire new_Jinkela_wire_4029;
    wire new_Jinkela_wire_4785;
    wire new_Jinkela_wire_4777;
    wire new_Jinkela_wire_5519;
    wire new_Jinkela_wire_6430;
    wire n_0232_;
    wire new_Jinkela_wire_2672;
    wire new_Jinkela_wire_2241;
    wire n_0626_;
    wire new_Jinkela_wire_6964;
    wire new_Jinkela_wire_9635;
    wire new_Jinkela_wire_1964;
    wire new_Jinkela_wire_3093;
    wire new_Jinkela_wire_2395;
    wire new_Jinkela_wire_6375;
    wire new_Jinkela_wire_9947;
    wire new_Jinkela_wire_1581;
    wire new_Jinkela_wire_1508;
    wire new_Jinkela_wire_9469;
    wire new_Jinkela_wire_2836;
    wire new_Jinkela_wire_6143;
    wire new_Jinkela_wire_8980;
    wire new_Jinkela_wire_2516;
    wire n_0950_;
    wire new_Jinkela_wire_5106;
    wire new_Jinkela_wire_8200;
    wire new_Jinkela_wire_956;
    wire new_Jinkela_wire_2032;
    wire new_Jinkela_wire_3121;
    wire new_Jinkela_wire_4294;
    wire n_0735_;
    wire new_Jinkela_wire_2056;
    wire new_Jinkela_wire_5943;
    wire new_Jinkela_wire_1955;
    wire n_0884_;
    wire new_Jinkela_wire_7297;
    wire new_Jinkela_wire_7577;
    wire n_0830_;
    wire new_Jinkela_wire_1416;
    wire new_Jinkela_wire_6155;
    wire new_Jinkela_wire_4708;
    wire new_Jinkela_wire_5172;
    wire new_Jinkela_wire_4068;
    wire new_Jinkela_wire_10393;
    wire new_Jinkela_wire_10226;
    wire new_Jinkela_wire_6385;
    wire new_Jinkela_wire_4415;
    wire new_Jinkela_wire_3039;
    wire new_Jinkela_wire_2292;
    wire new_Jinkela_wire_5009;
    wire new_Jinkela_wire_10216;
    wire new_Jinkela_wire_4549;
    wire new_net_2525;
    wire new_Jinkela_wire_4272;
    wire new_Jinkela_wire_7811;
    wire new_Jinkela_wire_3297;
    wire new_Jinkela_wire_604;
    wire new_Jinkela_wire_4880;
    wire new_Jinkela_wire_6383;
    wire new_Jinkela_wire_6451;
    wire n_0078_;
    wire new_Jinkela_wire_75;
    wire n_0233_;
    wire new_Jinkela_wire_8349;
    wire new_Jinkela_wire_7440;
    wire new_Jinkela_wire_7610;
    wire new_Jinkela_wire_1982;
    wire new_Jinkela_wire_692;
    wire new_Jinkela_wire_255;
    wire new_Jinkela_wire_1505;
    wire new_Jinkela_wire_4577;
    wire new_Jinkela_wire_1223;
    wire new_Jinkela_wire_7485;
    wire new_Jinkela_wire_7640;
    wire new_Jinkela_wire_10622;
    wire new_Jinkela_wire_6525;
    wire new_Jinkela_wire_6276;
    wire new_Jinkela_wire_8065;
    wire new_Jinkela_wire_2206;
    wire n_1295_;
    wire new_Jinkela_wire_290;
    wire new_Jinkela_wire_5958;
    wire n_0525_;
    wire new_Jinkela_wire_1477;
    wire new_Jinkela_wire_8805;
    wire new_Jinkela_wire_7491;
    wire new_Jinkela_wire_1750;
    wire new_Jinkela_wire_9948;
    wire n_0259_;
    wire new_Jinkela_wire_8876;
    wire new_Jinkela_wire_2310;
    wire new_Jinkela_wire_3342;
    wire new_Jinkela_wire_5203;
    wire new_Jinkela_wire_9813;
    wire new_Jinkela_wire_536;
    wire new_Jinkela_wire_4203;
    wire new_Jinkela_wire_4705;
    wire new_Jinkela_wire_5725;
    wire new_Jinkela_wire_9182;
    wire new_Jinkela_wire_1956;
    wire new_Jinkela_wire_8939;
    wire new_Jinkela_wire_3483;
    wire new_Jinkela_wire_1485;
    wire n_1369_;
    wire new_Jinkela_wire_8013;
    wire new_Jinkela_wire_7190;
    wire new_Jinkela_wire_3224;
    wire new_Jinkela_wire_8903;
    wire new_Jinkela_wire_7951;
    wire n_0771_;
    wire n_0713_;
    wire new_Jinkela_wire_6998;
    wire new_Jinkela_wire_6278;
    wire new_Jinkela_wire_3795;
    wire new_Jinkela_wire_6104;
    wire new_Jinkela_wire_8699;
    wire new_Jinkela_wire_2986;
    wire new_Jinkela_wire_875;
    wire new_Jinkela_wire_9089;
    wire new_Jinkela_wire_1751;
    wire new_Jinkela_wire_6078;
    wire new_Jinkela_wire_619;
    wire new_Jinkela_wire_6524;
    wire new_Jinkela_wire_578;
    wire new_Jinkela_wire_2219;
    wire new_Jinkela_wire_7473;
    wire new_Jinkela_wire_814;
    wire new_Jinkela_wire_4170;
    wire new_Jinkela_wire_3714;
    wire new_Jinkela_wire_6583;
    wire new_Jinkela_wire_5552;
    wire new_Jinkela_wire_2052;
    wire new_Jinkela_wire_7020;
    wire new_Jinkela_wire_2288;
    wire new_Jinkela_wire_1783;
    wire new_Jinkela_wire_2663;
    wire new_Jinkela_wire_9181;
    wire new_Jinkela_wire_3377;
    wire new_Jinkela_wire_4723;
    wire new_Jinkela_wire_860;
    wire new_Jinkela_wire_4279;
    wire new_Jinkela_wire_2075;
    wire new_Jinkela_wire_5507;
    wire n_0181_;
    wire new_Jinkela_wire_2914;
    wire new_Jinkela_wire_3794;
    wire new_Jinkela_wire_8899;
    wire new_Jinkela_wire_336;
    wire new_Jinkela_wire_5054;
    wire new_Jinkela_wire_150;
    wire new_Jinkela_wire_1655;
    wire new_Jinkela_wire_8444;
    wire new_Jinkela_wire_3422;
    wire new_Jinkela_wire_6761;
    wire new_Jinkela_wire_8934;
    wire new_Jinkela_wire_3049;
    wire new_Jinkela_wire_1274;
    wire new_Jinkela_wire_3518;
    wire new_Jinkela_wire_2265;
    wire n_0351_;
    wire new_Jinkela_wire_5666;
    wire new_Jinkela_wire_2386;
    wire new_Jinkela_wire_10339;
    wire n_0649_;
    wire new_Jinkela_wire_6927;
    wire new_Jinkela_wire_5380;
    wire n_1118_;
    wire new_Jinkela_wire_22;
    wire new_Jinkela_wire_8012;
    wire new_Jinkela_wire_5853;
    wire new_Jinkela_wire_8896;
    wire new_Jinkela_wire_10503;
    wire new_Jinkela_wire_996;
    wire new_Jinkela_wire_1293;
    wire new_Jinkela_wire_5073;
    wire new_Jinkela_wire_4154;
    wire new_Jinkela_wire_4255;
    wire new_Jinkela_wire_5329;
    wire new_Jinkela_wire_3823;
    wire new_Jinkela_wire_3608;
    wire new_Jinkela_wire_9133;
    wire new_Jinkela_wire_3161;
    wire new_Jinkela_wire_4751;
    wire new_Jinkela_wire_865;
    wire new_Jinkela_wire_7646;
    wire new_Jinkela_wire_8166;
    wire new_Jinkela_wire_9882;
    wire new_Jinkela_wire_9653;
    wire n_0184_;
    wire new_Jinkela_wire_1562;
    wire new_Jinkela_wire_6209;
    wire new_Jinkela_wire_7303;
    wire n_1235_;
    wire new_Jinkela_wire_3408;
    wire n_1184_;
    wire new_Jinkela_wire_3697;
    wire new_Jinkela_wire_7094;
    wire new_Jinkela_wire_4001;
    wire new_Jinkela_wire_3675;
    wire new_Jinkela_wire_2728;
    wire new_Jinkela_wire_8319;
    wire new_Jinkela_wire_9994;
    wire new_Jinkela_wire_1928;
    wire new_Jinkela_wire_1406;
    wire new_Jinkela_wire_6268;
    wire new_Jinkela_wire_3092;
    wire new_Jinkela_wire_8762;
    wire new_Jinkela_wire_6568;
    wire new_Jinkela_wire_5880;
    wire new_Jinkela_wire_2520;
    wire new_Jinkela_wire_3940;
    wire new_Jinkela_wire_364;
    wire new_Jinkela_wire_357;
    wire new_Jinkela_wire_3672;
    wire n_0792_;
    wire new_Jinkela_wire_5474;
    wire new_Jinkela_wire_2093;
    wire new_Jinkela_wire_5415;
    wire new_Jinkela_wire_8858;
    wire new_Jinkela_wire_3569;
    wire new_Jinkela_wire_7170;
    wire new_Jinkela_wire_2410;
    wire new_Jinkela_wire_9759;
    wire new_Jinkela_wire_1204;
    wire new_Jinkela_wire_7789;
    wire n_0628_;
    wire new_Jinkela_wire_2166;
    wire new_Jinkela_wire_763;
    wire new_Jinkela_wire_10183;
    wire new_Jinkela_wire_9642;
    wire new_Jinkela_wire_5733;
    wire new_Jinkela_wire_3375;
    wire new_Jinkela_wire_9120;
    wire n_0596_;
    wire new_Jinkela_wire_1980;
    wire new_Jinkela_wire_6114;
    wire new_Jinkela_wire_9032;
    wire new_Jinkela_wire_2251;
    wire new_Jinkela_wire_8963;
    wire new_Jinkela_wire_4627;
    wire n_0931_;
    wire new_Jinkela_wire_5153;
    wire n_0907_;
    wire new_Jinkela_wire_8982;
    wire new_Jinkela_wire_2844;
    wire new_Jinkela_wire_348;
    wire new_Jinkela_wire_9734;
    wire new_Jinkela_wire_8960;
    wire new_Jinkela_wire_6717;
    wire new_Jinkela_wire_6694;
    wire new_Jinkela_wire_3053;
    wire new_Jinkela_wire_3850;
    wire new_Jinkela_wire_3901;
    wire new_Jinkela_wire_7486;
    wire new_Jinkela_wire_366;
    wire new_Jinkela_wire_7353;
    wire new_Jinkela_wire_8710;
    wire n_0928_;
    wire new_Jinkela_wire_1742;
    wire new_Jinkela_wire_4269;
    wire new_Jinkela_wire_8322;
    wire new_Jinkela_wire_9188;
    wire n_0826_;
    wire new_Jinkela_wire_8007;
    wire new_Jinkela_wire_8069;
    wire new_Jinkela_wire_9147;
    wire new_Jinkela_wire_1567;
    wire n_1179_;
    wire new_Jinkela_wire_2228;
    wire new_Jinkela_wire_10526;
    wire new_Jinkela_wire_8093;
    wire new_Jinkela_wire_7739;
    wire n_1324_;
    wire n_0601_;
    wire new_Jinkela_wire_1297;
    wire new_Jinkela_wire_8656;
    wire new_Jinkela_wire_7677;
    wire new_Jinkela_wire_9798;
    wire new_Jinkela_wire_7613;
    wire new_Jinkela_wire_9632;
    wire new_Jinkela_wire_199;
    wire new_Jinkela_wire_4774;
    wire new_Jinkela_wire_9868;
    wire new_Jinkela_wire_8263;
    wire new_Jinkela_wire_1101;
    wire new_Jinkela_wire_7086;
    wire new_Jinkela_wire_9185;
    wire new_Jinkela_wire_3332;
    wire n_0637_;
    wire new_Jinkela_wire_2945;
    wire new_Jinkela_wire_2194;
    wire new_Jinkela_wire_6894;
    wire new_Jinkela_wire_537;
    wire new_Jinkela_wire_7446;
    wire new_Jinkela_wire_4652;
    wire new_Jinkela_wire_2838;
    wire new_Jinkela_wire_6976;
    wire new_Jinkela_wire_6752;
    wire new_Jinkela_wire_4499;
    wire new_Jinkela_wire_2389;
    wire new_Jinkela_wire_2560;
    wire new_Jinkela_wire_422;
    wire new_Jinkela_wire_228;
    wire n_0998_;
    wire n_0518_;
    wire new_Jinkela_wire_9748;
    wire new_Jinkela_wire_7405;
    wire new_Jinkela_wire_551;
    wire new_Jinkela_wire_4760;
    wire new_Jinkela_wire_2394;
    wire new_Jinkela_wire_3700;
    wire new_Jinkela_wire_2747;
    wire new_Jinkela_wire_8717;
    wire new_Jinkela_wire_8080;
    wire new_Jinkela_wire_7076;
    wire new_Jinkela_wire_9524;
    wire new_Jinkela_wire_3515;
    wire new_Jinkela_wire_6795;
    wire new_Jinkela_wire_5897;
    wire new_Jinkela_wire_479;
    wire new_Jinkela_wire_10285;
    wire new_Jinkela_wire_6021;
    wire new_Jinkela_wire_5001;
    wire new_Jinkela_wire_7070;
    wire new_Jinkela_wire_1936;
    wire new_Jinkela_wire_4813;
    wire n_0188_;
    wire new_Jinkela_wire_3310;
    wire new_Jinkela_wire_980;
    wire new_Jinkela_wire_5450;
    wire new_Jinkela_wire_1474;
    wire new_Jinkela_wire_4200;
    wire new_Jinkela_wire_4297;
    wire new_Jinkela_wire_7445;
    wire new_Jinkela_wire_6141;
    wire new_Jinkela_wire_4539;
    wire new_Jinkela_wire_8311;
    wire new_Jinkela_wire_5597;
    wire new_Jinkela_wire_3189;
    wire n_0066_;
    wire new_Jinkela_wire_1026;
    wire new_Jinkela_wire_6824;
    wire new_Jinkela_wire_10246;
    wire new_Jinkela_wire_6776;
    wire new_Jinkela_wire_7752;
    wire new_Jinkela_wire_9638;
    wire new_Jinkela_wire_3598;
    wire new_Jinkela_wire_3780;
    wire new_Jinkela_wire_5607;
    wire new_Jinkela_wire_9107;
    wire new_Jinkela_wire_5744;
    wire new_Jinkela_wire_7331;
    wire new_Jinkela_wire_5204;
    wire new_Jinkela_wire_8583;
    wire new_Jinkela_wire_8673;
    wire new_net_2497;
    wire new_Jinkela_wire_9831;
    wire new_Jinkela_wire_5821;
    wire new_Jinkela_wire_4453;
    wire new_Jinkela_wire_7414;
    wire new_Jinkela_wire_2358;
    wire new_Jinkela_wire_8104;
    wire new_Jinkela_wire_5982;
    wire new_Jinkela_wire_9940;
    wire new_Jinkela_wire_3991;
    wire new_Jinkela_wire_626;
    wire new_Jinkela_wire_2694;
    wire new_Jinkela_wire_6863;
    wire new_Jinkela_wire_2277;
    wire new_Jinkela_wire_7400;
    wire new_Jinkela_wire_2361;
    wire new_Jinkela_wire_8064;
    wire new_Jinkela_wire_9376;
    wire new_Jinkela_wire_1305;
    wire new_Jinkela_wire_1708;
    wire new_Jinkela_wire_6166;
    wire new_Jinkela_wire_7781;
    wire new_Jinkela_wire_9444;
    wire new_Jinkela_wire_10445;
    wire new_Jinkela_wire_7982;
    wire new_Jinkela_wire_10214;
    wire new_Jinkela_wire_762;
    wire new_Jinkela_wire_748;
    wire new_Jinkela_wire_7063;
    wire new_Jinkela_wire_4205;
    wire new_Jinkela_wire_1983;
    wire new_Jinkela_wire_8975;
    wire n_0015_;
    wire new_Jinkela_wire_7624;
    wire new_Jinkela_wire_10054;
    wire new_Jinkela_wire_4378;
    wire new_Jinkela_wire_7180;
    wire new_Jinkela_wire_4517;
    wire new_Jinkela_wire_7566;
    wire new_Jinkela_wire_9458;
    wire new_Jinkela_wire_4959;
    wire new_Jinkela_wire_4131;
    wire new_Jinkela_wire_3384;
    wire new_Jinkela_wire_2332;
    wire new_Jinkela_wire_9963;
    wire new_Jinkela_wire_4226;
    wire new_Jinkela_wire_8729;
    wire new_Jinkela_wire_892;
    wire new_Jinkela_wire_2270;
    wire new_Jinkela_wire_6182;
    wire new_Jinkela_wire_10017;
    wire new_Jinkela_wire_6794;
    wire new_Jinkela_wire_424;
    wire new_Jinkela_wire_6411;
    wire new_Jinkela_wire_10245;
    wire new_Jinkela_wire_6948;
    wire n_0005_;
    wire new_Jinkela_wire_1350;
    wire n_0718_;
    wire new_Jinkela_wire_8083;
    wire new_Jinkela_wire_9453;
    wire new_Jinkela_wire_7326;
    wire n_0235_;
    wire new_Jinkela_wire_3511;
    wire new_Jinkela_wire_8590;
    wire new_Jinkela_wire_4555;
    wire new_Jinkela_wire_6248;
    wire new_Jinkela_wire_8439;
    wire new_Jinkela_wire_8833;
    wire new_Jinkela_wire_3964;
    wire new_Jinkela_wire_8889;
    wire n_0887_;
    wire new_Jinkela_wire_6663;
    wire new_Jinkela_wire_928;
    wire new_Jinkela_wire_9079;
    wire new_Jinkela_wire_8118;
    wire new_Jinkela_wire_10248;
    wire new_Jinkela_wire_3997;
    wire new_Jinkela_wire_6482;
    wire new_Jinkela_wire_9819;
    wire new_Jinkela_wire_4401;
    wire new_Jinkela_wire_4195;
    wire new_Jinkela_wire_1271;
    wire new_Jinkela_wire_5177;
    wire new_Jinkela_wire_0;
    wire new_Jinkela_wire_654;
    wire new_Jinkela_wire_1330;
    wire new_Jinkela_wire_8136;
    wire new_Jinkela_wire_674;
    wire new_Jinkela_wire_3254;
    wire new_Jinkela_wire_6680;
    wire new_Jinkela_wire_3956;
    wire n_1209_;
    wire new_Jinkela_wire_4661;
    wire new_Jinkela_wire_1634;
    wire new_Jinkela_wire_7969;
    wire new_Jinkela_wire_925;
    wire n_1107_;
    wire new_Jinkela_wire_451;
    wire new_Jinkela_wire_9942;
    wire new_Jinkela_wire_1341;
    wire new_Jinkela_wire_3996;
    wire new_Jinkela_wire_6082;
    wire new_Jinkela_wire_4726;
    wire new_Jinkela_wire_62;
    wire new_Jinkela_wire_4930;
    wire n_0537_;
    wire n_0511_;
    wire new_Jinkela_wire_9068;
    wire new_Jinkela_wire_757;
    wire new_Jinkela_wire_7715;
    wire n_1038_;
    wire n_0582_;
    wire new_Jinkela_wire_4353;
    wire new_Jinkela_wire_7786;
    wire new_Jinkela_wire_9461;
    wire new_Jinkela_wire_6812;
    wire new_Jinkela_wire_1801;
    wire n_0295_;
    wire new_Jinkela_wire_2538;
    wire new_Jinkela_wire_6632;
    wire new_Jinkela_wire_7238;
    wire new_Jinkela_wire_9750;
    wire new_Jinkela_wire_5599;
    wire new_Jinkela_wire_3650;
    wire new_Jinkela_wire_4940;
    wire new_Jinkela_wire_689;
    wire new_Jinkela_wire_8950;
    wire new_Jinkela_wire_10602;
    wire new_Jinkela_wire_1215;
    wire new_Jinkela_wire_3752;
    wire new_Jinkela_wire_8023;
    wire new_Jinkela_wire_6432;
    wire new_Jinkela_wire_8991;
    wire new_Jinkela_wire_4278;
    wire new_Jinkela_wire_6322;
    wire new_Jinkela_wire_7263;
    wire new_Jinkela_wire_9477;
    wire new_Jinkela_wire_8686;
    wire new_Jinkela_wire_2132;
    wire new_Jinkela_wire_3262;
    wire new_Jinkela_wire_4136;
    wire n_1016_;
    wire new_Jinkela_wire_4749;
    wire new_Jinkela_wire_2403;
    wire new_Jinkela_wire_566;
    wire new_Jinkela_wire_4302;
    wire new_Jinkela_wire_7816;
    wire new_Jinkela_wire_344;
    wire new_Jinkela_wire_6404;
    wire new_Jinkela_wire_10455;
    wire new_Jinkela_wire_3984;
    wire new_Jinkela_wire_10217;
    wire new_Jinkela_wire_3830;
    wire new_Jinkela_wire_6833;
    wire n_0530_;
    wire new_Jinkela_wire_1392;
    wire new_Jinkela_wire_2300;
    wire new_Jinkela_wire_7363;
    wire new_Jinkela_wire_9006;
    wire new_Jinkela_wire_352;
    wire new_Jinkela_wire_5771;
    wire new_Jinkela_wire_5080;
    wire new_Jinkela_wire_2442;
    wire new_Jinkela_wire_4842;
    wire new_Jinkela_wire_7588;
    wire new_Jinkela_wire_2894;
    wire new_Jinkela_wire_9523;
    wire new_Jinkela_wire_5276;
    wire n_0014_;
    wire new_Jinkela_wire_2719;
    wire new_Jinkela_wire_893;
    wire new_Jinkela_wire_10153;
    wire new_Jinkela_wire_2511;
    wire new_Jinkela_wire_7810;
    wire new_Jinkela_wire_4082;
    wire new_Jinkela_wire_492;
    wire new_Jinkela_wire_1461;
    wire new_Jinkela_wire_826;
    wire new_Jinkela_wire_2263;
    wire new_Jinkela_wire_8519;
    wire new_Jinkela_wire_2509;
    wire new_Jinkela_wire_7547;
    wire new_Jinkela_wire_10112;
    wire new_Jinkela_wire_7697;
    wire new_Jinkela_wire_9473;
    wire new_Jinkela_wire_6635;
    wire new_Jinkela_wire_8112;
    wire new_Jinkela_wire_10520;
    wire n_1246_;
    wire new_Jinkela_wire_6109;
    wire new_Jinkela_wire_672;
    wire new_Jinkela_wire_1917;
    wire n_0778_;
    wire new_Jinkela_wire_2611;
    wire new_Jinkela_wire_6484;
    wire new_Jinkela_wire_9575;
    wire new_Jinkela_wire_4922;
    wire new_Jinkela_wire_7532;
    wire n_0269_;
    wire new_Jinkela_wire_3164;
    wire new_Jinkela_wire_669;
    wire new_Jinkela_wire_2211;
    wire new_Jinkela_wire_2623;
    wire new_Jinkela_wire_436;
    wire new_Jinkela_wire_1429;
    wire new_Jinkela_wire_4733;
    wire new_Jinkela_wire_1021;
    wire new_Jinkela_wire_7884;
    wire new_Jinkela_wire_114;
    wire new_Jinkela_wire_8781;
    wire new_Jinkela_wire_3942;
    wire new_Jinkela_wire_8821;
    wire n_1289_;
    wire new_Jinkela_wire_8281;
    wire new_Jinkela_wire_903;
    wire new_Jinkela_wire_8665;
    wire new_Jinkela_wire_2985;
    wire new_Jinkela_wire_307;
    wire n_1068_;
    wire new_Jinkela_wire_3831;
    wire new_Jinkela_wire_10199;
    wire new_Jinkela_wire_4303;
    wire new_Jinkela_wire_10628;
    wire new_Jinkela_wire_6810;
    wire new_Jinkela_wire_5520;
    wire new_Jinkela_wire_8500;
    wire new_Jinkela_wire_313;
    wire new_Jinkela_wire_1571;
    wire new_Jinkela_wire_1475;
    wire new_Jinkela_wire_7114;
    wire new_Jinkela_wire_2711;
    wire new_Jinkela_wire_7222;
    wire new_Jinkela_wire_9078;
    wire new_Jinkela_wire_2247;
    wire new_Jinkela_wire_8036;
    wire new_Jinkela_wire_9967;
    wire new_Jinkela_wire_3220;
    wire n_0947_;
    wire new_Jinkela_wire_4046;
    wire new_Jinkela_wire_10454;
    wire new_Jinkela_wire_4002;
    wire new_Jinkela_wire_5598;
    wire new_Jinkela_wire_9624;
    wire new_Jinkela_wire_1315;
    wire n_1083_;
    wire new_Jinkela_wire_1251;
    wire new_Jinkela_wire_3975;
    wire n_0021_;
    wire new_Jinkela_wire_4786;
    wire new_net_2578;
    wire new_Jinkela_wire_3957;
    wire new_Jinkela_wire_6080;
    wire new_Jinkela_wire_8360;
    wire new_Jinkela_wire_9879;
    wire new_Jinkela_wire_3264;
    wire new_net_2566;
    wire new_Jinkela_wire_1222;
    wire new_Jinkela_wire_4188;
    wire new_Jinkela_wire_200;
    wire new_Jinkela_wire_167;
    wire new_Jinkela_wire_7513;
    wire new_Jinkela_wire_6978;
    wire new_Jinkela_wire_6357;
    wire new_Jinkela_wire_4788;
    wire new_Jinkela_wire_1294;
    wire new_Jinkela_wire_2111;
    wire new_Jinkela_wire_2136;
    wire new_Jinkela_wire_10076;
    wire new_Jinkela_wire_6158;
    wire new_Jinkela_wire_7778;
    wire new_Jinkela_wire_605;
    wire n_0246_;
    wire new_Jinkela_wire_7757;
    wire new_Jinkela_wire_720;
    wire new_Jinkela_wire_4443;
    wire new_Jinkela_wire_7387;
    wire new_Jinkela_wire_522;
    wire n_0993_;
    wire new_Jinkela_wire_2998;
    wire n_0288_;
    wire new_Jinkela_wire_2693;
    wire new_Jinkela_wire_4587;
    wire new_Jinkela_wire_7162;
    wire new_Jinkela_wire_8050;
    wire n_0299_;
    wire new_Jinkela_wire_6954;
    wire n_1078_;
    wire new_Jinkela_wire_7527;
    wire new_Jinkela_wire_3;
    wire new_Jinkela_wire_8418;
    wire new_Jinkela_wire_6298;
    wire new_Jinkela_wire_9263;
    wire new_Jinkela_wire_5130;
    wire new_Jinkela_wire_644;
    wire new_Jinkela_wire_3730;
    wire new_Jinkela_wire_10365;
    wire new_Jinkela_wire_8987;
    wire new_Jinkela_wire_326;
    wire new_Jinkela_wire_5784;
    wire new_Jinkela_wire_5418;
    wire new_Jinkela_wire_9051;
    wire n_1252_;
    wire new_Jinkela_wire_8572;
    wire new_Jinkela_wire_3376;
    wire new_Jinkela_wire_9964;
    wire new_Jinkela_wire_2807;
    wire new_Jinkela_wire_2373;
    wire new_Jinkela_wire_1731;
    wire new_Jinkela_wire_5470;
    wire new_Jinkela_wire_7185;
    wire new_Jinkela_wire_1405;
    wire n_0756_;
    wire new_Jinkela_wire_817;
    wire new_Jinkela_wire_5086;
    wire n_0375_;
    wire new_Jinkela_wire_2846;
    wire new_Jinkela_wire_10200;
    wire new_Jinkela_wire_1041;
    wire new_Jinkela_wire_8148;
    wire new_Jinkela_wire_5482;
    wire new_Jinkela_wire_1681;
    wire new_Jinkela_wire_5151;
    wire new_Jinkela_wire_1132;
    wire new_Jinkela_wire_2790;
    wire new_Jinkela_wire_2770;
    wire new_Jinkela_wire_9245;
    wire new_Jinkela_wire_4642;
    wire new_Jinkela_wire_6533;
    wire new_Jinkela_wire_9896;
    wire new_Jinkela_wire_2275;
    wire new_Jinkela_wire_4801;
    wire new_Jinkela_wire_6279;
    wire new_Jinkela_wire_9958;
    wire new_Jinkela_wire_6181;
    wire new_Jinkela_wire_10405;
    wire new_Jinkela_wire_4759;
    wire new_Jinkela_wire_10465;
    wire new_Jinkela_wire_2757;
    wire new_Jinkela_wire_6033;
    wire new_Jinkela_wire_10071;
    wire new_Jinkela_wire_6793;
    wire new_Jinkela_wire_1160;
    wire new_Jinkela_wire_207;
    wire new_Jinkela_wire_8355;
    wire new_Jinkela_wire_1504;
    wire new_Jinkela_wire_5548;
    wire new_Jinkela_wire_10580;
    wire new_Jinkela_wire_5851;
    wire new_Jinkela_wire_7335;
    wire n_0436_;
    wire new_Jinkela_wire_1895;
    wire new_Jinkela_wire_7397;
    wire new_Jinkela_wire_10316;
    wire new_Jinkela_wire_5631;
    wire new_Jinkela_wire_6958;
    wire new_Jinkela_wire_6000;
    wire new_Jinkela_wire_6757;
    wire n_1189_;
    wire new_Jinkela_wire_416;
    wire new_Jinkela_wire_1347;
    wire new_Jinkela_wire_4985;
    wire n_0502_;
    wire new_Jinkela_wire_5306;
    wire new_Jinkela_wire_10418;
    wire new_Jinkela_wire_20;
    wire new_Jinkela_wire_5392;
    wire new_Jinkela_wire_3595;
    wire new_Jinkela_wire_7783;
    wire new_Jinkela_wire_3271;
    wire new_Jinkela_wire_2612;
    wire new_Jinkela_wire_8457;
    wire new_Jinkela_wire_3258;
    wire new_Jinkela_wire_9701;
    wire new_Jinkela_wire_1604;
    wire new_Jinkela_wire_3516;
    wire n_0989_;
    wire new_Jinkela_wire_6017;
    wire new_Jinkela_wire_463;
    wire n_0749_;
    wire new_Jinkela_wire_6673;
    wire new_Jinkela_wire_6502;
    wire new_Jinkela_wire_808;
    wire new_Jinkela_wire_2588;
    wire n_0137_;
    wire new_Jinkela_wire_3872;
    wire new_Jinkela_wire_7762;
    wire new_Jinkela_wire_1117;
    wire new_Jinkela_wire_9090;
    wire new_Jinkela_wire_6892;
    wire new_Jinkela_wire_1868;
    wire new_Jinkela_wire_6163;
    wire new_Jinkela_wire_6719;
    wire new_Jinkela_wire_8541;
    wire new_Jinkela_wire_5282;
    wire new_Jinkela_wire_1438;
    wire new_Jinkela_wire_4038;
    wire new_Jinkela_wire_8554;
    wire new_Jinkela_wire_8204;
    wire new_Jinkela_wire_1413;
    wire new_Jinkela_wire_3821;
    wire new_Jinkela_wire_3755;
    wire new_Jinkela_wire_2319;
    wire new_Jinkela_wire_8414;
    wire new_Jinkela_wire_6908;
    wire new_Jinkela_wire_1710;
    wire new_Jinkela_wire_1524;
    wire new_Jinkela_wire_9310;
    wire new_Jinkela_wire_3465;
    wire new_Jinkela_wire_7003;
    wire new_Jinkela_wire_3501;
    wire new_Jinkela_wire_7133;
    wire new_Jinkela_wire_10137;
    wire new_Jinkela_wire_9528;
    wire new_Jinkela_wire_7959;
    wire new_Jinkela_wire_6428;
    wire new_Jinkela_wire_3076;
    wire new_Jinkela_wire_10293;
    wire new_Jinkela_wire_109;
    wire new_Jinkela_wire_3970;
    wire new_Jinkela_wire_1313;
    wire n_1229_;
    wire new_Jinkela_wire_4166;
    wire new_Jinkela_wire_761;
    wire n_0744_;
    wire new_Jinkela_wire_4388;
    wire new_Jinkela_wire_420;
    wire new_Jinkela_wire_5393;
    wire new_Jinkela_wire_8695;
    wire new_Jinkela_wire_4714;
    wire n_1337_;
    wire new_Jinkela_wire_1872;
    wire new_Jinkela_wire_2447;
    wire new_Jinkela_wire_4515;
    wire new_Jinkela_wire_10601;
    wire new_Jinkela_wire_3356;
    wire new_Jinkela_wire_6977;
    wire new_Jinkela_wire_1552;
    wire n_0706_;
    wire new_Jinkela_wire_5966;
    wire new_Jinkela_wire_2967;
    wire new_Jinkela_wire_2690;
    wire new_Jinkela_wire_7479;
    wire new_Jinkela_wire_431;
    wire new_Jinkela_wire_10439;
    wire new_Jinkela_wire_1503;
    wire n_0070_;
    wire n_0143_;
    wire n_0865_;
    wire new_Jinkela_wire_3918;
    wire new_Jinkela_wire_7205;
    wire n_0141_;
    wire new_Jinkela_wire_4201;
    wire new_Jinkela_wire_7193;
    wire new_Jinkela_wire_9870;
    wire new_Jinkela_wire_8814;
    wire new_Jinkela_wire_9646;
    wire new_Jinkela_wire_8513;
    wire n_0796_;
    wire new_Jinkela_wire_4273;
    wire new_Jinkela_wire_1583;
    wire new_Jinkela_wire_3361;
    wire new_Jinkela_wire_9380;
    wire new_Jinkela_wire_5210;
    wire new_Jinkela_wire_6573;
    wire new_Jinkela_wire_8548;
    wire new_Jinkela_wire_8809;
    wire n_0227_;
    wire new_Jinkela_wire_7818;
    wire new_Jinkela_wire_3715;
    wire n_0024_;
    wire n_1110_;
    wire new_Jinkela_wire_4781;
    wire new_Jinkela_wire_3658;
    wire new_Jinkela_wire_7978;
    wire new_Jinkela_wire_2800;
    wire n_0786_;
    wire new_Jinkela_wire_682;
    wire new_Jinkela_wire_9448;
    wire new_Jinkela_wire_10023;
    wire new_Jinkela_wire_508;
    wire new_Jinkela_wire_5749;
    wire new_Jinkela_wire_8792;
    wire new_Jinkela_wire_2456;
    wire new_Jinkela_wire_2177;
    wire new_Jinkela_wire_4716;
    wire new_Jinkela_wire_9116;
    wire n_1044_;
    wire new_Jinkela_wire_3651;
    wire new_Jinkela_wire_7956;
    wire new_Jinkela_wire_1851;
    wire new_Jinkela_wire_26;
    wire new_Jinkela_wire_10225;
    wire n_0754_;
    wire new_Jinkela_wire_10559;
    wire n_0707_;
    wire new_Jinkela_wire_2354;
    wire n_0922_;
    wire n_0466_;
    wire new_Jinkela_wire_2108;
    wire new_Jinkela_wire_1526;
    wire new_Jinkela_wire_910;
    wire new_Jinkela_wire_9544;
    wire new_Jinkela_wire_4285;
    wire new_Jinkela_wire_4754;
    wire new_Jinkela_wire_4757;
    wire n_0348_;
    wire new_Jinkela_wire_6865;
    wire new_Jinkela_wire_301;
    wire n_0278_;
    wire new_Jinkela_wire_8864;
    wire new_Jinkela_wire_8142;
    wire new_Jinkela_wire_5271;
    wire new_Jinkela_wire_8398;
    wire new_Jinkela_wire_7033;
    wire new_Jinkela_wire_4900;
    wire new_Jinkela_wire_4849;
    wire new_Jinkela_wire_9044;
    wire new_Jinkela_wire_5565;
    wire n_0394_;
    wire new_Jinkela_wire_6702;
    wire n_0485_;
    wire new_Jinkela_wire_3358;
    wire n_1136_;
    wire new_Jinkela_wire_3591;
    wire new_Jinkela_wire_7695;
    wire new_Jinkela_wire_7418;
    wire new_Jinkela_wire_6830;
    wire new_Jinkela_wire_1863;
    wire new_Jinkela_wire_984;
    wire new_Jinkela_wire_3480;
    wire new_Jinkela_wire_1077;
    wire new_Jinkela_wire_2916;
    wire new_Jinkela_wire_8691;
    wire new_Jinkela_wire_2801;
    wire new_Jinkela_wire_7497;
    wire new_Jinkela_wire_800;
    wire new_Jinkela_wire_1455;
    wire new_Jinkela_wire_46;
    wire new_Jinkela_wire_8345;
    wire new_Jinkela_wire_2198;
    wire new_Jinkela_wire_1263;
    wire new_Jinkela_wire_7299;
    wire new_Jinkela_wire_7362;
    wire new_Jinkela_wire_7967;
    wire new_Jinkela_wire_1966;
    wire new_Jinkela_wire_6448;
    wire new_Jinkela_wire_8033;
    wire new_Jinkela_wire_8994;
    wire new_Jinkela_wire_5976;
    wire new_Jinkela_wire_6737;
    wire new_Jinkela_wire_6466;
    wire new_Jinkela_wire_189;
    wire new_Jinkela_wire_2053;
    wire n_0941_;
    wire new_Jinkela_wire_3136;
    wire new_Jinkela_wire_8260;
    wire new_Jinkela_wire_5942;
    wire new_Jinkela_wire_6409;
    wire new_Jinkela_wire_3877;
    wire new_Jinkela_wire_5849;
    wire new_Jinkela_wire_7602;
    wire new_Jinkela_wire_407;
    wire new_Jinkela_wire_2231;
    wire new_Jinkela_wire_86;
    wire n_0742_;
    wire new_Jinkela_wire_5524;
    wire new_Jinkela_wire_2651;
    wire new_Jinkela_wire_2333;
    wire new_Jinkela_wire_7553;
    wire new_Jinkela_wire_4914;
    wire new_Jinkela_wire_10585;
    wire n_1127_;
    wire new_Jinkela_wire_2983;
    wire n_0807_;
    wire n_1071_;
    wire new_Jinkela_wire_10271;
    wire new_Jinkela_wire_6882;
    wire new_Jinkela_wire_1595;
    wire new_Jinkela_wire_842;
    wire new_Jinkela_wire_8463;
    wire new_Jinkela_wire_1880;
    wire n_0500_;
    wire new_Jinkela_wire_898;
    wire new_Jinkela_wire_1031;
    wire new_Jinkela_wire_5702;
    wire new_Jinkela_wire_5901;
    wire new_Jinkela_wire_5010;
    wire new_Jinkela_wire_7933;
    wire new_Jinkela_wire_4829;
    wire new_Jinkela_wire_4942;
    wire n_0440_;
    wire new_Jinkela_wire_4929;
    wire new_Jinkela_wire_226;
    wire new_Jinkela_wire_10094;
    wire new_Jinkela_wire_10432;
    wire new_Jinkela_wire_1374;
    wire new_Jinkela_wire_683;
    wire n_0581_;
    wire new_Jinkela_wire_3641;
    wire new_Jinkela_wire_1034;
    wire new_Jinkela_wire_1375;
    wire new_Jinkela_wire_1449;
    wire new_Jinkela_wire_1705;
    wire new_Jinkela_wire_4671;
    wire new_Jinkela_wire_6509;
    wire new_Jinkela_wire_8352;
    wire new_Jinkela_wire_3085;
    wire new_Jinkela_wire_662;
    wire new_Jinkela_wire_2463;
    wire new_Jinkela_wire_4752;
    wire n_0337_;
    wire new_Jinkela_wire_5433;
    wire new_Jinkela_wire_1894;
    wire new_Jinkela_wire_7725;
    wire new_Jinkela_wire_2551;
    wire new_Jinkela_wire_4312;
    wire new_Jinkela_wire_5850;
    wire new_Jinkela_wire_7681;
    wire n_0775_;
    wire new_Jinkela_wire_2909;
    wire new_Jinkela_wire_899;
    wire new_Jinkela_wire_1394;
    wire new_Jinkela_wire_736;
    wire new_Jinkela_wire_4660;
    wire new_Jinkela_wire_2375;
    wire new_Jinkela_wire_9579;
    wire new_Jinkela_wire_5795;
    wire new_Jinkela_wire_2815;
    wire n_0810_;
    wire new_Jinkela_wire_5858;
    wire new_Jinkela_wire_5460;
    wire new_Jinkela_wire_8568;
    wire new_Jinkela_wire_8758;
    wire new_Jinkela_wire_3421;
    wire new_Jinkela_wire_990;
    wire new_Jinkela_wire_7784;
    wire new_Jinkela_wire_10348;
    wire new_Jinkela_wire_3913;
    wire new_Jinkela_wire_5629;
    wire n_0354_;
    wire n_0319_;
    wire new_Jinkela_wire_10621;
    wire new_Jinkela_wire_1719;
    wire new_Jinkela_wire_124;
    wire new_Jinkela_wire_2647;
    wire new_Jinkela_wire_1192;
    wire n_0940_;
    wire new_Jinkela_wire_6075;
    wire new_Jinkela_wire_3296;
    wire n_1052_;
    wire new_Jinkela_wire_5227;
    wire new_Jinkela_wire_139;
    wire new_Jinkela_wire_10048;
    wire new_Jinkela_wire_9166;
    wire new_Jinkela_wire_3790;
    wire new_Jinkela_wire_6916;
    wire new_Jinkela_wire_2828;
    wire new_Jinkela_wire_2339;
    wire new_Jinkela_wire_5662;
    wire new_Jinkela_wire_7531;
    wire new_Jinkela_wire_9285;
    wire new_Jinkela_wire_1570;
    wire new_Jinkela_wire_7753;
    wire new_Jinkela_wire_5980;
    wire n_1254_;
    wire new_Jinkela_wire_5963;
    wire new_Jinkela_wire_2291;
    wire new_Jinkela_wire_6234;
    wire new_Jinkela_wire_3407;
    wire new_Jinkela_wire_5522;
    wire new_Jinkela_wire_3878;
    wire new_Jinkela_wire_6192;
    wire new_Jinkela_wire_10041;
    wire new_Jinkela_wire_6707;
    wire n_0943_;
    wire new_Jinkela_wire_4820;
    wire new_Jinkela_wire_6605;
    wire new_Jinkela_wire_2335;
    wire new_Jinkela_wire_7946;
    wire new_Jinkela_wire_5924;
    wire new_Jinkela_wire_9307;
    wire new_Jinkela_wire_5431;
    wire n_1258_;
    wire new_Jinkela_wire_6187;
    wire new_Jinkela_wire_6120;
    wire new_Jinkela_wire_3128;
    wire new_Jinkela_wire_5077;
    wire new_Jinkela_wire_5544;
    wire n_1119_;
    wire new_Jinkela_wire_3077;
    wire new_Jinkela_wire_2276;
    wire new_Jinkela_wire_8206;
    wire new_Jinkela_wire_8379;
    wire n_0633_;
    wire new_Jinkela_wire_2134;
    wire n_0808_;
    wire new_Jinkela_wire_6736;
    wire new_Jinkela_wire_8362;
    wire new_Jinkela_wire_4495;
    wire new_Jinkela_wire_7194;
    wire new_Jinkela_wire_8827;
    wire new_Jinkela_wire_625;
    wire new_Jinkela_wire_3288;
    wire new_Jinkela_wire_876;
    wire new_Jinkela_wire_8553;
    wire new_Jinkela_wire_6418;
    wire n_0556_;
    wire new_Jinkela_wire_7570;
    wire new_Jinkela_wire_9619;
    wire new_Jinkela_wire_7164;
    wire n_0225_;
    wire new_Jinkela_wire_4531;
    wire new_Jinkela_wire_9474;
    wire new_Jinkela_wire_6868;
    wire new_Jinkela_wire_4996;
    wire new_Jinkela_wire_5515;
    wire new_Jinkela_wire_2756;
    wire new_Jinkela_wire_7537;
    wire new_Jinkela_wire_446;
    wire new_Jinkela_wire_9445;
    wire new_Jinkela_wire_5956;
    wire new_Jinkela_wire_6032;
    wire new_Jinkela_wire_829;
    wire new_Jinkela_wire_8018;
    wire new_Jinkela_wire_4371;
    wire new_Jinkela_wire_186;
    wire n_1011_;
    wire new_Jinkela_wire_9782;
    wire new_Jinkela_wire_3098;
    wire new_Jinkela_wire_3392;
    wire new_Jinkela_wire_4846;
    wire new_Jinkela_wire_6515;
    wire new_Jinkela_wire_3314;
    wire new_Jinkela_wire_8114;
    wire new_Jinkela_wire_5800;
    wire new_Jinkela_wire_10504;
    wire new_Jinkela_wire_5665;
    wire new_Jinkela_wire_4574;
    wire new_Jinkela_wire_9961;
    wire new_Jinkela_wire_4268;
    wire new_Jinkela_wire_6823;
    wire new_Jinkela_wire_4240;
    wire new_Jinkela_wire_9067;
    wire new_Jinkela_wire_8477;
    wire new_Jinkela_wire_9806;
    wire n_1166_;
    wire new_Jinkela_wire_2971;
    wire new_Jinkela_wire_4462;
    wire new_Jinkela_wire_8878;
    wire new_Jinkela_wire_6820;
    wire new_Jinkela_wire_4767;
    wire new_Jinkela_wire_1447;
    wire new_Jinkela_wire_2061;
    wire new_Jinkela_wire_4347;
    wire new_Jinkela_wire_4452;
    wire new_Jinkela_wire_6111;
    wire new_Jinkela_wire_7858;
    wire new_Jinkela_wire_3034;
    wire new_Jinkela_wire_693;
    wire new_Jinkela_wire_5532;
    wire new_Jinkela_wire_1775;
    wire new_Jinkela_wire_6162;
    wire new_Jinkela_wire_5033;
    wire new_Jinkela_wire_5667;
    wire new_Jinkela_wire_4121;
    wire n_0159_;
    wire new_Jinkela_wire_3104;
    wire new_Jinkela_wire_4730;
    wire n_0116_;
    wire new_Jinkela_wire_8768;
    wire new_Jinkela_wire_3601;
    wire new_Jinkela_wire_540;
    wire new_Jinkela_wire_732;
    wire new_Jinkela_wire_9589;
    wire n_0378_;
    wire new_Jinkela_wire_7365;
    wire n_0589_;
    wire new_Jinkela_wire_6165;
    wire new_Jinkela_wire_6494;
    wire new_Jinkela_wire_10412;
    wire new_Jinkela_wire_994;
    wire n_0533_;
    wire new_Jinkela_wire_5488;
    wire new_Jinkela_wire_6039;
    wire new_Jinkela_wire_4222;
    wire new_Jinkela_wire_1450;
    wire n_1219_;
    wire new_Jinkela_wire_85;
    wire n_1367_;
    wire new_Jinkela_wire_458;
    wire new_Jinkela_wire_5483;
    wire new_Jinkela_wire_2237;
    wire new_Jinkela_wire_6489;
    wire n_0779_;
    wire new_Jinkela_wire_4308;
    wire new_Jinkela_wire_3299;
    wire new_Jinkela_wire_183;
    wire new_Jinkela_wire_2576;
    wire new_Jinkela_wire_5914;
    wire new_Jinkela_wire_2099;
    wire n_0480_;
    wire new_Jinkela_wire_10572;
    wire new_Jinkela_wire_1334;
    wire new_Jinkela_wire_6285;
    wire new_Jinkela_wire_486;
    wire new_Jinkela_wire_2832;
    wire new_Jinkela_wire_8337;
    wire new_Jinkela_wire_5149;
    wire new_Jinkela_wire_7433;
    wire new_Jinkela_wire_3791;
    wire new_Jinkela_wire_235;
    wire new_Jinkela_wire_1988;
    wire new_Jinkela_wire_4949;
    wire new_Jinkela_wire_1057;
    wire n_0386_;
    wire new_Jinkela_wire_7288;
    wire new_Jinkela_wire_668;
    wire new_Jinkela_wire_3620;
    wire new_Jinkela_wire_5143;
    wire new_Jinkela_wire_7968;
    wire new_Jinkela_wire_6354;
    wire new_Jinkela_wire_3079;
    wire new_Jinkela_wire_6609;
    wire new_Jinkela_wire_8900;
    wire new_Jinkela_wire_8090;
    wire new_Jinkela_wire_6201;
    wire new_Jinkela_wire_5304;
    wire new_Jinkela_wire_7873;
    wire new_Jinkela_wire_9873;
    wire new_Jinkela_wire_850;
    wire new_Jinkela_wire_7221;
    wire new_Jinkela_wire_8564;
    wire new_Jinkela_wire_10179;
    wire new_Jinkela_wire_338;
    wire new_Jinkela_wire_5779;
    wire new_Jinkela_wire_3060;
    wire new_Jinkela_wire_8506;
    wire new_Jinkela_wire_5871;
    wire new_Jinkela_wire_10419;
    wire new_Jinkela_wire_1214;
    wire new_Jinkela_wire_8826;
    wire new_Jinkela_wire_5527;
    wire new_Jinkela_wire_5891;
    wire new_Jinkela_wire_6360;
    wire new_Jinkela_wire_6895;
    wire new_Jinkela_wire_9429;
    wire new_Jinkela_wire_9985;
    wire n_0465_;
    wire new_Jinkela_wire_4408;
    wire new_Jinkela_wire_10597;
    wire new_Jinkela_wire_2586;
    wire new_Jinkela_wire_3084;
    wire n_0680_;
    wire new_Jinkela_wire_3914;
    wire new_Jinkela_wire_3148;
    wire n_0673_;
    wire new_Jinkela_wire_4414;
    wire new_Jinkela_wire_1030;
    wire new_Jinkela_wire_9127;
    wire new_Jinkela_wire_1298;
    wire new_Jinkela_wire_1613;
    wire new_Jinkela_wire_3721;
    wire new_Jinkela_wire_6597;
    wire n_0435_;
    wire new_Jinkela_wire_8705;
    wire new_Jinkela_wire_2424;
    wire new_Jinkela_wire_10284;
    wire new_Jinkela_wire_1688;
    wire n_0221_;
    wire new_Jinkela_wire_1839;
    wire new_Jinkela_wire_3693;
    wire new_Jinkela_wire_9438;
    wire n_0927_;
    wire new_Jinkela_wire_7334;
    wire new_Jinkela_wire_2900;
    wire new_Jinkela_wire_2236;
    wire new_Jinkela_wire_5459;
    wire new_Jinkela_wire_7990;
    wire new_Jinkela_wire_6889;
    wire n_0200_;
    wire new_Jinkela_wire_6564;
    wire n_1139_;
    wire new_Jinkela_wire_3689;
    wire new_Jinkela_wire_4762;
    wire new_Jinkela_wire_6530;
    wire new_Jinkela_wire_5244;
    wire new_Jinkela_wire_5923;
    wire new_Jinkela_wire_3523;
    wire new_Jinkela_wire_7558;
    wire new_Jinkela_wire_8861;
    wire new_Jinkela_wire_2157;
    wire new_Jinkela_wire_157;
    wire new_Jinkela_wire_468;
    wire new_Jinkela_wire_5192;
    wire new_Jinkela_wire_6044;
    wire new_Jinkela_wire_4296;
    wire n_0773_;
    wire new_Jinkela_wire_9382;
    wire new_Jinkela_wire_6177;
    wire new_Jinkela_wire_981;
    wire n_1015_;
    wire n_0872_;
    wire new_Jinkela_wire_1458;
    wire new_Jinkela_wire_8871;
    wire new_Jinkela_wire_7863;
    wire new_Jinkela_wire_1993;
    wire n_0908_;
    wire new_Jinkela_wire_7691;
    wire new_Jinkela_wire_6108;
    wire new_Jinkela_wire_1635;
    wire new_Jinkela_wire_10416;
    wire new_Jinkela_wire_4124;
    wire new_Jinkela_wire_9487;
    wire new_Jinkela_wire_9957;
    wire new_Jinkela_wire_10382;
    wire new_Jinkela_wire_9660;
    wire new_Jinkela_wire_7317;
    wire new_Jinkela_wire_7245;
    wire n_0858_;
    wire new_Jinkela_wire_7612;
    wire new_Jinkela_wire_6094;
    wire new_Jinkela_wire_10237;
    wire n_0593_;
    wire new_Jinkela_wire_7767;
    wire new_Jinkela_wire_5601;
    wire new_Jinkela_wire_4583;
    wire n_0090_;
    wire n_1029_;
    wire new_Jinkela_wire_5551;
    wire new_Jinkela_wire_7042;
    wire new_Jinkela_wire_3248;
    wire new_Jinkela_wire_10077;
    wire n_0854_;
    wire new_Jinkela_wire_1484;
    wire new_Jinkela_wire_2150;
    wire new_Jinkela_wire_1663;
    wire new_Jinkela_wire_10630;
    wire new_Jinkela_wire_9839;
    wire new_Jinkela_wire_334;
    wire new_Jinkela_wire_464;
    wire n_0837_;
    wire new_Jinkela_wire_5410;
    wire new_Jinkela_wire_7034;
    wire new_Jinkela_wire_9742;
    wire new_Jinkela_wire_3334;
    wire n_0123_;
    wire new_Jinkela_wire_8800;
    wire new_Jinkela_wire_9884;
    wire new_Jinkela_wire_1460;
    wire new_Jinkela_wire_10549;
    wire new_Jinkela_wire_1242;
    wire new_Jinkela_wire_10436;
    wire new_Jinkela_wire_9152;
    wire new_Jinkela_wire_2328;
    wire new_Jinkela_wire_5078;
    wire new_Jinkela_wire_3204;
    wire n_1001_;
    wire new_Jinkela_wire_8924;
    wire new_Jinkela_wire_1565;
    wire n_0097_;
    wire new_Jinkela_wire_4725;
    wire new_Jinkela_wire_3363;
    wire new_Jinkela_wire_1683;
    wire new_Jinkela_wire_2135;
    wire n_1315_;
    wire n_0509_;
    wire new_Jinkela_wire_9706;
    wire new_Jinkela_wire_4591;
    wire new_Jinkela_wire_3798;
    wire n_0613_;
    wire n_1304_;
    wire new_Jinkela_wire_2472;
    wire new_Jinkela_wire_1502;
    wire new_Jinkela_wire_41;
    wire new_Jinkela_wire_3031;
    wire new_Jinkela_wire_1714;
    wire new_Jinkela_wire_8723;
    wire n_0780_;
    wire new_Jinkela_wire_8942;
    wire new_Jinkela_wire_6942;
    wire new_Jinkela_wire_9703;
    wire new_Jinkela_wire_1627;
    wire new_Jinkela_wire_2189;
    wire new_Jinkela_wire_4381;
    wire new_Jinkela_wire_9213;
    wire new_Jinkela_wire_6327;
    wire new_Jinkela_wire_3058;
    wire new_Jinkela_wire_5243;
    wire new_Jinkela_wire_3046;
    wire n_0173_;
    wire new_Jinkela_wire_3561;
    wire new_Jinkela_wire_296;
    wire n_0487_;
    wire new_Jinkela_wire_501;
    wire new_Jinkela_wire_6699;
    wire new_Jinkela_wire_9644;
    wire new_Jinkela_wire_1456;
    wire new_Jinkela_wire_3734;
    wire new_Jinkela_wire_7690;
    wire new_Jinkela_wire_10494;
    wire new_Jinkela_wire_10170;
    wire new_Jinkela_wire_3653;
    wire new_Jinkela_wire_8912;
    wire new_Jinkela_wire_7281;
    wire new_Jinkela_wire_4325;
    wire new_Jinkela_wire_5331;
    wire new_Jinkela_wire_4598;
    wire new_Jinkela_wire_9745;
    wire new_Jinkela_wire_392;
    wire new_Jinkela_wire_1452;
    wire new_Jinkela_wire_2569;
    wire n_0445_;
    wire new_Jinkela_wire_5339;
    wire new_Jinkela_wire_4678;
    wire new_Jinkela_wire_1003;
    wire new_Jinkela_wire_8038;
    wire new_Jinkela_wire_9358;
    wire new_Jinkela_wire_5790;
    wire n_1257_;
    wire n_0576_;
    wire new_Jinkela_wire_4497;
    wire new_Jinkela_wire_8742;
    wire n_0432_;
    wire new_Jinkela_wire_8055;
    wire new_Jinkela_wire_7225;
    wire new_Jinkela_wire_9891;
    wire new_Jinkela_wire_6237;
    wire new_Jinkela_wire_3141;
    wire new_Jinkela_wire_5366;
    wire new_Jinkela_wire_1004;
    wire new_Jinkela_wire_3179;
    wire new_Jinkela_wire_5443;
    wire new_Jinkela_wire_2170;
    wire n_0041_;
    wire new_Jinkela_wire_3560;
    wire new_Jinkela_wire_8135;
    wire new_Jinkela_wire_7772;
    wire new_Jinkela_wire_6553;
    wire new_Jinkela_wire_3042;
    wire new_Jinkela_wire_4112;
    wire new_Jinkela_wire_4734;
    wire new_Jinkela_wire_8632;
    wire new_Jinkela_wire_9542;
    wire new_Jinkela_wire_7264;
    wire new_Jinkela_wire_9014;
    wire new_Jinkela_wire_8557;
    wire new_Jinkela_wire_4665;
    wire new_Jinkela_wire_2888;
    wire new_Jinkela_wire_9441;
    wire new_Jinkela_wire_1693;
    wire n_1073_;
    wire new_Jinkela_wire_144;
    wire new_Jinkela_wire_1668;
    wire new_Jinkela_wire_6244;
    wire new_Jinkela_wire_3244;
    wire new_Jinkela_wire_7191;
    wire new_Jinkela_wire_3989;
    wire new_Jinkela_wire_930;
    wire new_Jinkela_wire_8138;
    wire new_Jinkela_wire_6897;
    wire n_0949_;
    wire new_Jinkela_wire_5927;
    wire new_Jinkela_wire_7512;
    wire new_Jinkela_wire_5731;
    wire new_Jinkela_wire_2244;
    wire new_Jinkela_wire_3257;
    wire new_Jinkela_wire_5382;
    wire new_Jinkela_wire_2957;
    wire new_Jinkela_wire_6440;
    wire new_Jinkela_wire_9301;
    wire new_Jinkela_wire_7897;
    wire new_Jinkela_wire_1284;
    wire new_Jinkela_wire_6837;
    wire new_Jinkela_wire_2649;
    wire new_Jinkela_wire_3857;
    wire n_0491_;
    wire new_Jinkela_wire_3955;
    wire new_Jinkela_wire_3151;
    wire n_0496_;
    wire n_1319_;
    wire new_Jinkela_wire_598;
    wire new_Jinkela_wire_4430;
    wire new_Jinkela_wire_8380;
    wire n_1130_;
    wire new_Jinkela_wire_8804;
    wire new_Jinkela_wire_5163;
    wire new_Jinkela_wire_3853;
    wire new_Jinkela_wire_5637;
    wire new_Jinkela_wire_1494;
    wire new_Jinkela_wire_4186;
    wire new_Jinkela_wire_3552;
    wire n_0048_;
    wire new_Jinkela_wire_9977;
    wire new_Jinkela_wire_10210;
    wire new_Jinkela_wire_10358;
    wire n_0860_;
    wire new_Jinkela_wire_9284;
    wire n_0212_;
    wire new_Jinkela_wire_6787;
    wire new_Jinkela_wire_3785;
    wire n_1320_;
    wire new_Jinkela_wire_6378;
    wire n_1225_;
    wire new_Jinkela_wire_879;
    wire new_Jinkela_wire_5878;
    wire new_Jinkela_wire_816;
    wire n_0363_;
    wire new_Jinkela_wire_588;
    wire new_Jinkela_wire_10031;
    wire n_1112_;
    wire new_Jinkela_wire_1230;
    wire new_Jinkela_wire_6985;
    wire new_Jinkela_wire_7330;
    wire new_Jinkela_wire_8626;
    wire n_0133_;
    wire n_1279_;
    wire new_Jinkela_wire_2000;
    wire new_Jinkela_wire_5547;
    wire new_Jinkela_wire_5238;
    wire new_Jinkela_wire_7490;
    wire new_Jinkela_wire_6138;
    wire new_Jinkela_wire_4346;
    wire new_Jinkela_wire_2069;
    wire new_Jinkela_wire_6454;
    wire new_Jinkela_wire_6784;
    wire new_Jinkela_wire_3710;
    wire new_Jinkela_wire_8343;
    wire new_Jinkela_wire_3581;
    wire n_0632_;
    wire new_Jinkela_wire_7992;
    wire new_Jinkela_wire_5476;
    wire n_0380_;
    wire n_0130_;
    wire new_Jinkela_wire_6674;
    wire new_Jinkela_wire_8778;
    wire new_Jinkela_wire_4053;
    wire n_0741_;
    wire new_Jinkela_wire_9195;
    wire new_Jinkela_wire_2257;
    wire new_Jinkela_wire_2901;
    wire new_Jinkela_wire_7341;
    wire new_Jinkela_wire_7966;
    wire new_Jinkela_wire_3398;
    wire n_0467_;
    wire new_Jinkela_wire_9591;
    wire new_Jinkela_wire_1995;
    wire new_Jinkela_wire_8940;
    wire new_Jinkela_wire_1080;
    wire new_Jinkela_wire_6753;
    wire new_Jinkela_wire_2487;
    wire new_Jinkela_wire_460;
    wire new_Jinkela_wire_7419;
    wire new_Jinkela_wire_5892;
    wire new_Jinkela_wire_5426;
    wire new_Jinkela_wire_9902;
    wire new_Jinkela_wire_559;
    wire new_Jinkela_wire_5107;
    wire new_Jinkela_wire_8877;
    wire new_Jinkela_wire_5584;
    wire new_Jinkela_wire_5817;
    wire new_Jinkela_wire_5628;
    wire new_Jinkela_wire_9486;
    wire new_Jinkela_wire_7871;
    wire new_Jinkela_wire_2242;
    wire new_Jinkela_wire_7845;
    wire new_Jinkela_wire_2097;
    wire new_Jinkela_wire_572;
    wire new_Jinkela_wire_5320;
    wire new_Jinkela_wire_10204;
    wire new_Jinkela_wire_8977;
    wire new_Jinkela_wire_4466;
    wire new_Jinkela_wire_8909;
    wire new_Jinkela_wire_827;
    wire new_Jinkela_wire_7919;
    wire new_Jinkela_wire_5215;
    wire new_Jinkela_wire_2607;
    wire new_Jinkela_wire_10298;
    wire new_Jinkela_wire_6915;
    wire new_Jinkela_wire_9498;
    wire new_Jinkela_wire_653;
    wire n_0060_;
    wire new_Jinkela_wire_10552;
    wire new_Jinkela_wire_7482;
    wire new_Jinkela_wire_3973;
    wire n_1259_;
    wire new_Jinkela_wire_10165;
    wire new_Jinkela_wire_613;
    wire new_Jinkela_wire_7448;
    wire n_0359_;
    wire new_Jinkela_wire_5806;
    wire n_0416_;
    wire new_Jinkela_wire_4680;
    wire new_Jinkela_wire_4411;
    wire new_net_4;
    wire new_Jinkela_wire_9651;
    wire new_Jinkela_wire_1098;
    wire new_Jinkela_wire_2027;
    wire new_Jinkela_wire_5070;
    wire n_0140_;
    wire new_Jinkela_wire_270;
    wire new_Jinkela_wire_2200;
    wire new_Jinkela_wire_9518;
    wire new_Jinkela_wire_5141;
    wire new_Jinkela_wire_10155;
    wire new_Jinkela_wire_10066;
    wire new_Jinkela_wire_5438;
    wire new_net_2499;
    wire new_Jinkela_wire_3811;
    wire new_Jinkela_wire_4631;
    wire new_Jinkela_wire_9264;
    wire new_Jinkela_wire_5011;
    wire new_Jinkela_wire_3002;
    wire new_Jinkela_wire_4724;
    wire new_Jinkela_wire_8031;
    wire n_1240_;
    wire new_Jinkela_wire_6213;
    wire new_Jinkela_wire_1615;
    wire n_0802_;
    wire new_Jinkela_wire_9752;
    wire new_Jinkela_wire_8996;
    wire new_Jinkela_wire_5730;
    wire n_1280_;
    wire new_Jinkela_wire_8164;
    wire new_Jinkela_wire_9415;
    wire new_Jinkela_wire_4109;
    wire new_Jinkela_wire_4373;
    wire n_1013_;
    wire new_Jinkela_wire_10460;
    wire new_Jinkela_wire_7298;
    wire new_Jinkela_wire_4869;
    wire new_Jinkela_wire_608;
    wire new_Jinkela_wire_1153;
    wire new_Jinkela_wire_4020;
    wire new_Jinkela_wire_3170;
    wire new_Jinkela_wire_7702;
    wire new_Jinkela_wire_8576;
    wire new_Jinkela_wire_3986;
    wire n_0629_;
    wire new_Jinkela_wire_10588;
    wire new_Jinkela_wire_8365;
    wire new_Jinkela_wire_8446;
    wire new_Jinkela_wire_8938;
    wire new_Jinkela_wire_4927;
    wire new_Jinkela_wire_2020;
    wire new_Jinkela_wire_3068;
    wire n_0036_;
    wire new_Jinkela_wire_9256;
    wire new_Jinkela_wire_6725;
    wire new_Jinkela_wire_9232;
    wire new_Jinkela_wire_10614;
    wire new_Jinkela_wire_3430;
    wire new_Jinkela_wire_3451;
    wire new_Jinkela_wire_1087;
    wire new_Jinkela_wire_2843;
    wire new_Jinkela_wire_3238;
    wire n_0267_;
    wire new_Jinkela_wire_4159;
    wire new_Jinkela_wire_4271;
    wire new_Jinkela_wire_3372;
    wire new_Jinkela_wire_3333;
    wire new_Jinkela_wire_240;
    wire new_Jinkela_wire_7817;
    wire new_Jinkela_wire_8341;
    wire n_1091_;
    wire new_Jinkela_wire_9268;
    wire new_Jinkela_wire_3761;
    wire new_Jinkela_wire_946;
    wire new_Jinkela_wire_6527;
    wire new_Jinkela_wire_381;
    wire n_0641_;
    wire new_Jinkela_wire_4333;
    wire new_Jinkela_wire_10590;
    wire new_Jinkela_wire_159;
    wire new_Jinkela_wire_9464;
    wire new_Jinkela_wire_7037;
    wire new_Jinkela_wire_7720;
    wire new_Jinkela_wire_6056;
    wire n_0848_;
    wire new_Jinkela_wire_9254;
    wire new_Jinkela_wire_2191;
    wire new_Jinkela_wire_6095;
    wire new_Jinkela_wire_1670;
    wire n_0506_;
    wire new_Jinkela_wire_5391;
    wire new_Jinkela_wire_10306;
    wire new_Jinkela_wire_4624;
    wire new_Jinkela_wire_5523;
    wire new_Jinkela_wire_5813;
    wire new_Jinkela_wire_5012;
    wire new_Jinkela_wire_9123;
    wire new_Jinkela_wire_615;
    wire new_Jinkela_wire_7393;
    wire new_Jinkela_wire_2252;
    wire new_Jinkela_wire_8894;
    wire new_Jinkela_wire_9128;
    wire new_Jinkela_wire_8497;
    wire new_Jinkela_wire_7385;
    wire new_Jinkela_wire_155;
    wire new_Jinkela_wire_6932;
    wire new_Jinkela_wire_2964;
    wire new_Jinkela_wire_5494;
    wire new_Jinkela_wire_6857;
    wire new_Jinkela_wire_8461;
    wire new_Jinkela_wire_3824;
    wire new_Jinkela_wire_4634;
    wire new_Jinkela_wire_1120;
    wire new_Jinkela_wire_1906;
    wire new_Jinkela_wire_3255;
    wire new_Jinkela_wire_3648;
    wire new_Jinkela_wire_6036;
    wire new_Jinkela_wire_9505;
    wire new_Jinkela_wire_4344;
    wire new_Jinkela_wire_4095;
    wire new_Jinkela_wire_7631;
    wire new_Jinkela_wire_3514;
    wire new_Jinkela_wire_3717;
    wire new_Jinkela_wire_2042;
    wire new_Jinkela_wire_8586;
    wire new_Jinkela_wire_2024;
    wire new_Jinkela_wire_4676;
    wire new_Jinkela_wire_2687;
    wire n_1323_;
    wire new_Jinkela_wire_3510;
    wire new_Jinkela_wire_8664;
    wire new_Jinkela_wire_3718;
    wire new_Jinkela_wire_9368;
    wire new_Jinkela_wire_10043;
    wire new_Jinkela_wire_471;
    wire new_Jinkela_wire_728;
    wire new_Jinkela_wire_1944;
    wire new_Jinkela_wire_4376;
    wire new_Jinkela_wire_8648;
    wire new_Jinkela_wire_3500;
    wire new_Jinkela_wire_6654;
    wire n_0102_;
    wire new_net_3;
    wire new_Jinkela_wire_782;
    wire n_0763_;
    wire new_Jinkela_wire_3232;
    wire new_Jinkela_wire_7805;
    wire new_Jinkela_wire_1161;
    wire new_Jinkela_wire_2213;
    wire new_Jinkela_wire_8661;
    wire n_0603_;
    wire n_1056_;
    wire new_Jinkela_wire_134;
    wire n_0150_;
    wire new_Jinkela_wire_7041;
    wire new_Jinkela_wire_7546;
    wire new_Jinkela_wire_4643;
    wire new_Jinkela_wire_4387;
    wire new_Jinkela_wire_10010;
    wire new_Jinkela_wire_6580;
    wire new_Jinkela_wire_391;
    wire new_Jinkela_wire_6636;
    wire new_Jinkela_wire_4984;
    wire new_Jinkela_wire_7717;
    wire new_Jinkela_wire_7920;
    wire new_Jinkela_wire_5792;
    wire new_Jinkela_wire_6935;
    wire new_Jinkela_wire_7492;
    wire new_Jinkela_wire_8767;
    wire new_Jinkela_wire_6734;
    wire n_0948_;
    wire new_Jinkela_wire_2833;
    wire new_Jinkela_wire_8220;
    wire new_Jinkela_wire_3464;
    wire new_Jinkela_wire_6875;
    wire new_Jinkela_wire_5752;
    wire new_Jinkela_wire_9417;
    wire new_Jinkela_wire_4237;
    wire new_Jinkela_wire_10116;
    wire new_Jinkela_wire_10480;
    wire new_Jinkela_wire_5213;
    wire new_Jinkela_wire_161;
    wire new_Jinkela_wire_754;
    wire new_Jinkela_wire_6644;
    wire new_Jinkela_wire_2716;
    wire n_1111_;
    wire new_Jinkela_wire_8546;
    wire new_Jinkela_wire_10164;
    wire new_Jinkela_wire_9196;
    wire new_Jinkela_wire_5609;
    wire new_Jinkela_wire_2625;
    wire new_Jinkela_wire_10294;
    wire new_Jinkela_wire_585;
    wire n_0864_;
    wire new_Jinkela_wire_2168;
    wire new_Jinkela_wire_10195;
    wire new_Jinkela_wire_8434;
    wire new_Jinkela_wire_5689;
    wire new_Jinkela_wire_8627;
    wire new_Jinkela_wire_4823;
    wire new_Jinkela_wire_7500;
    wire new_Jinkela_wire_5035;
    wire n_1061_;
    wire new_Jinkela_wire_960;
    wire new_Jinkela_wire_2235;
    wire new_Jinkela_wire_9888;
    wire new_Jinkela_wire_8842;
    wire new_Jinkela_wire_360;
    wire new_net_2;
    wire new_Jinkela_wire_6780;
    wire new_Jinkela_wire_4718;
    wire new_Jinkela_wire_198;
    wire new_Jinkela_wire_2878;
    wire new_Jinkela_wire_9815;
    wire new_Jinkela_wire_4772;
    wire n_0661_;
    wire new_Jinkela_wire_10385;
    wire new_net_6;
    wire new_Jinkela_wire_7426;
    wire new_Jinkela_wire_9712;
    wire new_Jinkela_wire_8400;
    wire new_Jinkela_wire_7149;
    wire n_0470_;
    wire new_Jinkela_wire_6514;
    wire new_Jinkela_wire_10576;
    wire new_Jinkela_wire_1665;
    wire new_Jinkela_wire_9526;
    wire new_Jinkela_wire_4815;
    wire new_Jinkela_wire_273;
    wire new_Jinkela_wire_5995;
    wire new_Jinkela_wire_6008;
    wire new_Jinkela_wire_10450;
    wire new_Jinkela_wire_1136;
    wire new_Jinkela_wire_7219;
    wire new_Jinkela_wire_3458;
    wire new_Jinkela_wire_3308;
    wire new_Jinkela_wire_6903;
    wire new_Jinkela_wire_7983;
    wire new_Jinkela_wire_9328;
    wire new_Jinkela_wire_3826;
    wire n_0586_;
    wire new_Jinkela_wire_7432;
    wire new_Jinkela_wire_6425;
    wire new_Jinkela_wire_94;
    wire new_Jinkela_wire_8674;
    wire new_Jinkela_wire_10440;
    wire new_Jinkela_wire_10351;
    wire new_Jinkela_wire_4125;
    wire new_Jinkela_wire_4659;
    wire new_Jinkela_wire_2434;
    wire new_Jinkela_wire_2821;
    wire n_1200_;
    wire new_Jinkela_wire_7616;
    wire new_Jinkela_wire_4711;
    wire new_Jinkela_wire_1253;
    wire new_Jinkela_wire_193;
    wire new_Jinkela_wire_8578;
    wire new_Jinkela_wire_6735;
    wire new_Jinkela_wire_1902;
    wire new_Jinkela_wire_3941;
    wire new_Jinkela_wire_8344;
    wire new_Jinkela_wire_1191;
    wire new_Jinkela_wire_5533;
    wire new_Jinkela_wire_1470;
    wire new_Jinkela_wire_10030;
    wire new_Jinkela_wire_6715;
    wire new_Jinkela_wire_1986;
    wire new_Jinkela_wire_3491;
    wire new_Jinkela_wire_1281;
    wire new_Jinkela_wire_2761;
    wire new_Jinkela_wire_4890;
    wire new_Jinkela_wire_2521;
    wire new_Jinkela_wire_546;
    wire new_Jinkela_wire_7484;
    wire new_Jinkela_wire_6551;
    wire new_Jinkela_wire_3327;
    wire n_0952_;
    wire new_Jinkela_wire_5907;
    wire new_Jinkela_wire_136;
    wire new_Jinkela_wire_1967;
    wire new_Jinkela_wire_10525;
    wire new_Jinkela_wire_9308;
    wire new_Jinkela_wire_3866;
    wire new_Jinkela_wire_7562;
    wire new_Jinkela_wire_4933;
    wire new_Jinkela_wire_8766;
    wire new_Jinkela_wire_69;
    wire new_Jinkela_wire_5112;
    wire new_Jinkela_wire_1629;
    wire new_Jinkela_wire_9773;
    wire new_net_2517;
    wire new_Jinkela_wire_5240;
    wire new_Jinkela_wire_1579;
    wire new_Jinkela_wire_5478;
    wire new_Jinkela_wire_6068;
    wire new_Jinkela_wire_2351;
    wire new_Jinkela_wire_6230;
    wire new_Jinkela_wire_6321;
    wire n_1074_;
    wire new_Jinkela_wire_132;
    wire new_Jinkela_wire_9108;
    wire new_Jinkela_wire_3716;
    wire new_Jinkela_wire_8334;
    wire new_Jinkela_wire_1419;
    wire new_Jinkela_wire_1290;
    wire new_Jinkela_wire_372;
    wire new_Jinkela_wire_5284;
    wire new_Jinkela_wire_3434;
    wire new_Jinkela_wire_7246;
    wire new_Jinkela_wire_9895;
    wire new_Jinkela_wire_7633;
    wire new_Jinkela_wire_10406;
    wire new_Jinkela_wire_6957;
    wire new_Jinkela_wire_7991;
    wire new_Jinkela_wire_7087;
    wire new_Jinkela_wire_8026;
    wire new_Jinkela_wire_9913;
    wire new_Jinkela_wire_10086;
    wire new_Jinkela_wire_5081;
    wire new_Jinkela_wire_9613;
    wire new_Jinkela_wire_3099;
    wire new_Jinkela_wire_1975;
    wire n_0823_;
    wire n_0857_;
    wire n_0395_;
    wire new_Jinkela_wire_10528;
    wire new_Jinkela_wire_5294;
    wire new_Jinkela_wire_10557;
    wire new_Jinkela_wire_9349;
    wire new_Jinkela_wire_3911;
    wire new_Jinkela_wire_9534;
    wire new_Jinkela_wire_5390;
    wire new_Jinkela_wire_1122;
    wire n_0098_;
    wire new_Jinkela_wire_7174;
    wire new_Jinkela_wire_8549;
    wire new_Jinkela_wire_8473;
    wire new_Jinkela_wire_5363;
    wire n_0527_;
    wire new_Jinkela_wire_6619;
    wire new_Jinkela_wire_576;
    wire new_Jinkela_wire_7311;
    wire new_Jinkela_wire_8700;
    wire new_Jinkela_wire_6885;
    wire new_Jinkela_wire_823;
    wire new_Jinkela_wire_8973;
    wire new_Jinkela_wire_7257;
    wire new_Jinkela_wire_2609;
    wire new_Jinkela_wire_9576;
    wire new_Jinkela_wire_2385;
    wire new_Jinkela_wire_6382;
    wire new_Jinkela_wire_9304;
    wire new_Jinkela_wire_1661;
    wire new_Jinkela_wire_7947;
    wire new_Jinkela_wire_3482;
    wire new_Jinkela_wire_4522;
    wire new_Jinkela_wire_6603;
    wire new_Jinkela_wire_1033;
    wire new_Jinkela_wire_10368;
    wire new_Jinkela_wire_1878;
    wire n_0817_;
    wire new_Jinkela_wire_10172;
    wire new_Jinkela_wire_10127;
    wire new_Jinkela_wire_9194;
    wire new_Jinkela_wire_8149;
    wire new_Jinkela_wire_6180;
    wire new_Jinkela_wire_4087;
    wire new_Jinkela_wire_2066;
    wire new_Jinkela_wire_1658;
    wire new_Jinkela_wire_3960;
    wire new_Jinkela_wire_3528;
    wire new_Jinkela_wire_1052;
    wire new_Jinkela_wire_8005;
    wire new_Jinkela_wire_5994;
    wire n_0619_;
    wire new_Jinkela_wire_9042;
    wire new_Jinkela_wire_3094;
    wire new_Jinkela_wire_9887;
    wire new_Jinkela_wire_4263;
    wire new_Jinkela_wire_10239;
    wire new_Jinkela_wire_8102;
    wire new_Jinkela_wire_5464;
    wire new_Jinkela_wire_4386;
    wire new_Jinkela_wire_8074;
    wire new_Jinkela_wire_4078;
    wire new_Jinkela_wire_2485;
    wire new_Jinkela_wire_5268;
    wire new_Jinkela_wire_7937;
    wire new_Jinkela_wire_7928;
    wire new_Jinkela_wire_275;
    wire new_Jinkela_wire_1157;
    wire new_Jinkela_wire_2848;
    wire new_Jinkela_wire_3163;
    wire new_Jinkela_wire_3321;
    wire new_Jinkela_wire_430;
    wire new_Jinkela_wire_5895;
    wire new_Jinkela_wire_1994;
    wire n_1027_;
    wire new_Jinkela_wire_8487;
    wire new_Jinkela_wire_8743;
    wire new_Jinkela_wire_4695;
    wire new_Jinkela_wire_5837;
    wire new_Jinkela_wire_7793;
    wire n_0224_;
    wire new_Jinkela_wire_7794;
    wire new_Jinkela_wire_702;
    wire n_1192_;
    wire new_Jinkela_wire_6646;
    wire new_Jinkela_wire_351;
    wire new_Jinkela_wire_3983;
    wire new_Jinkela_wire_6688;
    wire new_Jinkela_wire_4031;
    wire new_Jinkela_wire_4490;
    wire new_Jinkela_wire_3379;
    wire new_Jinkela_wire_5946;
    wire n_0020_;
    wire n_0755_;
    wire n_0187_;
    wire new_Jinkela_wire_922;
    wire new_Jinkela_wire_4746;
    wire new_Jinkela_wire_3211;
    wire new_Jinkela_wire_1675;
    wire new_Jinkela_wire_5913;
    wire new_Jinkela_wire_942;
    wire new_Jinkela_wire_982;
    wire new_Jinkela_wire_3593;
    wire new_Jinkela_wire_8043;
    wire new_Jinkela_wire_6051;
    wire new_Jinkela_wire_1471;
    wire new_Jinkela_wire_5223;
    wire new_Jinkela_wire_6436;
    wire new_Jinkela_wire_10521;
    wire new_Jinkela_wire_8251;
    wire new_Jinkela_wire_3074;
    wire new_Jinkela_wire_1860;
    wire new_Jinkela_wire_8125;
    wire new_Jinkela_wire_7306;
    wire new_Jinkela_wire_4554;
    wire new_Jinkela_wire_6724;
    wire new_Jinkela_wire_8458;
    wire new_Jinkela_wire_5511;
    wire new_Jinkela_wire_7713;
    wire new_Jinkela_wire_9623;
    wire new_Jinkela_wire_5955;
    wire new_Jinkela_wire_1111;
    wire new_Jinkela_wire_1288;
    wire new_Jinkela_wire_2934;
    wire new_Jinkela_wire_2243;
    wire new_Jinkela_wire_5867;
    wire new_Jinkela_wire_2839;
    wire new_Jinkela_wire_5134;
    wire new_Jinkela_wire_10384;
    wire new_Jinkela_wire_6196;
    wire new_Jinkela_wire_77;
    wire new_Jinkela_wire_9532;
    wire new_Jinkela_wire_1761;
    wire new_Jinkela_wire_10110;
    wire new_Jinkela_wire_3609;
    wire new_Jinkela_wire_2556;
    wire new_Jinkela_wire_2762;
    wire new_Jinkela_wire_5591;
    wire new_Jinkela_wire_5017;
    wire new_Jinkela_wire_7729;
    wire n_0720_;
    wire new_Jinkela_wire_258;
    wire new_Jinkela_wire_9511;
    wire n_1316_;
    wire new_Jinkela_wire_7964;
    wire new_Jinkela_wire_3764;
    wire new_Jinkela_wire_8247;
    wire new_Jinkela_wire_106;
    wire new_Jinkela_wire_8071;
    wire new_Jinkela_wire_5406;
    wire new_Jinkela_wire_7645;
    wire new_Jinkela_wire_7110;
    wire new_Jinkela_wire_6373;
    wire new_Jinkela_wire_8615;
    wire new_Jinkela_wire_1231;
    wire new_Jinkela_wire_3725;
    wire new_Jinkela_wire_7807;
    wire new_Jinkela_wire_1479;
    wire new_Jinkela_wire_5940;
    wire new_Jinkela_wire_10026;
    wire n_0067_;
    wire new_Jinkela_wire_6063;
    wire new_Jinkela_wire_4326;
    wire new_Jinkela_wire_2990;
    wire new_Jinkela_wire_9946;
    wire new_Jinkela_wire_3276;
    wire new_Jinkela_wire_636;
    wire new_Jinkela_wire_5233;
    wire new_Jinkela_wire_3934;
    wire new_Jinkela_wire_9164;
    wire new_Jinkela_wire_4573;
    wire new_Jinkela_wire_789;
    wire new_Jinkela_wire_897;
    wire new_Jinkela_wire_2026;
    wire new_Jinkela_wire_1720;
    wire new_Jinkela_wire_10499;
    wire new_Jinkela_wire_4622;
    wire new_Jinkela_wire_5900;
    wire new_Jinkela_wire_3703;
    wire new_Jinkela_wire_4055;
    wire new_Jinkela_wire_1989;
    wire new_Jinkela_wire_9077;
    wire n_0955_;
    wire new_Jinkela_wire_7922;
    wire new_Jinkela_wire_2680;
    wire new_Jinkela_wire_5824;
    wire new_Jinkela_wire_10230;
    wire new_Jinkela_wire_1828;
    wire new_Jinkela_wire_5222;
    wire new_Jinkela_wire_8287;
    wire new_Jinkela_wire_9971;
    wire n_0984_;
    wire new_Jinkela_wire_10215;
    wire new_Jinkela_wire_532;
    wire new_Jinkela_wire_4889;
    wire new_Jinkela_wire_9547;
    wire new_Jinkela_wire_5862;
    wire new_Jinkela_wire_3202;
    wire new_Jinkela_wire_9088;
    wire n_0651_;
    wire new_Jinkela_wire_5959;
    wire new_Jinkela_wire_1;
    wire new_Jinkela_wire_4484;
    wire new_Jinkela_wire_6928;
    wire new_Jinkela_wire_1010;
    wire new_Jinkela_wire_6770;
    wire new_Jinkela_wire_2058;
    wire new_Jinkela_wire_6061;
    wire new_Jinkela_wire_1133;
    wire new_Jinkela_wire_1254;
    wire new_Jinkela_wire_8182;
    wire new_Jinkela_wire_5803;
    wire new_Jinkela_wire_405;
    wire new_Jinkela_wire_7745;
    wire new_Jinkela_wire_2176;
    wire new_Jinkela_wire_6251;
    wire new_Jinkela_wire_5843;
    wire new_Jinkela_wire_8210;
    wire new_Jinkela_wire_9005;
    wire new_Jinkela_wire_346;
    wire n_1260_;
    wire new_Jinkela_wire_10608;
    wire new_Jinkela_wire_239;
    wire new_Jinkela_wire_1382;
    wire new_Jinkela_wire_6214;
    wire new_Jinkela_wire_10496;
    wire new_Jinkela_wire_9595;
    wire new_Jinkela_wire_3306;
    wire new_Jinkela_wire_9139;
    wire new_Jinkela_wire_3888;
    wire new_Jinkela_wire_328;
    wire new_Jinkela_wire_5085;
    wire new_Jinkela_wire_3583;
    wire new_Jinkela_wire_119;
    wire new_Jinkela_wire_1576;
    wire new_Jinkela_wire_2374;
    wire new_Jinkela_wire_4313;
    wire new_Jinkela_wire_9058;
    wire new_Jinkela_wire_1908;
    wire new_Jinkela_wire_148;
    wire new_Jinkela_wire_8666;
    wire new_Jinkela_wire_1550;
    wire new_Jinkela_wire_8830;
    wire n_0028_;
    wire new_Jinkela_wire_195;
    wire new_Jinkela_wire_7986;
    wire n_0381_;
    wire new_Jinkela_wire_10318;
    wire new_Jinkela_wire_10052;
    wire new_Jinkela_wire_3152;
    wire new_Jinkela_wire_1963;
    wire n_0047_;
    wire new_Jinkela_wire_3640;
    wire new_Jinkela_wire_2810;
    wire new_Jinkela_wire_2530;
    wire new_Jinkela_wire_2513;
    wire n_0412_;
    wire n_1250_;
    wire new_Jinkela_wire_6587;
    wire new_Jinkela_wire_91;
    wire new_Jinkela_wire_2837;
    wire new_Jinkela_wire_5288;
    wire new_Jinkela_wire_7336;
    wire new_Jinkela_wire_737;
    wire new_Jinkela_wire_8237;
    wire new_Jinkela_wire_2785;
    wire new_Jinkela_wire_6532;
    wire new_Jinkela_wire_7733;
    wire new_Jinkela_wire_2230;
    wire new_Jinkela_wire_7957;
    wire new_Jinkela_wire_6112;
    wire new_Jinkela_wire_2376;
    wire new_Jinkela_wire_10338;
    wire new_Jinkela_wire_2483;
    wire new_Jinkela_wire_1875;
    wire new_Jinkela_wire_3606;
    wire new_Jinkela_wire_2452;
    wire new_Jinkela_wire_6303;
    wire new_Jinkela_wire_9282;
    wire new_Jinkela_wire_656;
    wire new_Jinkela_wire_3615;
    wire new_Jinkela_wire_1945;
    wire new_Jinkela_wire_3362;
    wire new_Jinkela_wire_9622;
    wire new_Jinkela_wire_1853;
    wire new_Jinkela_wire_10042;
    wire new_Jinkela_wire_2633;
    wire new_Jinkela_wire_3694;
    wire new_Jinkela_wire_9003;
    wire new_net_2493;
    wire new_Jinkela_wire_4403;
    wire new_Jinkela_wire_1431;
    wire new_Jinkela_wire_2303;
    wire new_Jinkela_wire_5783;
    wire n_0286_;
    wire new_Jinkela_wire_1255;
    wire new_Jinkela_wire_3147;
    wire new_Jinkela_wire_5883;
    wire new_Jinkela_wire_6671;
    wire new_Jinkela_wire_5945;
    wire new_Jinkela_wire_2819;
    wire new_Jinkela_wire_2055;
    wire new_Jinkela_wire_8584;
    wire n_0882_;
    wire new_Jinkela_wire_10037;
    wire new_Jinkela_wire_5358;
    wire new_Jinkela_wire_3695;
    wire new_Jinkela_wire_222;
    wire new_Jinkela_wire_10335;
    wire new_Jinkela_wire_8035;
    wire new_Jinkela_wire_6668;
    wire new_Jinkela_wire_5289;
    wire new_Jinkela_wire_9313;
    wire new_Jinkela_wire_2404;
    wire new_Jinkela_wire_4184;
    wire new_Jinkela_wire_4824;
    wire n_0338_;
    wire new_Jinkela_wire_2713;
    wire new_Jinkela_wire_2126;
    wire new_Jinkela_wire_9846;
    wire n_0766_;
    wire new_Jinkela_wire_3587;
    wire new_Jinkela_wire_9249;
    wire new_Jinkela_wire_5132;
    wire new_Jinkela_wire_1328;
    wire new_Jinkela_wire_10479;
    wire new_Jinkela_wire_2197;
    wire new_Jinkela_wire_3040;
    wire new_Jinkela_wire_4540;
    wire new_Jinkela_wire_744;
    wire new_Jinkela_wire_1537;
    wire new_Jinkela_wire_587;
    wire new_Jinkela_wire_10258;
    wire new_Jinkela_wire_5756;
    wire new_Jinkela_wire_3388;
    wire new_net_2505;
    wire new_Jinkela_wire_9615;
    wire new_Jinkela_wire_9959;
    wire new_Jinkela_wire_4799;
    wire new_Jinkela_wire_699;
    wire new_Jinkela_wire_6190;
    wire n_1368_;
    wire new_Jinkela_wire_9791;
    wire new_Jinkela_wire_5224;
    wire new_Jinkela_wire_9433;
    wire new_Jinkela_wire_1970;
    wire new_Jinkela_wire_5688;
    wire new_Jinkela_wire_2896;
    wire new_Jinkela_wire_3320;
    wire new_Jinkela_wire_3006;
    wire new_Jinkela_wire_547;
    wire new_Jinkela_wire_7925;
    wire new_Jinkela_wire_4158;
    wire new_Jinkela_wire_10483;
    wire new_Jinkela_wire_2493;
    wire new_Jinkela_wire_5715;
    wire new_Jinkela_wire_4794;
    wire new_Jinkela_wire_7014;
    wire new_Jinkela_wire_6077;
    wire new_Jinkela_wire_8086;
    wire new_Jinkela_wire_935;
    wire new_Jinkela_wire_2666;
    wire new_Jinkela_wire_1078;
    wire new_Jinkela_wire_691;
    wire new_Jinkela_wire_7657;
    wire new_Jinkela_wire_516;
    wire new_Jinkela_wire_7395;
    wire new_Jinkela_wire_3486;
    wire new_Jinkela_wire_6097;
    wire new_Jinkela_wire_5864;
    wire new_Jinkela_wire_1921;
    wire new_Jinkela_wire_4257;
    wire new_Jinkela_wire_1671;
    wire new_Jinkela_wire_9351;
    wire new_Jinkela_wire_772;
    wire new_Jinkela_wire_4771;
    wire new_Jinkela_wire_9923;
    wire new_Jinkela_wire_5452;
    wire new_Jinkela_wire_6655;
    wire new_Jinkela_wire_2233;
    wire new_Jinkela_wire_4113;
    wire new_Jinkela_wire_525;
    wire new_Jinkela_wire_138;
    wire new_Jinkela_wire_2624;
    wire new_Jinkela_wire_4340;
    wire new_Jinkela_wire_5619;
    wire new_Jinkela_wire_7848;
    wire new_Jinkela_wire_8440;
    wire new_Jinkela_wire_7234;
    wire new_Jinkela_wire_110;
    wire new_Jinkela_wire_1574;
    wire new_Jinkela_wire_9715;
    wire new_Jinkela_wire_1115;
    wire new_Jinkela_wire_7187;
    wire new_Jinkela_wire_3097;
    wire new_Jinkela_wire_6236;
    wire new_Jinkela_wire_10536;
    wire new_Jinkela_wire_5700;
    wire new_Jinkela_wire_6405;
    wire new_Jinkela_wire_9063;
    wire new_Jinkela_wire_2344;
    wire new_Jinkela_wire_2542;
    wire new_Jinkela_wire_8959;
    wire new_Jinkela_wire_5692;
    wire new_Jinkela_wire_225;
    wire new_Jinkela_wire_7310;
    wire new_Jinkela_wire_1735;
    wire new_Jinkela_wire_6959;
    wire new_Jinkela_wire_5695;
    wire new_Jinkela_wire_7240;
    wire n_1264_;
    wire new_Jinkela_wire_6250;
    wire n_0704_;
    wire new_Jinkela_wire_7459;
    wire new_Jinkela_wire_477;
    wire new_Jinkela_wire_10231;
    wire new_Jinkela_wire_6412;
    wire new_Jinkela_wire_10065;
    wire new_Jinkela_wire_8474;
    wire new_Jinkela_wire_7860;
    wire new_Jinkela_wire_3283;
    wire new_Jinkela_wire_9449;
    wire n_0843_;
    wire new_Jinkela_wire_219;
    wire new_Jinkela_wire_4048;
    wire new_Jinkela_wire_3051;
    wire new_Jinkela_wire_7359;
    wire new_Jinkela_wire_3468;
    wire new_Jinkela_wire_2752;
    wire new_Jinkela_wire_4192;
    wire n_1165_;
    wire new_Jinkela_wire_2142;
    wire new_Jinkela_wire_4538;
    wire new_Jinkela_wire_5739;
    wire new_Jinkela_wire_6626;
    wire new_Jinkela_wire_418;
    wire new_Jinkela_wire_1488;
    wire new_Jinkela_wire_5826;
    wire new_Jinkela_wire_2446;
    wire new_Jinkela_wire_8194;
    wire n_1310_;
    wire new_Jinkela_wire_176;
    wire new_Jinkela_wire_8371;
    wire new_Jinkela_wire_371;
    wire new_Jinkela_wire_7797;
    wire new_Jinkela_wire_2248;
    wire n_0369_;
    wire n_0578_;
    wire new_Jinkela_wire_2229;
    wire new_Jinkela_wire_3933;
    wire new_Jinkela_wire_3723;
    wire new_Jinkela_wire_1032;
    wire new_Jinkela_wire_8753;
    wire new_Jinkela_wire_771;
    wire new_Jinkela_wire_9698;
    wire new_Jinkela_wire_5639;
    wire n_1230_;
    wire new_Jinkela_wire_9818;
    wire new_Jinkela_wire_2941;
    wire new_Jinkela_wire_5019;
    wire new_Jinkela_wire_8620;
    wire new_Jinkela_wire_6179;
    wire new_Jinkela_wire_10162;
    wire new_Jinkela_wire_9747;
    wire n_0915_;
    wire new_Jinkela_wire_7142;
    wire new_Jinkela_wire_9669;
    wire new_Jinkela_wire_5068;
    wire new_Jinkela_wire_8883;
    wire n_1213_;
    wire new_Jinkela_wire_7916;
    wire new_Jinkela_wire_2668;
    wire new_Jinkela_wire_2124;
    wire new_Jinkela_wire_6705;
    wire new_Jinkela_wire_5234;
    wire new_Jinkela_wire_5555;
    wire new_Jinkela_wire_2630;
    wire new_Jinkela_wire_9787;
    wire new_Jinkela_wire_7392;
    wire new_Jinkela_wire_9040;
    wire new_Jinkela_wire_10168;
    wire n_0446_;
    wire n_1359_;
    wire new_Jinkela_wire_4948;
    wire new_Jinkela_wire_7672;
    wire new_Jinkela_wire_4885;
    wire new_Jinkela_wire_648;
    wire new_Jinkela_wire_9566;
    wire new_Jinkela_wire_4698;
    wire new_Jinkela_wire_2143;
    wire new_Jinkela_wire_4307;
    wire new_Jinkela_wire_10259;
    wire new_Jinkela_wire_8199;
    wire new_Jinkela_wire_8663;
    wire new_Jinkela_wire_121;
    wire new_Jinkela_wire_4162;
    wire new_Jinkela_wire_9612;
    wire n_0799_;
    wire new_Jinkela_wire_1185;
    wire new_Jinkela_wire_4126;
    wire new_Jinkela_wire_3688;
    wire new_Jinkela_wire_3261;
    wire new_Jinkela_wire_1551;
    wire new_Jinkela_wire_8228;
    wire new_Jinkela_wire_3294;
    wire new_Jinkela_wire_5229;
    wire new_Jinkela_wire_9683;
    wire n_0163_;
    wire new_Jinkela_wire_8348;
    wire n_0407_;
    wire new_Jinkela_wire_10434;
    wire new_Jinkela_wire_5651;
    wire new_Jinkela_wire_7232;
    wire new_Jinkela_wire_4107;
    wire new_Jinkela_wire_4473;
    wire new_Jinkela_wire_203;
    wire new_Jinkela_wire_6661;
    wire n_0728_;
    wire new_Jinkela_wire_3749;
    wire new_Jinkela_wire_6664;
    wire new_Jinkela_wire_2060;
    wire new_Jinkela_wire_1778;
    wire new_Jinkela_wire_8818;
    wire new_Jinkela_wire_5558;
    wire new_Jinkela_wire_8317;
    wire new_Jinkela_wire_5808;
    wire new_Jinkela_wire_5777;
    wire n_0800_;
    wire new_Jinkela_wire_863;
    wire new_Jinkela_wire_3707;
    wire new_Jinkela_wire_3727;
    wire new_Jinkela_wire_6085;
    wire new_Jinkela_wire_3240;
    wire new_Jinkela_wire_2399;
    wire new_Jinkela_wire_1009;
    wire new_Jinkela_wire_9978;
    wire new_Jinkela_wire_4291;
    wire new_Jinkela_wire_8682;
    wire new_Jinkela_wire_9766;
    wire new_Jinkela_wire_7364;
    wire new_Jinkela_wire_7742;
    wire new_Jinkela_wire_6968;
    wire new_Jinkela_wire_146;
    wire new_Jinkela_wire_9812;
    wire new_Jinkela_wire_10095;
    wire new_Jinkela_wire_2835;
    wire new_Jinkela_wire_5014;
    wire n_1144_;
    wire n_0460_;
    input N1;
    input N164;
    input N160;
    input N82;
    input N188;
    input N152;
    input N84;
    input N174;
    input N180;
    input N55;
    input N57;
    input N65;
    input N144;
    input N343;
    input N85;
    input N41;
    input N151;
    input N211;
    input N175;
    input N183;
    input N207;
    input N210;
    input N26;
    input N162;
    input N150;
    input N346;
    input N166;
    input N319;
    input N59;
    input N156;
    input N182;
    input N38;
    input N115;
    input N337;
    input N87;
    input N219;
    input N229;
    input N289;
    input N69;
    input N352;
    input N44;
    input N133;
    input N214;
    input N109;
    input N97;
    input N240;
    input N271;
    input N88;
    input N86;
    input N242;
    input N260;
    input N189;
    input N199;
    input N186;
    input N158;
    input N198;
    input N334;
    input N118;
    input N89;
    input N212;
    input N168;
    input N205;
    input N224;
    input N64;
    input N208;
    input N155;
    input N94;
    input N9;
    input N361;
    input N195;
    input N231;
    input N124;
    input N316;
    input N293;
    input N364;
    input N232;
    input N121;
    input N78;
    input N307;
    input N245;
    input N18;
    input N179;
    input N141;
    input N280;
    input N328;
    input N358;
    input N134;
    input N239;
    input N296;
    input N81;
    input N202;
    input N29;
    input N79;
    input N163;
    input N165;
    input N217;
    input N254;
    input N193;
    input N53;
    input N80;
    input N157;
    input N154;
    input N197;
    input N218;
    input N181;
    input N196;
    input N111;
    input N167;
    input N237;
    input N112;
    input N113;
    input N172;
    input N223;
    input N106;
    input N73;
    input N263;
    input N74;
    input N203;
    input N206;
    input N76;
    input N213;
    input N135;
    input N248;
    input N32;
    input N12;
    input N226;
    input N77;
    input N201;
    input N286;
    input N170;
    input N227;
    input N236;
    input N331;
    input N184;
    input N176;
    input N310;
    input N355;
    input N173;
    input N349;
    input N190;
    input N235;
    input N47;
    input N221;
    input N153;
    input N178;
    input N191;
    input N130;
    input N257;
    input N62;
    input N200;
    input N228;
    input N230;
    input N367;
    input N66;
    input N70;
    input N185;
    input N277;
    input N233;
    input N299;
    input N234;
    input N313;
    input N83;
    input N159;
    input N177;
    input N251;
    input N103;
    input N58;
    input N216;
    input N220;
    input N241_I;
    input N187;
    input N60;
    input N267;
    input N204;
    input N325;
    input N15;
    input N75;
    input N303;
    input N61;
    input N171;
    input N56;
    input N340;
    input N322;
    input N138;
    input N194;
    input N23;
    input N161;
    input N54;
    input N225;
    input N283;
    input N147;
    input N127;
    input N110;
    input N274;
    input N100;
    input N222;
    input N382;
    input N238;
    input N169;
    input N35;
    input N5;
    input N114;
    input N50;
    input N209;
    input N215;
    input N192;
    input N63;
    output N707;
    output N492;
    output N10714;
    output N10576;
    output N884;
    output N505;
    output N10907;
    output N10869;
    output N10101;
    output N10350;
    output N387;
    output N10762;
    output N567;
    output N11334;
    output N10704;
    output N509;
    output N10104;
    output N10760;
    output N535;
    output N10871;
    output N1110;
    output N10870;
    output N10632;
    output N11333;
    output N545;
    output N513;
    output N882;
    output N10759;
    output N11342;
    output N10110;
    output N482;
    output N10575;
    output N10908;
    output N10717;
    output N569;
    output N11340;
    output N10641;
    output N10868;
    output N241_O;
    output N889;
    output N515;
    output N563;
    output N10713;
    output N10905;
    output N10729;
    output N10712;
    output N582;
    output N10574;
    output N541;
    output N561;
    output N883;
    output N881;
    output N553;
    output N10906;
    output N10761;
    output N556;
    output N10025;
    output N10353;
    output N1111;
    output N10112;
    output N486;
    output N571;
    output N10711;
    output N813;
    output N559;
    output N1114;
    output N1781;
    output N10715;
    output N10352;
    output N478;
    output N551;
    output N388;
    output N1112;
    output N489;
    output N517;
    output N10839;
    output N10763;
    output N10111;
    output N539;
    output N10840;
    output N543;
    output N10718;
    output N507;
    output N10109;
    output N501;
    output N565;
    output N10837;
    output N10716;
    output N643;
    output N1490;
    output N537;
    output N10838;
    output N10102;
    output N547;
    output N549;
    output N10628;
    output N10706;
    output N519;
    output N10103;
    output N885;
    output N484;
    output N10827;
    output N1489;
    output N10351;
    output N511;
    output N945;
    output N573;
    output N1113;

    bfr new_Jinkela_buffer_8112 (
        .din(new_Jinkela_wire_10206),
        .dout(new_Jinkela_wire_10207)
    );

    bfr new_Jinkela_buffer_8202 (
        .din(new_Jinkela_wire_10305),
        .dout(new_Jinkela_wire_10306)
    );

    bfr new_Jinkela_buffer_2784 (
        .din(new_Jinkela_wire_3198),
        .dout(new_Jinkela_wire_3199)
    );

    bfr new_Jinkela_buffer_8113 (
        .din(new_Jinkela_wire_10207),
        .dout(new_Jinkela_wire_10208)
    );

    bfr new_Jinkela_buffer_8151 (
        .din(new_Jinkela_wire_10252),
        .dout(new_Jinkela_wire_10253)
    );

    bfr new_Jinkela_buffer_8114 (
        .din(new_Jinkela_wire_10208),
        .dout(new_Jinkela_wire_10209)
    );

    bfr new_Jinkela_buffer_8244 (
        .din(new_Jinkela_wire_10347),
        .dout(new_Jinkela_wire_10348)
    );

    bfr new_Jinkela_buffer_8115 (
        .din(new_Jinkela_wire_10209),
        .dout(new_Jinkela_wire_10210)
    );

    bfr new_Jinkela_buffer_8152 (
        .din(new_Jinkela_wire_10253),
        .dout(new_Jinkela_wire_10254)
    );

    bfr new_Jinkela_buffer_8116 (
        .din(new_Jinkela_wire_10210),
        .dout(new_Jinkela_wire_10211)
    );

    bfr new_Jinkela_buffer_8203 (
        .din(new_Jinkela_wire_10306),
        .dout(new_Jinkela_wire_10307)
    );

    bfr new_Jinkela_buffer_8117 (
        .din(new_Jinkela_wire_10211),
        .dout(new_Jinkela_wire_10212)
    );

    bfr new_Jinkela_buffer_8153 (
        .din(new_Jinkela_wire_10254),
        .dout(new_Jinkela_wire_10255)
    );

    bfr new_Jinkela_buffer_2663 (
        .din(new_Jinkela_wire_3072),
        .dout(new_Jinkela_wire_3073)
    );

    bfr new_Jinkela_buffer_8118 (
        .din(new_Jinkela_wire_10212),
        .dout(new_Jinkela_wire_10213)
    );

    spl2 new_Jinkela_splitter_849 (
        .a(n_0020_),
        .b(new_Jinkela_wire_10382),
        .c(new_Jinkela_wire_10383)
    );

    bfr new_Jinkela_buffer_8119 (
        .din(new_Jinkela_wire_10213),
        .dout(new_Jinkela_wire_10214)
    );

    bfr new_Jinkela_buffer_8154 (
        .din(new_Jinkela_wire_10255),
        .dout(new_Jinkela_wire_10256)
    );

    bfr new_Jinkela_buffer_8120 (
        .din(new_Jinkela_wire_10214),
        .dout(new_Jinkela_wire_10215)
    );

    bfr new_Jinkela_buffer_8204 (
        .din(new_Jinkela_wire_10307),
        .dout(new_Jinkela_wire_10308)
    );

    bfr new_Jinkela_buffer_8121 (
        .din(new_Jinkela_wire_10215),
        .dout(new_Jinkela_wire_10216)
    );

    bfr new_Jinkela_buffer_8155 (
        .din(new_Jinkela_wire_10256),
        .dout(new_Jinkela_wire_10257)
    );

    bfr new_Jinkela_buffer_8122 (
        .din(new_Jinkela_wire_10216),
        .dout(new_Jinkela_wire_10217)
    );

    bfr new_Jinkela_buffer_8256 (
        .din(new_Jinkela_wire_10368),
        .dout(new_Jinkela_wire_10369)
    );

    bfr new_Jinkela_buffer_8245 (
        .din(new_Jinkela_wire_10348),
        .dout(new_Jinkela_wire_10349)
    );

    bfr new_Jinkela_buffer_2718 (
        .din(new_Jinkela_wire_3132),
        .dout(new_Jinkela_wire_3133)
    );

    bfr new_Jinkela_buffer_8123 (
        .din(new_Jinkela_wire_10217),
        .dout(new_Jinkela_wire_10218)
    );

    bfr new_Jinkela_buffer_8156 (
        .din(new_Jinkela_wire_10257),
        .dout(new_Jinkela_wire_10258)
    );

    bfr new_Jinkela_buffer_8205 (
        .din(new_Jinkela_wire_10308),
        .dout(new_Jinkela_wire_10309)
    );

    bfr new_Jinkela_buffer_8157 (
        .din(new_Jinkela_wire_10258),
        .dout(new_Jinkela_wire_10259)
    );

    spl2 new_Jinkela_splitter_850 (
        .a(n_0755_),
        .b(new_Jinkela_wire_10384),
        .c(new_Jinkela_wire_10385)
    );

    bfr new_Jinkela_buffer_8158 (
        .din(new_Jinkela_wire_10259),
        .dout(new_Jinkela_wire_10260)
    );

    bfr new_Jinkela_buffer_8206 (
        .din(new_Jinkela_wire_10309),
        .dout(new_Jinkela_wire_10310)
    );

    bfr new_Jinkela_buffer_8159 (
        .din(new_Jinkela_wire_10260),
        .dout(new_Jinkela_wire_10261)
    );

    bfr new_Jinkela_buffer_8257 (
        .din(new_Jinkela_wire_10369),
        .dout(new_Jinkela_wire_10370)
    );

    bfr new_Jinkela_buffer_8246 (
        .din(new_Jinkela_wire_10349),
        .dout(new_Jinkela_wire_10350)
    );

    bfr new_Jinkela_buffer_8160 (
        .din(new_Jinkela_wire_10261),
        .dout(new_Jinkela_wire_10262)
    );

    bfr new_Jinkela_buffer_8207 (
        .din(new_Jinkela_wire_10310),
        .dout(new_Jinkela_wire_10311)
    );

    bfr new_Jinkela_buffer_8161 (
        .din(new_Jinkela_wire_10262),
        .dout(new_Jinkela_wire_10263)
    );

    bfr new_Jinkela_buffer_8162 (
        .din(new_Jinkela_wire_10263),
        .dout(new_Jinkela_wire_10264)
    );

    bfr new_Jinkela_buffer_8208 (
        .din(new_Jinkela_wire_10311),
        .dout(new_Jinkela_wire_10312)
    );

    bfr new_Jinkela_buffer_8163 (
        .din(new_Jinkela_wire_10264),
        .dout(new_Jinkela_wire_10265)
    );

    bfr new_Jinkela_buffer_8247 (
        .din(new_Jinkela_wire_10350),
        .dout(new_Jinkela_wire_10351)
    );

    bfr new_Jinkela_buffer_8164 (
        .din(new_Jinkela_wire_10265),
        .dout(new_Jinkela_wire_10266)
    );

    bfr new_Jinkela_buffer_8209 (
        .din(new_Jinkela_wire_10312),
        .dout(new_Jinkela_wire_10313)
    );

    bfr new_Jinkela_buffer_8165 (
        .din(new_Jinkela_wire_10266),
        .dout(new_Jinkela_wire_10267)
    );

    bfr new_Jinkela_buffer_3691 (
        .din(new_Jinkela_wire_4305),
        .dout(new_Jinkela_wire_4306)
    );

    bfr new_Jinkela_buffer_3772 (
        .din(new_Jinkela_wire_4394),
        .dout(new_Jinkela_wire_4395)
    );

    spl2 new_Jinkela_splitter_805 (
        .a(new_Jinkela_wire_9752),
        .b(new_Jinkela_wire_9753),
        .c(new_Jinkela_wire_9754)
    );

    bfr new_Jinkela_buffer_3696 (
        .din(new_Jinkela_wire_4314),
        .dout(new_Jinkela_wire_4315)
    );

    bfr new_Jinkela_buffer_7686 (
        .din(new_Jinkela_wire_9672),
        .dout(new_Jinkela_wire_9673)
    );

    bfr new_Jinkela_buffer_3720 (
        .din(new_Jinkela_wire_4340),
        .dout(new_Jinkela_wire_4341)
    );

    bfr new_Jinkela_buffer_7722 (
        .din(new_Jinkela_wire_9718),
        .dout(new_Jinkela_wire_9719)
    );

    bfr new_Jinkela_buffer_3697 (
        .din(new_Jinkela_wire_4315),
        .dout(new_Jinkela_wire_4316)
    );

    bfr new_Jinkela_buffer_7687 (
        .din(new_Jinkela_wire_9673),
        .dout(new_Jinkela_wire_9674)
    );

    spl2 new_Jinkela_splitter_808 (
        .a(n_1015_),
        .b(new_Jinkela_wire_9761),
        .c(new_Jinkela_wire_9762)
    );

    bfr new_Jinkela_buffer_3805 (
        .din(n_0969_),
        .dout(new_Jinkela_wire_4428)
    );

    bfr new_Jinkela_buffer_7738 (
        .din(new_Jinkela_wire_9736),
        .dout(new_Jinkela_wire_9737)
    );

    bfr new_Jinkela_buffer_3698 (
        .din(new_Jinkela_wire_4316),
        .dout(new_Jinkela_wire_4317)
    );

    bfr new_Jinkela_buffer_7688 (
        .din(new_Jinkela_wire_9674),
        .dout(new_Jinkela_wire_9675)
    );

    bfr new_Jinkela_buffer_3721 (
        .din(new_Jinkela_wire_4341),
        .dout(new_Jinkela_wire_4342)
    );

    bfr new_Jinkela_buffer_7723 (
        .din(new_Jinkela_wire_9719),
        .dout(new_Jinkela_wire_9720)
    );

    bfr new_Jinkela_buffer_3699 (
        .din(new_Jinkela_wire_4317),
        .dout(new_Jinkela_wire_4318)
    );

    bfr new_Jinkela_buffer_7689 (
        .din(new_Jinkela_wire_9675),
        .dout(new_Jinkela_wire_9676)
    );

    spl3L new_Jinkela_splitter_226 (
        .a(n_0072_),
        .d(new_Jinkela_wire_4432),
        .b(new_Jinkela_wire_4433),
        .c(new_Jinkela_wire_4434)
    );

    bfr new_Jinkela_buffer_3773 (
        .din(new_Jinkela_wire_4395),
        .dout(new_Jinkela_wire_4396)
    );

    bfr new_Jinkela_buffer_3700 (
        .din(new_Jinkela_wire_4318),
        .dout(new_Jinkela_wire_4319)
    );

    bfr new_Jinkela_buffer_7690 (
        .din(new_Jinkela_wire_9676),
        .dout(new_Jinkela_wire_9677)
    );

    bfr new_Jinkela_buffer_3722 (
        .din(new_Jinkela_wire_4342),
        .dout(new_Jinkela_wire_4343)
    );

    bfr new_Jinkela_buffer_7724 (
        .din(new_Jinkela_wire_9720),
        .dout(new_Jinkela_wire_9721)
    );

    bfr new_Jinkela_buffer_3701 (
        .din(new_Jinkela_wire_4319),
        .dout(new_Jinkela_wire_4320)
    );

    bfr new_Jinkela_buffer_7691 (
        .din(new_Jinkela_wire_9677),
        .dout(new_Jinkela_wire_9678)
    );

    bfr new_Jinkela_buffer_3789 (
        .din(new_Jinkela_wire_4411),
        .dout(new_Jinkela_wire_4412)
    );

    spl2 new_Jinkela_splitter_801 (
        .a(new_Jinkela_wire_9737),
        .b(new_Jinkela_wire_9738),
        .c(new_Jinkela_wire_9739)
    );

    bfr new_Jinkela_buffer_3702 (
        .din(new_Jinkela_wire_4320),
        .dout(new_Jinkela_wire_4321)
    );

    bfr new_Jinkela_buffer_7692 (
        .din(new_Jinkela_wire_9678),
        .dout(new_Jinkela_wire_9679)
    );

    bfr new_Jinkela_buffer_3723 (
        .din(new_Jinkela_wire_4343),
        .dout(new_Jinkela_wire_4344)
    );

    bfr new_Jinkela_buffer_7725 (
        .din(new_Jinkela_wire_9721),
        .dout(new_Jinkela_wire_9722)
    );

    bfr new_Jinkela_buffer_3703 (
        .din(new_Jinkela_wire_4321),
        .dout(new_Jinkela_wire_4322)
    );

    bfr new_Jinkela_buffer_7693 (
        .din(new_Jinkela_wire_9679),
        .dout(new_Jinkela_wire_9680)
    );

    bfr new_Jinkela_buffer_3774 (
        .din(new_Jinkela_wire_4396),
        .dout(new_Jinkela_wire_4397)
    );

    bfr new_Jinkela_buffer_7739 (
        .din(new_Jinkela_wire_9739),
        .dout(new_Jinkela_wire_9740)
    );

    bfr new_Jinkela_buffer_3704 (
        .din(new_Jinkela_wire_4322),
        .dout(new_Jinkela_wire_4323)
    );

    bfr new_Jinkela_buffer_7694 (
        .din(new_Jinkela_wire_9680),
        .dout(new_Jinkela_wire_9681)
    );

    bfr new_Jinkela_buffer_3724 (
        .din(new_Jinkela_wire_4344),
        .dout(new_Jinkela_wire_4345)
    );

    bfr new_Jinkela_buffer_7726 (
        .din(new_Jinkela_wire_9722),
        .dout(new_Jinkela_wire_9723)
    );

    bfr new_Jinkela_buffer_3705 (
        .din(new_Jinkela_wire_4323),
        .dout(new_Jinkela_wire_4324)
    );

    bfr new_Jinkela_buffer_7695 (
        .din(new_Jinkela_wire_9681),
        .dout(new_Jinkela_wire_9682)
    );

    bfr new_Jinkela_buffer_3806 (
        .din(new_Jinkela_wire_4428),
        .dout(new_Jinkela_wire_4429)
    );

    bfr new_Jinkela_buffer_7743 (
        .din(new_Jinkela_wire_9758),
        .dout(new_Jinkela_wire_9759)
    );

    bfr new_Jinkela_buffer_3706 (
        .din(new_Jinkela_wire_4324),
        .dout(new_Jinkela_wire_4325)
    );

    bfr new_Jinkela_buffer_7696 (
        .din(new_Jinkela_wire_9682),
        .dout(new_Jinkela_wire_9683)
    );

    bfr new_Jinkela_buffer_3725 (
        .din(new_Jinkela_wire_4345),
        .dout(new_Jinkela_wire_4346)
    );

    bfr new_Jinkela_buffer_7727 (
        .din(new_Jinkela_wire_9723),
        .dout(new_Jinkela_wire_9724)
    );

    bfr new_Jinkela_buffer_3707 (
        .din(new_Jinkela_wire_4325),
        .dout(new_Jinkela_wire_4326)
    );

    bfr new_Jinkela_buffer_7697 (
        .din(new_Jinkela_wire_9683),
        .dout(new_Jinkela_wire_9684)
    );

    bfr new_Jinkela_buffer_3775 (
        .din(new_Jinkela_wire_4397),
        .dout(new_Jinkela_wire_4398)
    );

    bfr new_Jinkela_buffer_3708 (
        .din(new_Jinkela_wire_4326),
        .dout(new_Jinkela_wire_4327)
    );

    bfr new_Jinkela_buffer_7698 (
        .din(new_Jinkela_wire_9684),
        .dout(new_Jinkela_wire_9685)
    );

    bfr new_Jinkela_buffer_3726 (
        .din(new_Jinkela_wire_4346),
        .dout(new_Jinkela_wire_4347)
    );

    bfr new_Jinkela_buffer_7728 (
        .din(new_Jinkela_wire_9724),
        .dout(new_Jinkela_wire_9725)
    );

    bfr new_Jinkela_buffer_3709 (
        .din(new_Jinkela_wire_4327),
        .dout(new_Jinkela_wire_4328)
    );

    bfr new_Jinkela_buffer_7699 (
        .din(new_Jinkela_wire_9685),
        .dout(new_Jinkela_wire_9686)
    );

    spl4L new_Jinkela_splitter_809 (
        .a(n_0872_),
        .d(new_Jinkela_wire_9763),
        .b(new_Jinkela_wire_9764),
        .e(new_Jinkela_wire_9765),
        .c(new_Jinkela_wire_9766)
    );

    bfr new_Jinkela_buffer_3790 (
        .din(new_Jinkela_wire_4412),
        .dout(new_Jinkela_wire_4413)
    );

    spl2 new_Jinkela_splitter_802 (
        .a(new_Jinkela_wire_9740),
        .b(new_Jinkela_wire_9741),
        .c(new_Jinkela_wire_9742)
    );

    bfr new_Jinkela_buffer_3710 (
        .din(new_Jinkela_wire_4328),
        .dout(new_Jinkela_wire_4329)
    );

    bfr new_Jinkela_buffer_7700 (
        .din(new_Jinkela_wire_9686),
        .dout(new_Jinkela_wire_9687)
    );

    bfr new_Jinkela_buffer_3727 (
        .din(new_Jinkela_wire_4347),
        .dout(new_Jinkela_wire_4348)
    );

    bfr new_Jinkela_buffer_7729 (
        .din(new_Jinkela_wire_9725),
        .dout(new_Jinkela_wire_9726)
    );

    bfr new_Jinkela_buffer_3711 (
        .din(new_Jinkela_wire_4329),
        .dout(new_Jinkela_wire_4330)
    );

    bfr new_Jinkela_buffer_7701 (
        .din(new_Jinkela_wire_9687),
        .dout(new_Jinkela_wire_9688)
    );

    bfr new_Jinkela_buffer_3776 (
        .din(new_Jinkela_wire_4398),
        .dout(new_Jinkela_wire_4399)
    );

    bfr new_Jinkela_buffer_7740 (
        .din(new_Jinkela_wire_9742),
        .dout(new_Jinkela_wire_9743)
    );

    bfr new_Jinkela_buffer_3712 (
        .din(new_Jinkela_wire_4330),
        .dout(new_Jinkela_wire_4331)
    );

    bfr new_Jinkela_buffer_7702 (
        .din(new_Jinkela_wire_9688),
        .dout(new_Jinkela_wire_9689)
    );

    bfr new_Jinkela_buffer_3728 (
        .din(new_Jinkela_wire_4348),
        .dout(new_Jinkela_wire_4349)
    );

    bfr new_Jinkela_buffer_7730 (
        .din(new_Jinkela_wire_9726),
        .dout(new_Jinkela_wire_9727)
    );

    bfr new_Jinkela_buffer_3713 (
        .din(new_Jinkela_wire_4331),
        .dout(new_Jinkela_wire_4332)
    );

    bfr new_Jinkela_buffer_7703 (
        .din(new_Jinkela_wire_9689),
        .dout(new_Jinkela_wire_9690)
    );

    spl2 new_Jinkela_splitter_227 (
        .a(n_1335_),
        .b(new_Jinkela_wire_4435),
        .c(new_Jinkela_wire_4436)
    );

    bfr new_Jinkela_buffer_7745 (
        .din(n_0858_),
        .dout(new_Jinkela_wire_9767)
    );

    bfr new_Jinkela_buffer_3714 (
        .din(new_Jinkela_wire_4332),
        .dout(new_Jinkela_wire_4333)
    );

    bfr new_Jinkela_buffer_7704 (
        .din(new_Jinkela_wire_9690),
        .dout(new_Jinkela_wire_9691)
    );

    bfr new_Jinkela_buffer_3729 (
        .din(new_Jinkela_wire_4349),
        .dout(new_Jinkela_wire_4350)
    );

    bfr new_Jinkela_buffer_7731 (
        .din(new_Jinkela_wire_9727),
        .dout(new_Jinkela_wire_9728)
    );

    bfr new_Jinkela_buffer_3715 (
        .din(new_Jinkela_wire_4333),
        .dout(new_Jinkela_wire_4334)
    );

    bfr new_Jinkela_buffer_7705 (
        .din(new_Jinkela_wire_9691),
        .dout(new_Jinkela_wire_9692)
    );

    bfr new_Jinkela_buffer_3777 (
        .din(new_Jinkela_wire_4399),
        .dout(new_Jinkela_wire_4400)
    );

    bfr new_Jinkela_buffer_7744 (
        .din(new_Jinkela_wire_9759),
        .dout(new_Jinkela_wire_9760)
    );

    bfr new_Jinkela_buffer_3716 (
        .din(new_Jinkela_wire_4334),
        .dout(new_Jinkela_wire_4335)
    );

    bfr new_Jinkela_buffer_7706 (
        .din(new_Jinkela_wire_9692),
        .dout(new_Jinkela_wire_9693)
    );

    bfr new_Jinkela_buffer_2930 (
        .din(new_Jinkela_wire_3353),
        .dout(new_Jinkela_wire_3354)
    );

    or_bb n_1485_ (
        .a(new_Jinkela_wire_5101),
        .b(new_Jinkela_wire_6252),
        .c(n_0753_)
    );

    and_bi n_2199_ (
        .a(new_Jinkela_wire_7304),
        .b(new_Jinkela_wire_3768),
        .c(n_0089_)
    );

    bfr new_Jinkela_buffer_2821 (
        .din(new_Jinkela_wire_3240),
        .dout(new_Jinkela_wire_3241)
    );

    and_bb n_1486_ (
        .a(new_Jinkela_wire_5100),
        .b(new_Jinkela_wire_6251),
        .c(n_0754_)
    );

    and_bi n_2200_ (
        .a(new_Jinkela_wire_3767),
        .b(new_Jinkela_wire_7303),
        .c(n_0090_)
    );

    bfr new_Jinkela_buffer_2867 (
        .din(new_Jinkela_wire_3290),
        .dout(new_Jinkela_wire_3291)
    );

    and_bi n_1487_ (
        .a(n_0753_),
        .b(n_0754_),
        .c(n_0755_)
    );

    or_bb n_2201_ (
        .a(n_0090_),
        .b(n_0089_),
        .c(new_net_2517)
    );

    bfr new_Jinkela_buffer_2822 (
        .din(new_Jinkela_wire_3241),
        .dout(new_Jinkela_wire_3242)
    );

    and_bi n_1488_ (
        .a(new_Jinkela_wire_3342),
        .b(new_Jinkela_wire_1212),
        .c(n_0756_)
    );

    and_bi n_2202_ (
        .a(new_Jinkela_wire_7446),
        .b(new_Jinkela_wire_8381),
        .c(n_0091_)
    );

    spl2 new_Jinkela_splitter_144 (
        .a(N283),
        .b(new_Jinkela_wire_3363),
        .c(new_Jinkela_wire_3364)
    );

    and_bb n_1489_ (
        .a(new_Jinkela_wire_75),
        .b(new_Jinkela_wire_1335),
        .c(n_0757_)
    );

    and_bi n_2203_ (
        .a(new_Jinkela_wire_7803),
        .b(n_0091_),
        .c(n_0092_)
    );

    bfr new_Jinkela_buffer_3003 (
        .din(N147),
        .dout(new_Jinkela_wire_3431)
    );

    bfr new_Jinkela_buffer_2823 (
        .din(new_Jinkela_wire_3242),
        .dout(new_Jinkela_wire_3243)
    );

    and_ii n_1490_ (
        .a(new_Jinkela_wire_6767),
        .b(new_Jinkela_wire_9550),
        .c(n_0758_)
    );

    and_bi n_2204_ (
        .a(new_Jinkela_wire_5968),
        .b(new_Jinkela_wire_7448),
        .c(n_0093_)
    );

    bfr new_Jinkela_buffer_2868 (
        .din(new_Jinkela_wire_3291),
        .dout(new_Jinkela_wire_3292)
    );

    and_bi n_1491_ (
        .a(new_Jinkela_wire_104),
        .b(new_Jinkela_wire_1294),
        .c(n_0759_)
    );

    and_bi n_2205_ (
        .a(new_Jinkela_wire_7447),
        .b(new_Jinkela_wire_5969),
        .c(n_0094_)
    );

    bfr new_Jinkela_buffer_2824 (
        .din(new_Jinkela_wire_3243),
        .dout(new_Jinkela_wire_3244)
    );

    bfr new_Jinkela_buffer_2667 (
        .din(new_Jinkela_wire_3076),
        .dout(new_Jinkela_wire_3077)
    );

    and_bb n_1492_ (
        .a(new_Jinkela_wire_2812),
        .b(new_Jinkela_wire_1383),
        .c(n_0760_)
    );

    or_bb n_2206_ (
        .a(n_0094_),
        .b(n_0093_),
        .c(new_net_2564)
    );

    bfr new_Jinkela_buffer_2933 (
        .din(new_Jinkela_wire_3356),
        .dout(new_Jinkela_wire_3357)
    );

    and_ii n_1493_ (
        .a(new_Jinkela_wire_7541),
        .b(new_Jinkela_wire_4338),
        .c(n_0761_)
    );

    and_ii n_2207_ (
        .a(new_Jinkela_wire_10382),
        .b(new_Jinkela_wire_7499),
        .c(n_0095_)
    );

    bfr new_Jinkela_buffer_2825 (
        .din(new_Jinkela_wire_3244),
        .dout(new_Jinkela_wire_3245)
    );

    and_ii n_1494_ (
        .a(new_Jinkela_wire_3864),
        .b(new_Jinkela_wire_5159),
        .c(n_0762_)
    );

    or_ii n_2208_ (
        .a(new_Jinkela_wire_7841),
        .b(new_Jinkela_wire_9289),
        .c(n_0096_)
    );

    bfr new_Jinkela_buffer_2869 (
        .din(new_Jinkela_wire_3292),
        .dout(new_Jinkela_wire_3293)
    );

    and_bb n_1495_ (
        .a(new_Jinkela_wire_3863),
        .b(new_Jinkela_wire_5160),
        .c(n_0763_)
    );

    or_bb n_2209_ (
        .a(new_Jinkela_wire_7840),
        .b(new_Jinkela_wire_9290),
        .c(n_0097_)
    );

    bfr new_Jinkela_buffer_2826 (
        .din(new_Jinkela_wire_3245),
        .dout(new_Jinkela_wire_3246)
    );

    or_bb n_1496_ (
        .a(n_0763_),
        .b(n_0762_),
        .c(n_0764_)
    );

    or_ii n_2210_ (
        .a(n_0097_),
        .b(n_0096_),
        .c(new_net_2495)
    );

    bfr new_Jinkela_buffer_2936 (
        .din(new_Jinkela_wire_3359),
        .dout(new_Jinkela_wire_3360)
    );

    and_ii n_1497_ (
        .a(new_Jinkela_wire_3854),
        .b(new_Jinkela_wire_10385),
        .c(n_0765_)
    );

    and_bi n_2211_ (
        .a(new_Jinkela_wire_4173),
        .b(new_Jinkela_wire_2488),
        .c(n_0098_)
    );

    bfr new_Jinkela_buffer_2827 (
        .din(new_Jinkela_wire_3246),
        .dout(new_Jinkela_wire_3247)
    );

    and_bb n_1498_ (
        .a(new_Jinkela_wire_3853),
        .b(new_Jinkela_wire_10384),
        .c(n_0766_)
    );

    and_bi n_2212_ (
        .a(new_Jinkela_wire_2487),
        .b(new_Jinkela_wire_4174),
        .c(n_0099_)
    );

    bfr new_Jinkela_buffer_2870 (
        .din(new_Jinkela_wire_3293),
        .dout(new_Jinkela_wire_3294)
    );

    and_ii n_1499_ (
        .a(n_0766_),
        .b(n_0765_),
        .c(n_0767_)
    );

    and_bi n_2213_ (
        .a(new_Jinkela_wire_7090),
        .b(new_Jinkela_wire_1840),
        .c(n_0100_)
    );

    bfr new_Jinkela_buffer_2828 (
        .din(new_Jinkela_wire_3247),
        .dout(new_Jinkela_wire_3248)
    );

    and_bb n_1500_ (
        .a(new_Jinkela_wire_3933),
        .b(new_Jinkela_wire_4964),
        .c(n_0768_)
    );

    inv n_2214_ (
        .din(new_Jinkela_wire_8178),
        .dout(n_0101_)
    );

    bfr new_Jinkela_buffer_2934 (
        .din(new_Jinkela_wire_3357),
        .dout(new_Jinkela_wire_3358)
    );

    and_bi n_2215_ (
        .a(new_Jinkela_wire_1839),
        .b(new_Jinkela_wire_7089),
        .c(n_0102_)
    );

    and_bi n_1501_ (
        .a(new_Jinkela_wire_1298),
        .b(new_Jinkela_wire_3550),
        .c(n_0769_)
    );

    bfr new_Jinkela_buffer_2829 (
        .din(new_Jinkela_wire_3248),
        .dout(new_Jinkela_wire_3249)
    );

    bfr new_Jinkela_buffer_2720 (
        .din(new_Jinkela_wire_3134),
        .dout(new_Jinkela_wire_3135)
    );

    and_bi n_2216_ (
        .a(new_Jinkela_wire_1714),
        .b(new_Jinkela_wire_7069),
        .c(n_0103_)
    );

    and_bi n_1502_ (
        .a(new_Jinkela_wire_4528),
        .b(new_Jinkela_wire_9457),
        .c(n_0770_)
    );

    bfr new_Jinkela_buffer_2871 (
        .din(new_Jinkela_wire_3294),
        .dout(new_Jinkela_wire_3295)
    );

    and_bi n_2217_ (
        .a(new_Jinkela_wire_7070),
        .b(new_Jinkela_wire_1715),
        .c(n_0104_)
    );

    and_bi n_1503_ (
        .a(new_Jinkela_wire_1263),
        .b(new_Jinkela_wire_590),
        .c(n_0771_)
    );

    bfr new_Jinkela_buffer_2830 (
        .din(new_Jinkela_wire_3249),
        .dout(new_Jinkela_wire_3250)
    );

    and_ii n_2218_ (
        .a(new_Jinkela_wire_5571),
        .b(new_Jinkela_wire_6436),
        .c(n_0105_)
    );

    and_ii n_1504_ (
        .a(new_Jinkela_wire_9366),
        .b(new_Jinkela_wire_9442),
        .c(n_0772_)
    );

    or_bb n_2219_ (
        .a(new_Jinkela_wire_9142),
        .b(new_Jinkela_wire_8269),
        .c(n_0106_)
    );

    and_bi n_1505_ (
        .a(new_Jinkela_wire_1256),
        .b(new_Jinkela_wire_1993),
        .c(n_0773_)
    );

    bfr new_Jinkela_buffer_3004 (
        .din(new_Jinkela_wire_3431),
        .dout(new_Jinkela_wire_3432)
    );

    bfr new_Jinkela_buffer_2831 (
        .din(new_Jinkela_wire_3250),
        .dout(new_Jinkela_wire_3251)
    );

    and_ii n_2220_ (
        .a(new_Jinkela_wire_6016),
        .b(new_Jinkela_wire_10153),
        .c(n_0107_)
    );

    and_bb n_1506_ (
        .a(new_Jinkela_wire_9760),
        .b(new_Jinkela_wire_4175),
        .c(n_0774_)
    );

    bfr new_Jinkela_buffer_2872 (
        .din(new_Jinkela_wire_3295),
        .dout(new_Jinkela_wire_3296)
    );

    and_bi n_2221_ (
        .a(new_Jinkela_wire_4180),
        .b(n_0107_),
        .c(n_0108_)
    );

    and_ii n_1507_ (
        .a(new_Jinkela_wire_9757),
        .b(new_Jinkela_wire_9454),
        .c(n_0775_)
    );

    bfr new_Jinkela_buffer_2832 (
        .din(new_Jinkela_wire_3251),
        .dout(new_Jinkela_wire_3252)
    );

    and_ii n_2222_ (
        .a(new_Jinkela_wire_6194),
        .b(new_Jinkela_wire_5892),
        .c(n_0109_)
    );

    and_bb n_1508_ (
        .a(new_Jinkela_wire_9619),
        .b(new_Jinkela_wire_9369),
        .c(n_0776_)
    );

    bfr new_Jinkela_buffer_2937 (
        .din(new_Jinkela_wire_3360),
        .dout(new_Jinkela_wire_3361)
    );

    and_ii n_2223_ (
        .a(n_0109_),
        .b(new_Jinkela_wire_10377),
        .c(n_0110_)
    );

    and_ii n_1509_ (
        .a(n_0776_),
        .b(n_0774_),
        .c(n_0777_)
    );

    bfr new_Jinkela_buffer_2833 (
        .din(new_Jinkela_wire_3252),
        .dout(new_Jinkela_wire_3253)
    );

    and_ii n_2224_ (
        .a(new_Jinkela_wire_10148),
        .b(new_Jinkela_wire_8177),
        .c(n_0111_)
    );

    or_bi n_1510_ (
        .a(new_Jinkela_wire_7363),
        .b(new_Jinkela_wire_8295),
        .c(n_0778_)
    );

    bfr new_Jinkela_buffer_2873 (
        .din(new_Jinkela_wire_3296),
        .dout(new_Jinkela_wire_3297)
    );

    and_ii n_2225_ (
        .a(new_Jinkela_wire_8266),
        .b(new_Jinkela_wire_5570),
        .c(n_0112_)
    );

    and_bi n_1511_ (
        .a(new_Jinkela_wire_7362),
        .b(new_Jinkela_wire_8294),
        .c(n_0779_)
    );

    bfr new_Jinkela_buffer_2834 (
        .din(new_Jinkela_wire_3253),
        .dout(new_Jinkela_wire_3254)
    );

    or_ii n_2226_ (
        .a(new_Jinkela_wire_5756),
        .b(new_Jinkela_wire_9201),
        .c(n_0113_)
    );

    and_bi n_1512_ (
        .a(n_0778_),
        .b(n_0779_),
        .c(n_0780_)
    );

    and_bi n_2227_ (
        .a(new_Jinkela_wire_9043),
        .b(new_Jinkela_wire_7025),
        .c(n_0114_)
    );

    and_bi n_1513_ (
        .a(new_Jinkela_wire_1220),
        .b(new_Jinkela_wire_2897),
        .c(n_0781_)
    );

    bfr new_Jinkela_buffer_3007 (
        .din(N127),
        .dout(new_Jinkela_wire_3435)
    );

    bfr new_Jinkela_buffer_2835 (
        .din(new_Jinkela_wire_3254),
        .dout(new_Jinkela_wire_3255)
    );

    and_bi n_2228_ (
        .a(new_Jinkela_wire_7585),
        .b(new_Jinkela_wire_4529),
        .c(n_0115_)
    );

    and_ii n_1514_ (
        .a(new_Jinkela_wire_5288),
        .b(new_Jinkela_wire_9463),
        .c(n_0782_)
    );

    bfr new_Jinkela_buffer_2874 (
        .din(new_Jinkela_wire_3297),
        .dout(new_Jinkela_wire_3298)
    );

    and_ii n_2229_ (
        .a(new_Jinkela_wire_5883),
        .b(new_Jinkela_wire_10366),
        .c(n_0116_)
    );

    and_bi n_1515_ (
        .a(new_Jinkela_wire_1320),
        .b(new_Jinkela_wire_3554),
        .c(n_0783_)
    );

    bfr new_Jinkela_buffer_2836 (
        .din(new_Jinkela_wire_3255),
        .dout(new_Jinkela_wire_3256)
    );

    or_ii n_2230_ (
        .a(new_Jinkela_wire_9698),
        .b(new_Jinkela_wire_5878),
        .c(n_0117_)
    );

    and_bb n_1516_ (
        .a(new_Jinkela_wire_8096),
        .b(new_Jinkela_wire_7071),
        .c(n_0784_)
    );

    bfr new_Jinkela_buffer_2938 (
        .din(new_Jinkela_wire_3361),
        .dout(new_Jinkela_wire_3362)
    );

    or_ii n_2231_ (
        .a(n_0117_),
        .b(new_Jinkela_wire_4276),
        .c(n_0118_)
    );

    and_ii n_1517_ (
        .a(new_Jinkela_wire_8093),
        .b(new_Jinkela_wire_9444),
        .c(n_0785_)
    );

    bfr new_Jinkela_buffer_2837 (
        .din(new_Jinkela_wire_3256),
        .dout(new_Jinkela_wire_3257)
    );

    and_bb n_1518_ (
        .a(new_Jinkela_wire_7091),
        .b(new_Jinkela_wire_5291),
        .c(n_0786_)
    );

    and_bi n_2232_ (
        .a(new_Jinkela_wire_9618),
        .b(new_Jinkela_wire_619),
        .c(n_0119_)
    );

    bfr new_Jinkela_buffer_2875 (
        .din(new_Jinkela_wire_3298),
        .dout(new_Jinkela_wire_3299)
    );

    and_ii n_1519_ (
        .a(n_0786_),
        .b(n_0784_),
        .c(n_0787_)
    );

    and_bi n_2233_ (
        .a(new_Jinkela_wire_618),
        .b(new_Jinkela_wire_9617),
        .c(n_0120_)
    );

    bfr new_Jinkela_buffer_2838 (
        .din(new_Jinkela_wire_3257),
        .dout(new_Jinkela_wire_3258)
    );

    or_bi n_1520_ (
        .a(new_Jinkela_wire_9440),
        .b(new_Jinkela_wire_1391),
        .c(n_0788_)
    );

    and_ii n_2234_ (
        .a(new_Jinkela_wire_8479),
        .b(new_Jinkela_wire_3870),
        .c(n_0121_)
    );

    bfr new_Jinkela_buffer_2939 (
        .din(new_Jinkela_wire_3364),
        .dout(new_Jinkela_wire_3365)
    );

    and_ii n_1521_ (
        .a(new_Jinkela_wire_187),
        .b(new_Jinkela_wire_771),
        .c(n_0789_)
    );

    and_bi n_2235_ (
        .a(new_Jinkela_wire_5729),
        .b(new_Jinkela_wire_7991),
        .c(n_0122_)
    );

    bfr new_Jinkela_buffer_2839 (
        .din(new_Jinkela_wire_3258),
        .dout(new_Jinkela_wire_3259)
    );

    and_bb n_1522_ (
        .a(new_Jinkela_wire_186),
        .b(new_Jinkela_wire_770),
        .c(n_0790_)
    );

    and_bi n_2236_ (
        .a(new_Jinkela_wire_7990),
        .b(new_Jinkela_wire_5728),
        .c(n_0123_)
    );

    bfr new_Jinkela_buffer_2876 (
        .din(new_Jinkela_wire_3299),
        .dout(new_Jinkela_wire_3300)
    );

    or_bb n_1523_ (
        .a(n_0790_),
        .b(n_0789_),
        .c(n_0791_)
    );

    or_bb n_2237_ (
        .a(n_0123_),
        .b(n_0122_),
        .c(new_net_2556)
    );

    bfr new_Jinkela_buffer_2840 (
        .din(new_Jinkela_wire_3259),
        .dout(new_Jinkela_wire_3260)
    );

    and_ii n_1524_ (
        .a(new_Jinkela_wire_6397),
        .b(new_Jinkela_wire_6263),
        .c(n_0792_)
    );

    or_bi n_2238_ (
        .a(new_Jinkela_wire_5876),
        .b(new_Jinkela_wire_6237),
        .c(n_0124_)
    );

    and_bb n_1525_ (
        .a(new_Jinkela_wire_9389),
        .b(new_Jinkela_wire_8174),
        .c(n_0793_)
    );

    and_bi n_2239_ (
        .a(new_Jinkela_wire_9156),
        .b(new_Jinkela_wire_9702),
        .c(n_0125_)
    );

    bfr new_Jinkela_buffer_2841 (
        .din(new_Jinkela_wire_3260),
        .dout(new_Jinkela_wire_3261)
    );

    and_ii n_1526_ (
        .a(new_Jinkela_wire_9388),
        .b(new_Jinkela_wire_8173),
        .c(n_0794_)
    );

    and_bi n_2240_ (
        .a(new_Jinkela_wire_9701),
        .b(new_Jinkela_wire_9155),
        .c(n_0126_)
    );

    bfr new_Jinkela_buffer_7027 (
        .din(new_Jinkela_wire_8679),
        .dout(new_Jinkela_wire_8680)
    );

    bfr new_Jinkela_buffer_1210 (
        .din(new_Jinkela_wire_1526),
        .dout(new_Jinkela_wire_1527)
    );

    bfr new_Jinkela_buffer_5377 (
        .din(new_Jinkela_wire_6456),
        .dout(new_Jinkela_wire_6457)
    );

    bfr new_Jinkela_buffer_7052 (
        .din(new_Jinkela_wire_8712),
        .dout(new_Jinkela_wire_8713)
    );

    bfr new_Jinkela_buffer_1248 (
        .din(new_Jinkela_wire_1568),
        .dout(new_Jinkela_wire_1569)
    );

    spl2 new_Jinkela_splitter_420 (
        .a(new_Jinkela_wire_6521),
        .b(new_Jinkela_wire_6522),
        .c(new_Jinkela_wire_6523)
    );

    bfr new_Jinkela_buffer_7028 (
        .din(new_Jinkela_wire_8680),
        .dout(new_Jinkela_wire_8681)
    );

    bfr new_Jinkela_buffer_5415 (
        .din(new_Jinkela_wire_6494),
        .dout(new_Jinkela_wire_6495)
    );

    bfr new_Jinkela_buffer_1211 (
        .din(new_Jinkela_wire_1527),
        .dout(new_Jinkela_wire_1528)
    );

    bfr new_Jinkela_buffer_5378 (
        .din(new_Jinkela_wire_6457),
        .dout(new_Jinkela_wire_6458)
    );

    bfr new_Jinkela_buffer_7055 (
        .din(new_Jinkela_wire_8719),
        .dout(new_Jinkela_wire_8720)
    );

    bfr new_Jinkela_buffer_1373 (
        .din(N163),
        .dout(new_Jinkela_wire_1699)
    );

    bfr new_Jinkela_buffer_7029 (
        .din(new_Jinkela_wire_8681),
        .dout(new_Jinkela_wire_8682)
    );

    bfr new_Jinkela_buffer_1212 (
        .din(new_Jinkela_wire_1528),
        .dout(new_Jinkela_wire_1529)
    );

    bfr new_Jinkela_buffer_5379 (
        .din(new_Jinkela_wire_6458),
        .dout(new_Jinkela_wire_6459)
    );

    bfr new_Jinkela_buffer_7053 (
        .din(new_Jinkela_wire_8713),
        .dout(new_Jinkela_wire_8714)
    );

    bfr new_Jinkela_buffer_1249 (
        .din(new_Jinkela_wire_1569),
        .dout(new_Jinkela_wire_1570)
    );

    bfr new_Jinkela_buffer_7030 (
        .din(new_Jinkela_wire_8682),
        .dout(new_Jinkela_wire_8683)
    );

    bfr new_Jinkela_buffer_5416 (
        .din(new_Jinkela_wire_6495),
        .dout(new_Jinkela_wire_6496)
    );

    bfr new_Jinkela_buffer_1213 (
        .din(new_Jinkela_wire_1529),
        .dout(new_Jinkela_wire_1530)
    );

    bfr new_Jinkela_buffer_5380 (
        .din(new_Jinkela_wire_6459),
        .dout(new_Jinkela_wire_6460)
    );

    bfr new_Jinkela_buffer_1302 (
        .din(new_Jinkela_wire_1627),
        .dout(new_Jinkela_wire_1628)
    );

    spl4L new_Jinkela_splitter_671 (
        .a(n_0909_),
        .d(new_Jinkela_wire_8763),
        .b(new_Jinkela_wire_8764),
        .e(new_Jinkela_wire_8765),
        .c(new_Jinkela_wire_8766)
    );

    bfr new_Jinkela_buffer_7031 (
        .din(new_Jinkela_wire_8683),
        .dout(new_Jinkela_wire_8684)
    );

    bfr new_Jinkela_buffer_5442 (
        .din(n_0503_),
        .dout(new_Jinkela_wire_6536)
    );

    bfr new_Jinkela_buffer_1214 (
        .din(new_Jinkela_wire_1530),
        .dout(new_Jinkela_wire_1531)
    );

    bfr new_Jinkela_buffer_5381 (
        .din(new_Jinkela_wire_6460),
        .dout(new_Jinkela_wire_6461)
    );

    bfr new_Jinkela_buffer_7056 (
        .din(new_Jinkela_wire_8720),
        .dout(new_Jinkela_wire_8721)
    );

    bfr new_Jinkela_buffer_1250 (
        .din(new_Jinkela_wire_1570),
        .dout(new_Jinkela_wire_1571)
    );

    bfr new_Jinkela_buffer_7032 (
        .din(new_Jinkela_wire_8684),
        .dout(new_Jinkela_wire_8685)
    );

    bfr new_Jinkela_buffer_5417 (
        .din(new_Jinkela_wire_6496),
        .dout(new_Jinkela_wire_6497)
    );

    bfr new_Jinkela_buffer_1215 (
        .din(new_Jinkela_wire_1531),
        .dout(new_Jinkela_wire_1532)
    );

    bfr new_Jinkela_buffer_5382 (
        .din(new_Jinkela_wire_6461),
        .dout(new_Jinkela_wire_6462)
    );

    spl2 new_Jinkela_splitter_668 (
        .a(n_0685_),
        .b(new_Jinkela_wire_8754),
        .c(new_Jinkela_wire_8755)
    );

    bfr new_Jinkela_buffer_1367 (
        .din(new_Jinkela_wire_1692),
        .dout(new_Jinkela_wire_1693)
    );

    bfr new_Jinkela_buffer_7033 (
        .din(new_Jinkela_wire_8685),
        .dout(new_Jinkela_wire_8686)
    );

    bfr new_Jinkela_buffer_5438 (
        .din(new_Jinkela_wire_6525),
        .dout(new_Jinkela_wire_6526)
    );

    bfr new_Jinkela_buffer_1216 (
        .din(new_Jinkela_wire_1532),
        .dout(new_Jinkela_wire_1533)
    );

    bfr new_Jinkela_buffer_5383 (
        .din(new_Jinkela_wire_6462),
        .dout(new_Jinkela_wire_6463)
    );

    bfr new_Jinkela_buffer_7057 (
        .din(new_Jinkela_wire_8721),
        .dout(new_Jinkela_wire_8722)
    );

    bfr new_Jinkela_buffer_1251 (
        .din(new_Jinkela_wire_1571),
        .dout(new_Jinkela_wire_1572)
    );

    bfr new_Jinkela_buffer_7034 (
        .din(new_Jinkela_wire_8686),
        .dout(new_Jinkela_wire_8687)
    );

    bfr new_Jinkela_buffer_5418 (
        .din(new_Jinkela_wire_6497),
        .dout(new_Jinkela_wire_6498)
    );

    bfr new_Jinkela_buffer_1217 (
        .din(new_Jinkela_wire_1533),
        .dout(new_Jinkela_wire_1534)
    );

    bfr new_Jinkela_buffer_5384 (
        .din(new_Jinkela_wire_6463),
        .dout(new_Jinkela_wire_6464)
    );

    bfr new_Jinkela_buffer_7082 (
        .din(n_0879_),
        .dout(new_Jinkela_wire_8753)
    );

    bfr new_Jinkela_buffer_1303 (
        .din(new_Jinkela_wire_1628),
        .dout(new_Jinkela_wire_1629)
    );

    bfr new_Jinkela_buffer_7035 (
        .din(new_Jinkela_wire_8687),
        .dout(new_Jinkela_wire_8688)
    );

    bfr new_Jinkela_buffer_5439 (
        .din(new_Jinkela_wire_6526),
        .dout(new_Jinkela_wire_6527)
    );

    bfr new_Jinkela_buffer_1218 (
        .din(new_Jinkela_wire_1534),
        .dout(new_Jinkela_wire_1535)
    );

    bfr new_Jinkela_buffer_5385 (
        .din(new_Jinkela_wire_6464),
        .dout(new_Jinkela_wire_6465)
    );

    bfr new_Jinkela_buffer_7058 (
        .din(new_Jinkela_wire_8722),
        .dout(new_Jinkela_wire_8723)
    );

    bfr new_Jinkela_buffer_1252 (
        .din(new_Jinkela_wire_1572),
        .dout(new_Jinkela_wire_1573)
    );

    bfr new_Jinkela_buffer_7036 (
        .din(new_Jinkela_wire_8688),
        .dout(new_Jinkela_wire_8689)
    );

    bfr new_Jinkela_buffer_5419 (
        .din(new_Jinkela_wire_6498),
        .dout(new_Jinkela_wire_6499)
    );

    bfr new_Jinkela_buffer_1219 (
        .din(new_Jinkela_wire_1535),
        .dout(new_Jinkela_wire_1536)
    );

    bfr new_Jinkela_buffer_5386 (
        .din(new_Jinkela_wire_6465),
        .dout(new_Jinkela_wire_6466)
    );

    bfr new_Jinkela_buffer_1370 (
        .din(new_Jinkela_wire_1695),
        .dout(new_Jinkela_wire_1696)
    );

    bfr new_Jinkela_buffer_7083 (
        .din(n_0562_),
        .dout(new_Jinkela_wire_8756)
    );

    bfr new_Jinkela_buffer_7037 (
        .din(new_Jinkela_wire_8689),
        .dout(new_Jinkela_wire_8690)
    );

    spl2 new_Jinkela_splitter_423 (
        .a(n_1302_),
        .b(new_Jinkela_wire_6534),
        .c(new_Jinkela_wire_6535)
    );

    bfr new_Jinkela_buffer_1220 (
        .din(new_Jinkela_wire_1536),
        .dout(new_Jinkela_wire_1537)
    );

    bfr new_Jinkela_buffer_5387 (
        .din(new_Jinkela_wire_6466),
        .dout(new_Jinkela_wire_6467)
    );

    bfr new_Jinkela_buffer_7059 (
        .din(new_Jinkela_wire_8723),
        .dout(new_Jinkela_wire_8724)
    );

    bfr new_Jinkela_buffer_1253 (
        .din(new_Jinkela_wire_1573),
        .dout(new_Jinkela_wire_1574)
    );

    bfr new_Jinkela_buffer_5441 (
        .din(new_Jinkela_wire_6530),
        .dout(new_Jinkela_wire_6531)
    );

    bfr new_Jinkela_buffer_7038 (
        .din(new_Jinkela_wire_8690),
        .dout(new_Jinkela_wire_8691)
    );

    bfr new_Jinkela_buffer_5420 (
        .din(new_Jinkela_wire_6499),
        .dout(new_Jinkela_wire_6500)
    );

    bfr new_Jinkela_buffer_1221 (
        .din(new_Jinkela_wire_1537),
        .dout(new_Jinkela_wire_1538)
    );

    bfr new_Jinkela_buffer_5388 (
        .din(new_Jinkela_wire_6467),
        .dout(new_Jinkela_wire_6468)
    );

    bfr new_Jinkela_buffer_7084 (
        .din(new_Jinkela_wire_8756),
        .dout(new_Jinkela_wire_8757)
    );

    bfr new_Jinkela_buffer_1304 (
        .din(new_Jinkela_wire_1629),
        .dout(new_Jinkela_wire_1630)
    );

    bfr new_Jinkela_buffer_7039 (
        .din(new_Jinkela_wire_8691),
        .dout(new_Jinkela_wire_8692)
    );

    bfr new_Jinkela_buffer_5443 (
        .din(n_1357_),
        .dout(new_Jinkela_wire_6541)
    );

    bfr new_Jinkela_buffer_1222 (
        .din(new_Jinkela_wire_1538),
        .dout(new_Jinkela_wire_1539)
    );

    bfr new_Jinkela_buffer_5389 (
        .din(new_Jinkela_wire_6468),
        .dout(new_Jinkela_wire_6469)
    );

    bfr new_Jinkela_buffer_7060 (
        .din(new_Jinkela_wire_8724),
        .dout(new_Jinkela_wire_8725)
    );

    bfr new_Jinkela_buffer_1254 (
        .din(new_Jinkela_wire_1574),
        .dout(new_Jinkela_wire_1575)
    );

    bfr new_Jinkela_buffer_7040 (
        .din(new_Jinkela_wire_8692),
        .dout(new_Jinkela_wire_8693)
    );

    bfr new_Jinkela_buffer_5421 (
        .din(new_Jinkela_wire_6500),
        .dout(new_Jinkela_wire_6501)
    );

    bfr new_Jinkela_buffer_1223 (
        .din(new_Jinkela_wire_1539),
        .dout(new_Jinkela_wire_1540)
    );

    bfr new_Jinkela_buffer_5390 (
        .din(new_Jinkela_wire_6469),
        .dout(new_Jinkela_wire_6470)
    );

    spl3L new_Jinkela_splitter_669 (
        .a(n_1325_),
        .d(new_Jinkela_wire_8758),
        .b(new_Jinkela_wire_8759),
        .c(new_Jinkela_wire_8760)
    );

    bfr new_Jinkela_buffer_1368 (
        .din(new_Jinkela_wire_1693),
        .dout(new_Jinkela_wire_1694)
    );

    bfr new_Jinkela_buffer_7041 (
        .din(new_Jinkela_wire_8693),
        .dout(new_Jinkela_wire_8694)
    );

    bfr new_Jinkela_buffer_1255 (
        .din(new_Jinkela_wire_1575),
        .dout(new_Jinkela_wire_1576)
    );

    bfr new_Jinkela_buffer_5391 (
        .din(new_Jinkela_wire_6470),
        .dout(new_Jinkela_wire_6471)
    );

    bfr new_Jinkela_buffer_7061 (
        .din(new_Jinkela_wire_8725),
        .dout(new_Jinkela_wire_8726)
    );

    bfr new_Jinkela_buffer_1305 (
        .din(new_Jinkela_wire_1630),
        .dout(new_Jinkela_wire_1631)
    );

    spl2 new_Jinkela_splitter_422 (
        .a(new_Jinkela_wire_6531),
        .b(new_Jinkela_wire_6532),
        .c(new_Jinkela_wire_6533)
    );

    bfr new_Jinkela_buffer_7042 (
        .din(new_Jinkela_wire_8694),
        .dout(new_Jinkela_wire_8695)
    );

    bfr new_Jinkela_buffer_5422 (
        .din(new_Jinkela_wire_6501),
        .dout(new_Jinkela_wire_6502)
    );

    bfr new_Jinkela_buffer_1256 (
        .din(new_Jinkela_wire_1576),
        .dout(new_Jinkela_wire_1577)
    );

    bfr new_Jinkela_buffer_5392 (
        .din(new_Jinkela_wire_6471),
        .dout(new_Jinkela_wire_6472)
    );

    spl2 new_Jinkela_splitter_102 (
        .a(N165),
        .b(new_Jinkela_wire_1700),
        .c(new_Jinkela_wire_1701)
    );

    bfr new_Jinkela_buffer_1374 (
        .din(N217),
        .dout(new_Jinkela_wire_1702)
    );

    spl2 new_Jinkela_splitter_672 (
        .a(n_0026_),
        .b(new_Jinkela_wire_8767),
        .c(new_Jinkela_wire_8768)
    );

    spl2 new_Jinkela_splitter_660 (
        .a(new_Jinkela_wire_8695),
        .b(new_Jinkela_wire_8696),
        .c(new_Jinkela_wire_8697)
    );

    bfr new_Jinkela_buffer_1257 (
        .din(new_Jinkela_wire_1577),
        .dout(new_Jinkela_wire_1578)
    );

    bfr new_Jinkela_buffer_5393 (
        .din(new_Jinkela_wire_6472),
        .dout(new_Jinkela_wire_6473)
    );

    bfr new_Jinkela_buffer_1306 (
        .din(new_Jinkela_wire_1631),
        .dout(new_Jinkela_wire_1632)
    );

    bfr new_Jinkela_buffer_7085 (
        .din(new_Jinkela_wire_8768),
        .dout(new_Jinkela_wire_8769)
    );

    bfr new_Jinkela_buffer_7062 (
        .din(new_Jinkela_wire_8726),
        .dout(new_Jinkela_wire_8727)
    );

    bfr new_Jinkela_buffer_5423 (
        .din(new_Jinkela_wire_6502),
        .dout(new_Jinkela_wire_6503)
    );

    bfr new_Jinkela_buffer_1258 (
        .din(new_Jinkela_wire_1578),
        .dout(new_Jinkela_wire_1579)
    );

    bfr new_Jinkela_buffer_5394 (
        .din(new_Jinkela_wire_6473),
        .dout(new_Jinkela_wire_6474)
    );

    bfr new_Jinkela_buffer_7063 (
        .din(new_Jinkela_wire_8727),
        .dout(new_Jinkela_wire_8728)
    );

    bfr new_Jinkela_buffer_1371 (
        .din(new_Jinkela_wire_1696),
        .dout(new_Jinkela_wire_1697)
    );

    spl2 new_Jinkela_splitter_670 (
        .a(new_Jinkela_wire_8760),
        .b(new_Jinkela_wire_8761),
        .c(new_Jinkela_wire_8762)
    );

    bfr new_Jinkela_buffer_1259 (
        .din(new_Jinkela_wire_1579),
        .dout(new_Jinkela_wire_1580)
    );

    bfr new_Jinkela_buffer_5395 (
        .din(new_Jinkela_wire_6474),
        .dout(new_Jinkela_wire_6475)
    );

    bfr new_Jinkela_buffer_7127 (
        .din(n_0846_),
        .dout(new_Jinkela_wire_8820)
    );

    bfr new_Jinkela_buffer_7064 (
        .din(new_Jinkela_wire_8728),
        .dout(new_Jinkela_wire_8729)
    );

    bfr new_Jinkela_buffer_1307 (
        .din(new_Jinkela_wire_1632),
        .dout(new_Jinkela_wire_1633)
    );

    spl2 new_Jinkela_splitter_424 (
        .a(new_Jinkela_wire_6536),
        .b(new_Jinkela_wire_6537),
        .c(new_Jinkela_wire_6538)
    );

    bfr new_Jinkela_buffer_5424 (
        .din(new_Jinkela_wire_6503),
        .dout(new_Jinkela_wire_6504)
    );

    bfr new_Jinkela_buffer_1260 (
        .din(new_Jinkela_wire_1580),
        .dout(new_Jinkela_wire_1581)
    );

    bfr new_Jinkela_buffer_5396 (
        .din(new_Jinkela_wire_6475),
        .dout(new_Jinkela_wire_6476)
    );

    spl3L new_Jinkela_splitter_674 (
        .a(n_0686_),
        .d(new_Jinkela_wire_8812),
        .b(new_Jinkela_wire_8813),
        .c(new_Jinkela_wire_8814)
    );

    bfr new_Jinkela_buffer_7065 (
        .din(new_Jinkela_wire_8729),
        .dout(new_Jinkela_wire_8730)
    );

    spl2 new_Jinkela_splitter_425 (
        .a(n_0548_),
        .b(new_Jinkela_wire_6539),
        .c(new_Jinkela_wire_6540)
    );

    bfr new_Jinkela_buffer_1261 (
        .din(new_Jinkela_wire_1581),
        .dout(new_Jinkela_wire_1582)
    );

    bfr new_Jinkela_buffer_5397 (
        .din(new_Jinkela_wire_6476),
        .dout(new_Jinkela_wire_6477)
    );

    bfr new_Jinkela_buffer_7066 (
        .din(new_Jinkela_wire_8730),
        .dout(new_Jinkela_wire_8731)
    );

    bfr new_Jinkela_buffer_1308 (
        .din(new_Jinkela_wire_1633),
        .dout(new_Jinkela_wire_1634)
    );

    bfr new_Jinkela_buffer_6205 (
        .din(new_Jinkela_wire_7578),
        .dout(new_Jinkela_wire_7579)
    );

    bfr new_Jinkela_buffer_6282 (
        .din(new_Jinkela_wire_7659),
        .dout(new_Jinkela_wire_7660)
    );

    bfr new_Jinkela_buffer_6206 (
        .din(new_Jinkela_wire_7579),
        .dout(new_Jinkela_wire_7580)
    );

    bfr new_Jinkela_buffer_6229 (
        .din(new_Jinkela_wire_7602),
        .dout(new_Jinkela_wire_7603)
    );

    bfr new_Jinkela_buffer_6207 (
        .din(new_Jinkela_wire_7580),
        .dout(new_Jinkela_wire_7581)
    );

    bfr new_Jinkela_buffer_6308 (
        .din(new_Jinkela_wire_7689),
        .dout(new_Jinkela_wire_7690)
    );

    bfr new_Jinkela_buffer_6208 (
        .din(new_Jinkela_wire_7581),
        .dout(new_Jinkela_wire_7582)
    );

    bfr new_Jinkela_buffer_6230 (
        .din(new_Jinkela_wire_7603),
        .dout(new_Jinkela_wire_7604)
    );

    bfr new_Jinkela_buffer_6209 (
        .din(new_Jinkela_wire_7582),
        .dout(new_Jinkela_wire_7583)
    );

    bfr new_Jinkela_buffer_6283 (
        .din(new_Jinkela_wire_7660),
        .dout(new_Jinkela_wire_7661)
    );

    bfr new_Jinkela_buffer_6210 (
        .din(new_Jinkela_wire_7583),
        .dout(new_Jinkela_wire_7584)
    );

    bfr new_Jinkela_buffer_6231 (
        .din(new_Jinkela_wire_7604),
        .dout(new_Jinkela_wire_7605)
    );

    bfr new_Jinkela_buffer_6211 (
        .din(new_Jinkela_wire_7584),
        .dout(new_Jinkela_wire_7585)
    );

    bfr new_Jinkela_buffer_6346 (
        .din(new_Jinkela_wire_7731),
        .dout(new_Jinkela_wire_7732)
    );

    bfr new_Jinkela_buffer_6232 (
        .din(new_Jinkela_wire_7605),
        .dout(new_Jinkela_wire_7606)
    );

    bfr new_Jinkela_buffer_6284 (
        .din(new_Jinkela_wire_7661),
        .dout(new_Jinkela_wire_7662)
    );

    bfr new_Jinkela_buffer_6233 (
        .din(new_Jinkela_wire_7606),
        .dout(new_Jinkela_wire_7607)
    );

    bfr new_Jinkela_buffer_6309 (
        .din(new_Jinkela_wire_7690),
        .dout(new_Jinkela_wire_7691)
    );

    bfr new_Jinkela_buffer_6234 (
        .din(new_Jinkela_wire_7607),
        .dout(new_Jinkela_wire_7608)
    );

    bfr new_Jinkela_buffer_6285 (
        .din(new_Jinkela_wire_7662),
        .dout(new_Jinkela_wire_7663)
    );

    bfr new_Jinkela_buffer_6235 (
        .din(new_Jinkela_wire_7608),
        .dout(new_Jinkela_wire_7609)
    );

    bfr new_Jinkela_buffer_6236 (
        .din(new_Jinkela_wire_7609),
        .dout(new_Jinkela_wire_7610)
    );

    bfr new_Jinkela_buffer_6286 (
        .din(new_Jinkela_wire_7663),
        .dout(new_Jinkela_wire_7664)
    );

    bfr new_Jinkela_buffer_6237 (
        .din(new_Jinkela_wire_7610),
        .dout(new_Jinkela_wire_7611)
    );

    bfr new_Jinkela_buffer_6310 (
        .din(new_Jinkela_wire_7691),
        .dout(new_Jinkela_wire_7692)
    );

    bfr new_Jinkela_buffer_6238 (
        .din(new_Jinkela_wire_7611),
        .dout(new_Jinkela_wire_7612)
    );

    bfr new_Jinkela_buffer_6287 (
        .din(new_Jinkela_wire_7664),
        .dout(new_Jinkela_wire_7665)
    );

    bfr new_Jinkela_buffer_6239 (
        .din(new_Jinkela_wire_7612),
        .dout(new_Jinkela_wire_7613)
    );

    spl4L new_Jinkela_splitter_549 (
        .a(n_0691_),
        .d(new_Jinkela_wire_7747),
        .b(new_Jinkela_wire_7748),
        .e(new_Jinkela_wire_7749),
        .c(new_Jinkela_wire_7750)
    );

    bfr new_Jinkela_buffer_6240 (
        .din(new_Jinkela_wire_7613),
        .dout(new_Jinkela_wire_7614)
    );

    bfr new_Jinkela_buffer_6288 (
        .din(new_Jinkela_wire_7665),
        .dout(new_Jinkela_wire_7666)
    );

    bfr new_Jinkela_buffer_6241 (
        .din(new_Jinkela_wire_7614),
        .dout(new_Jinkela_wire_7615)
    );

    bfr new_Jinkela_buffer_6311 (
        .din(new_Jinkela_wire_7692),
        .dout(new_Jinkela_wire_7693)
    );

    bfr new_Jinkela_buffer_6242 (
        .din(new_Jinkela_wire_7615),
        .dout(new_Jinkela_wire_7616)
    );

    bfr new_Jinkela_buffer_6289 (
        .din(new_Jinkela_wire_7666),
        .dout(new_Jinkela_wire_7667)
    );

    bfr new_Jinkela_buffer_6243 (
        .din(new_Jinkela_wire_7616),
        .dout(new_Jinkela_wire_7617)
    );

    bfr new_Jinkela_buffer_6347 (
        .din(new_Jinkela_wire_7732),
        .dout(new_Jinkela_wire_7733)
    );

    bfr new_Jinkela_buffer_6244 (
        .din(new_Jinkela_wire_7617),
        .dout(new_Jinkela_wire_7618)
    );

    bfr new_Jinkela_buffer_6290 (
        .din(new_Jinkela_wire_7667),
        .dout(new_Jinkela_wire_7668)
    );

    bfr new_Jinkela_buffer_6245 (
        .din(new_Jinkela_wire_7618),
        .dout(new_Jinkela_wire_7619)
    );

    bfr new_Jinkela_buffer_6312 (
        .din(new_Jinkela_wire_7693),
        .dout(new_Jinkela_wire_7694)
    );

    spl2 new_Jinkela_splitter_25 (
        .a(N361),
        .b(new_Jinkela_wire_800),
        .c(new_Jinkela_wire_801)
    );

    bfr new_Jinkela_buffer_807 (
        .din(N195),
        .dout(new_Jinkela_wire_868)
    );

    bfr new_Jinkela_buffer_3730 (
        .din(new_Jinkela_wire_4350),
        .dout(new_Jinkela_wire_4351)
    );

    bfr new_Jinkela_buffer_8266 (
        .din(new_Jinkela_wire_10380),
        .dout(new_Jinkela_wire_10381)
    );

    bfr new_Jinkela_buffer_8166 (
        .din(new_Jinkela_wire_10267),
        .dout(new_Jinkela_wire_10268)
    );

    bfr new_Jinkela_buffer_674 (
        .din(new_Jinkela_wire_726),
        .dout(new_Jinkela_wire_727)
    );

    bfr new_Jinkela_buffer_3717 (
        .din(new_Jinkela_wire_4335),
        .dout(new_Jinkela_wire_4336)
    );

    bfr new_Jinkela_buffer_8210 (
        .din(new_Jinkela_wire_10313),
        .dout(new_Jinkela_wire_10314)
    );

    bfr new_Jinkela_buffer_737 (
        .din(new_Jinkela_wire_793),
        .dout(new_Jinkela_wire_794)
    );

    bfr new_Jinkela_buffer_8167 (
        .din(new_Jinkela_wire_10268),
        .dout(new_Jinkela_wire_10269)
    );

    bfr new_Jinkela_buffer_3791 (
        .din(new_Jinkela_wire_4413),
        .dout(new_Jinkela_wire_4414)
    );

    bfr new_Jinkela_buffer_675 (
        .din(new_Jinkela_wire_727),
        .dout(new_Jinkela_wire_728)
    );

    bfr new_Jinkela_buffer_3731 (
        .din(new_Jinkela_wire_4351),
        .dout(new_Jinkela_wire_4352)
    );

    bfr new_Jinkela_buffer_8258 (
        .din(new_Jinkela_wire_10370),
        .dout(new_Jinkela_wire_10371)
    );

    bfr new_Jinkela_buffer_740 (
        .din(new_Jinkela_wire_796),
        .dout(new_Jinkela_wire_797)
    );

    bfr new_Jinkela_buffer_8248 (
        .din(new_Jinkela_wire_10351),
        .dout(new_Jinkela_wire_10352)
    );

    bfr new_Jinkela_buffer_8168 (
        .din(new_Jinkela_wire_10269),
        .dout(new_Jinkela_wire_10270)
    );

    bfr new_Jinkela_buffer_3778 (
        .din(new_Jinkela_wire_4400),
        .dout(new_Jinkela_wire_4401)
    );

    bfr new_Jinkela_buffer_676 (
        .din(new_Jinkela_wire_728),
        .dout(new_Jinkela_wire_729)
    );

    bfr new_Jinkela_buffer_3732 (
        .din(new_Jinkela_wire_4352),
        .dout(new_Jinkela_wire_4353)
    );

    bfr new_Jinkela_buffer_8211 (
        .din(new_Jinkela_wire_10314),
        .dout(new_Jinkela_wire_10315)
    );

    bfr new_Jinkela_buffer_738 (
        .din(new_Jinkela_wire_794),
        .dout(new_Jinkela_wire_795)
    );

    bfr new_Jinkela_buffer_8169 (
        .din(new_Jinkela_wire_10270),
        .dout(new_Jinkela_wire_10271)
    );

    bfr new_Jinkela_buffer_677 (
        .din(new_Jinkela_wire_729),
        .dout(new_Jinkela_wire_730)
    );

    bfr new_Jinkela_buffer_3733 (
        .din(new_Jinkela_wire_4353),
        .dout(new_Jinkela_wire_4354)
    );

    bfr new_Jinkela_buffer_808 (
        .din(new_Jinkela_wire_868),
        .dout(new_Jinkela_wire_869)
    );

    bfr new_Jinkela_buffer_3807 (
        .din(new_Jinkela_wire_4436),
        .dout(new_Jinkela_wire_4437)
    );

    bfr new_Jinkela_buffer_8170 (
        .din(new_Jinkela_wire_10271),
        .dout(new_Jinkela_wire_10272)
    );

    bfr new_Jinkela_buffer_3779 (
        .din(new_Jinkela_wire_4401),
        .dout(new_Jinkela_wire_4402)
    );

    bfr new_Jinkela_buffer_678 (
        .din(new_Jinkela_wire_730),
        .dout(new_Jinkela_wire_731)
    );

    bfr new_Jinkela_buffer_3734 (
        .din(new_Jinkela_wire_4354),
        .dout(new_Jinkela_wire_4355)
    );

    bfr new_Jinkela_buffer_8212 (
        .din(new_Jinkela_wire_10315),
        .dout(new_Jinkela_wire_10316)
    );

    bfr new_Jinkela_buffer_741 (
        .din(new_Jinkela_wire_797),
        .dout(new_Jinkela_wire_798)
    );

    bfr new_Jinkela_buffer_8171 (
        .din(new_Jinkela_wire_10272),
        .dout(new_Jinkela_wire_10273)
    );

    bfr new_Jinkela_buffer_3792 (
        .din(new_Jinkela_wire_4414),
        .dout(new_Jinkela_wire_4415)
    );

    bfr new_Jinkela_buffer_679 (
        .din(new_Jinkela_wire_731),
        .dout(new_Jinkela_wire_732)
    );

    bfr new_Jinkela_buffer_3735 (
        .din(new_Jinkela_wire_4355),
        .dout(new_Jinkela_wire_4356)
    );

    bfr new_Jinkela_buffer_811 (
        .din(N231),
        .dout(new_Jinkela_wire_872)
    );

    bfr new_Jinkela_buffer_8249 (
        .din(new_Jinkela_wire_10352),
        .dout(new_Jinkela_wire_10353)
    );

    bfr new_Jinkela_buffer_8172 (
        .din(new_Jinkela_wire_10273),
        .dout(new_Jinkela_wire_10274)
    );

    bfr new_Jinkela_buffer_3780 (
        .din(new_Jinkela_wire_4402),
        .dout(new_Jinkela_wire_4403)
    );

    bfr new_Jinkela_buffer_680 (
        .din(new_Jinkela_wire_732),
        .dout(new_Jinkela_wire_733)
    );

    bfr new_Jinkela_buffer_3736 (
        .din(new_Jinkela_wire_4356),
        .dout(new_Jinkela_wire_4357)
    );

    bfr new_Jinkela_buffer_8213 (
        .din(new_Jinkela_wire_10316),
        .dout(new_Jinkela_wire_10317)
    );

    bfr new_Jinkela_buffer_742 (
        .din(new_Jinkela_wire_798),
        .dout(new_Jinkela_wire_799)
    );

    bfr new_Jinkela_buffer_8173 (
        .din(new_Jinkela_wire_10274),
        .dout(new_Jinkela_wire_10275)
    );

    bfr new_Jinkela_buffer_681 (
        .din(new_Jinkela_wire_733),
        .dout(new_Jinkela_wire_734)
    );

    bfr new_Jinkela_buffer_3737 (
        .din(new_Jinkela_wire_4357),
        .dout(new_Jinkela_wire_4358)
    );

    bfr new_Jinkela_buffer_743 (
        .din(new_Jinkela_wire_801),
        .dout(new_Jinkela_wire_802)
    );

    spl2 new_Jinkela_splitter_225 (
        .a(new_Jinkela_wire_4429),
        .b(new_Jinkela_wire_4430),
        .c(new_Jinkela_wire_4431)
    );

    bfr new_Jinkela_buffer_8174 (
        .din(new_Jinkela_wire_10275),
        .dout(new_Jinkela_wire_10276)
    );

    bfr new_Jinkela_buffer_3781 (
        .din(new_Jinkela_wire_4403),
        .dout(new_Jinkela_wire_4404)
    );

    bfr new_Jinkela_buffer_682 (
        .din(new_Jinkela_wire_734),
        .dout(new_Jinkela_wire_735)
    );

    bfr new_Jinkela_buffer_3738 (
        .din(new_Jinkela_wire_4358),
        .dout(new_Jinkela_wire_4359)
    );

    bfr new_Jinkela_buffer_8214 (
        .din(new_Jinkela_wire_10317),
        .dout(new_Jinkela_wire_10318)
    );

    bfr new_Jinkela_buffer_8175 (
        .din(new_Jinkela_wire_10276),
        .dout(new_Jinkela_wire_10277)
    );

    bfr new_Jinkela_buffer_3793 (
        .din(new_Jinkela_wire_4415),
        .dout(new_Jinkela_wire_4416)
    );

    bfr new_Jinkela_buffer_683 (
        .din(new_Jinkela_wire_735),
        .dout(new_Jinkela_wire_736)
    );

    bfr new_Jinkela_buffer_3739 (
        .din(new_Jinkela_wire_4359),
        .dout(new_Jinkela_wire_4360)
    );

    bfr new_Jinkela_buffer_8259 (
        .din(new_Jinkela_wire_10371),
        .dout(new_Jinkela_wire_10372)
    );

    bfr new_Jinkela_buffer_744 (
        .din(new_Jinkela_wire_802),
        .dout(new_Jinkela_wire_803)
    );

    bfr new_Jinkela_buffer_8250 (
        .din(new_Jinkela_wire_10353),
        .dout(new_Jinkela_wire_10354)
    );

    bfr new_Jinkela_buffer_8176 (
        .din(new_Jinkela_wire_10277),
        .dout(new_Jinkela_wire_10278)
    );

    bfr new_Jinkela_buffer_3782 (
        .din(new_Jinkela_wire_4404),
        .dout(new_Jinkela_wire_4405)
    );

    bfr new_Jinkela_buffer_684 (
        .din(new_Jinkela_wire_736),
        .dout(new_Jinkela_wire_737)
    );

    bfr new_Jinkela_buffer_3740 (
        .din(new_Jinkela_wire_4360),
        .dout(new_Jinkela_wire_4361)
    );

    bfr new_Jinkela_buffer_8215 (
        .din(new_Jinkela_wire_10318),
        .dout(new_Jinkela_wire_10319)
    );

    bfr new_Jinkela_buffer_815 (
        .din(N124),
        .dout(new_Jinkela_wire_876)
    );

    bfr new_Jinkela_buffer_8177 (
        .din(new_Jinkela_wire_10278),
        .dout(new_Jinkela_wire_10279)
    );

    bfr new_Jinkela_buffer_685 (
        .din(new_Jinkela_wire_737),
        .dout(new_Jinkela_wire_738)
    );

    bfr new_Jinkela_buffer_3741 (
        .din(new_Jinkela_wire_4361),
        .dout(new_Jinkela_wire_4362)
    );

    spl2 new_Jinkela_splitter_26 (
        .a(new_Jinkela_wire_803),
        .b(new_Jinkela_wire_804),
        .c(new_Jinkela_wire_805)
    );

    bfr new_Jinkela_buffer_8178 (
        .din(new_Jinkela_wire_10279),
        .dout(new_Jinkela_wire_10280)
    );

    bfr new_Jinkela_buffer_3783 (
        .din(new_Jinkela_wire_4405),
        .dout(new_Jinkela_wire_4406)
    );

    bfr new_Jinkela_buffer_686 (
        .din(new_Jinkela_wire_738),
        .dout(new_Jinkela_wire_739)
    );

    bfr new_Jinkela_buffer_3742 (
        .din(new_Jinkela_wire_4362),
        .dout(new_Jinkela_wire_4363)
    );

    bfr new_Jinkela_buffer_8216 (
        .din(new_Jinkela_wire_10319),
        .dout(new_Jinkela_wire_10320)
    );

    bfr new_Jinkela_buffer_745 (
        .din(new_Jinkela_wire_805),
        .dout(new_Jinkela_wire_806)
    );

    bfr new_Jinkela_buffer_8179 (
        .din(new_Jinkela_wire_10280),
        .dout(new_Jinkela_wire_10281)
    );

    bfr new_Jinkela_buffer_3794 (
        .din(new_Jinkela_wire_4416),
        .dout(new_Jinkela_wire_4417)
    );

    bfr new_Jinkela_buffer_687 (
        .din(new_Jinkela_wire_739),
        .dout(new_Jinkela_wire_740)
    );

    bfr new_Jinkela_buffer_3743 (
        .din(new_Jinkela_wire_4363),
        .dout(new_Jinkela_wire_4364)
    );

    bfr new_Jinkela_buffer_8267 (
        .din(n_0187_),
        .dout(new_Jinkela_wire_10386)
    );

    bfr new_Jinkela_buffer_809 (
        .din(new_Jinkela_wire_869),
        .dout(new_Jinkela_wire_870)
    );

    bfr new_Jinkela_buffer_8251 (
        .din(new_Jinkela_wire_10354),
        .dout(new_Jinkela_wire_10355)
    );

    bfr new_Jinkela_buffer_8180 (
        .din(new_Jinkela_wire_10281),
        .dout(new_Jinkela_wire_10282)
    );

    bfr new_Jinkela_buffer_3784 (
        .din(new_Jinkela_wire_4406),
        .dout(new_Jinkela_wire_4407)
    );

    bfr new_Jinkela_buffer_688 (
        .din(new_Jinkela_wire_740),
        .dout(new_Jinkela_wire_741)
    );

    bfr new_Jinkela_buffer_3744 (
        .din(new_Jinkela_wire_4364),
        .dout(new_Jinkela_wire_4365)
    );

    bfr new_Jinkela_buffer_8217 (
        .din(new_Jinkela_wire_10320),
        .dout(new_Jinkela_wire_10321)
    );

    bfr new_Jinkela_buffer_812 (
        .din(new_Jinkela_wire_872),
        .dout(new_Jinkela_wire_873)
    );

    bfr new_Jinkela_buffer_8181 (
        .din(new_Jinkela_wire_10282),
        .dout(new_Jinkela_wire_10283)
    );

    spl4L new_Jinkela_splitter_228 (
        .a(n_0031_),
        .d(new_Jinkela_wire_4438),
        .b(new_Jinkela_wire_4439),
        .e(new_Jinkela_wire_4440),
        .c(new_Jinkela_wire_4441)
    );

    bfr new_Jinkela_buffer_689 (
        .din(new_Jinkela_wire_741),
        .dout(new_Jinkela_wire_742)
    );

    bfr new_Jinkela_buffer_3745 (
        .din(new_Jinkela_wire_4365),
        .dout(new_Jinkela_wire_4366)
    );

    bfr new_Jinkela_buffer_746 (
        .din(new_Jinkela_wire_806),
        .dout(new_Jinkela_wire_807)
    );

    bfr new_Jinkela_buffer_8182 (
        .din(new_Jinkela_wire_10283),
        .dout(new_Jinkela_wire_10284)
    );

    bfr new_Jinkela_buffer_3785 (
        .din(new_Jinkela_wire_4407),
        .dout(new_Jinkela_wire_4408)
    );

    bfr new_Jinkela_buffer_690 (
        .din(new_Jinkela_wire_742),
        .dout(new_Jinkela_wire_743)
    );

    bfr new_Jinkela_buffer_3746 (
        .din(new_Jinkela_wire_4366),
        .dout(new_Jinkela_wire_4367)
    );

    bfr new_Jinkela_buffer_8218 (
        .din(new_Jinkela_wire_10321),
        .dout(new_Jinkela_wire_10322)
    );

    bfr new_Jinkela_buffer_810 (
        .din(new_Jinkela_wire_870),
        .dout(new_Jinkela_wire_871)
    );

    bfr new_Jinkela_buffer_8183 (
        .din(new_Jinkela_wire_10284),
        .dout(new_Jinkela_wire_10285)
    );

    bfr new_Jinkela_buffer_3795 (
        .din(new_Jinkela_wire_4417),
        .dout(new_Jinkela_wire_4418)
    );

    bfr new_Jinkela_buffer_691 (
        .din(new_Jinkela_wire_743),
        .dout(new_Jinkela_wire_744)
    );

    bfr new_Jinkela_buffer_3747 (
        .din(new_Jinkela_wire_4367),
        .dout(new_Jinkela_wire_4368)
    );

    bfr new_Jinkela_buffer_8260 (
        .din(new_Jinkela_wire_10372),
        .dout(new_Jinkela_wire_10373)
    );

    bfr new_Jinkela_buffer_747 (
        .din(new_Jinkela_wire_807),
        .dout(new_Jinkela_wire_808)
    );

    bfr new_Jinkela_buffer_8252 (
        .din(new_Jinkela_wire_10355),
        .dout(new_Jinkela_wire_10356)
    );

    bfr new_Jinkela_buffer_8184 (
        .din(new_Jinkela_wire_10285),
        .dout(new_Jinkela_wire_10286)
    );

    bfr new_Jinkela_buffer_3786 (
        .din(new_Jinkela_wire_4408),
        .dout(new_Jinkela_wire_4409)
    );

    bfr new_Jinkela_buffer_692 (
        .din(new_Jinkela_wire_744),
        .dout(new_Jinkela_wire_745)
    );

    bfr new_Jinkela_buffer_3748 (
        .din(new_Jinkela_wire_4368),
        .dout(new_Jinkela_wire_4369)
    );

    bfr new_Jinkela_buffer_8219 (
        .din(new_Jinkela_wire_10322),
        .dout(new_Jinkela_wire_10323)
    );

    bfr new_Jinkela_buffer_819 (
        .din(N316),
        .dout(new_Jinkela_wire_880)
    );

    bfr new_Jinkela_buffer_883 (
        .din(N293),
        .dout(new_Jinkela_wire_949)
    );

    bfr new_Jinkela_buffer_8185 (
        .din(new_Jinkela_wire_10286),
        .dout(new_Jinkela_wire_10287)
    );

    bfr new_Jinkela_buffer_3810 (
        .din(new_net_2570),
        .dout(new_Jinkela_wire_4444)
    );

    bfr new_Jinkela_buffer_693 (
        .din(new_Jinkela_wire_745),
        .dout(new_Jinkela_wire_746)
    );

    bfr new_Jinkela_buffer_3749 (
        .din(new_Jinkela_wire_4369),
        .dout(new_Jinkela_wire_4370)
    );

    bfr new_Jinkela_buffer_748 (
        .din(new_Jinkela_wire_808),
        .dout(new_Jinkela_wire_809)
    );

    bfr new_Jinkela_buffer_3808 (
        .din(new_Jinkela_wire_4441),
        .dout(new_Jinkela_wire_4442)
    );

    bfr new_Jinkela_buffer_8186 (
        .din(new_Jinkela_wire_10287),
        .dout(new_Jinkela_wire_10288)
    );

    bfr new_Jinkela_buffer_3787 (
        .din(new_Jinkela_wire_4409),
        .dout(new_Jinkela_wire_4410)
    );

    bfr new_Jinkela_buffer_694 (
        .din(new_Jinkela_wire_746),
        .dout(new_Jinkela_wire_747)
    );

    bfr new_Jinkela_buffer_3750 (
        .din(new_Jinkela_wire_4370),
        .dout(new_Jinkela_wire_4371)
    );

    bfr new_Jinkela_buffer_2877 (
        .din(new_Jinkela_wire_3300),
        .dout(new_Jinkela_wire_3301)
    );

    spl2 new_Jinkela_splitter_330 (
        .a(new_Jinkela_wire_5452),
        .b(new_Jinkela_wire_5453),
        .c(new_Jinkela_wire_5454)
    );

    bfr new_Jinkela_buffer_2842 (
        .din(new_Jinkela_wire_3261),
        .dout(new_Jinkela_wire_3262)
    );

    bfr new_Jinkela_buffer_4554 (
        .din(new_Jinkela_wire_5426),
        .dout(new_Jinkela_wire_5427)
    );

    bfr new_Jinkela_buffer_2940 (
        .din(new_Jinkela_wire_3365),
        .dout(new_Jinkela_wire_3366)
    );

    bfr new_Jinkela_buffer_4578 (
        .din(new_Jinkela_wire_5454),
        .dout(new_Jinkela_wire_5455)
    );

    bfr new_Jinkela_buffer_2843 (
        .din(new_Jinkela_wire_3262),
        .dout(new_Jinkela_wire_3263)
    );

    bfr new_Jinkela_buffer_4555 (
        .din(new_Jinkela_wire_5427),
        .dout(new_Jinkela_wire_5428)
    );

    bfr new_Jinkela_buffer_2878 (
        .din(new_Jinkela_wire_3301),
        .dout(new_Jinkela_wire_3302)
    );

    bfr new_Jinkela_buffer_4622 (
        .din(new_Jinkela_wire_5500),
        .dout(new_Jinkela_wire_5501)
    );

    bfr new_Jinkela_buffer_2844 (
        .din(new_Jinkela_wire_3263),
        .dout(new_Jinkela_wire_3264)
    );

    bfr new_Jinkela_buffer_4556 (
        .din(new_Jinkela_wire_5428),
        .dout(new_Jinkela_wire_5429)
    );

    bfr new_Jinkela_buffer_3011 (
        .din(N110),
        .dout(new_Jinkela_wire_3439)
    );

    bfr new_Jinkela_buffer_4582 (
        .din(new_Jinkela_wire_5460),
        .dout(new_Jinkela_wire_5461)
    );

    bfr new_Jinkela_buffer_2845 (
        .din(new_Jinkela_wire_3264),
        .dout(new_Jinkela_wire_3265)
    );

    bfr new_Jinkela_buffer_4557 (
        .din(new_Jinkela_wire_5429),
        .dout(new_Jinkela_wire_5430)
    );

    bfr new_Jinkela_buffer_2879 (
        .din(new_Jinkela_wire_3302),
        .dout(new_Jinkela_wire_3303)
    );

    bfr new_Jinkela_buffer_4579 (
        .din(new_Jinkela_wire_5455),
        .dout(new_Jinkela_wire_5456)
    );

    bfr new_Jinkela_buffer_2846 (
        .din(new_Jinkela_wire_3265),
        .dout(new_Jinkela_wire_3266)
    );

    bfr new_Jinkela_buffer_4558 (
        .din(new_Jinkela_wire_5430),
        .dout(new_Jinkela_wire_5431)
    );

    spl2 new_Jinkela_splitter_145 (
        .a(new_Jinkela_wire_3366),
        .b(new_Jinkela_wire_3367),
        .c(new_Jinkela_wire_3368)
    );

    spl2 new_Jinkela_splitter_332 (
        .a(new_net_8),
        .b(new_Jinkela_wire_5503),
        .c(new_Jinkela_wire_5504)
    );

    bfr new_Jinkela_buffer_2847 (
        .din(new_Jinkela_wire_3266),
        .dout(new_Jinkela_wire_3267)
    );

    bfr new_Jinkela_buffer_4559 (
        .din(new_Jinkela_wire_5431),
        .dout(new_Jinkela_wire_5432)
    );

    bfr new_Jinkela_buffer_2880 (
        .din(new_Jinkela_wire_3303),
        .dout(new_Jinkela_wire_3304)
    );

    bfr new_Jinkela_buffer_4583 (
        .din(new_Jinkela_wire_5461),
        .dout(new_Jinkela_wire_5462)
    );

    bfr new_Jinkela_buffer_4580 (
        .din(new_Jinkela_wire_5456),
        .dout(new_Jinkela_wire_5457)
    );

    bfr new_Jinkela_buffer_2848 (
        .din(new_Jinkela_wire_3267),
        .dout(new_Jinkela_wire_3268)
    );

    bfr new_Jinkela_buffer_4560 (
        .din(new_Jinkela_wire_5432),
        .dout(new_Jinkela_wire_5433)
    );

    bfr new_Jinkela_buffer_2941 (
        .din(new_Jinkela_wire_3368),
        .dout(new_Jinkela_wire_3369)
    );

    bfr new_Jinkela_buffer_2849 (
        .din(new_Jinkela_wire_3268),
        .dout(new_Jinkela_wire_3269)
    );

    bfr new_Jinkela_buffer_4561 (
        .din(new_Jinkela_wire_5433),
        .dout(new_Jinkela_wire_5434)
    );

    bfr new_Jinkela_buffer_2881 (
        .din(new_Jinkela_wire_3304),
        .dout(new_Jinkela_wire_3305)
    );

    bfr new_Jinkela_buffer_4624 (
        .din(new_net_2558),
        .dout(new_Jinkela_wire_5505)
    );

    bfr new_Jinkela_buffer_2850 (
        .din(new_Jinkela_wire_3269),
        .dout(new_Jinkela_wire_3270)
    );

    bfr new_Jinkela_buffer_4562 (
        .din(new_Jinkela_wire_5434),
        .dout(new_Jinkela_wire_5435)
    );

    bfr new_Jinkela_buffer_3005 (
        .din(new_Jinkela_wire_3432),
        .dout(new_Jinkela_wire_3433)
    );

    bfr new_Jinkela_buffer_4584 (
        .din(new_Jinkela_wire_5462),
        .dout(new_Jinkela_wire_5463)
    );

    bfr new_Jinkela_buffer_2882 (
        .din(new_Jinkela_wire_3305),
        .dout(new_Jinkela_wire_3306)
    );

    bfr new_Jinkela_buffer_4563 (
        .din(new_Jinkela_wire_5435),
        .dout(new_Jinkela_wire_5436)
    );

    bfr new_Jinkela_buffer_3008 (
        .din(new_Jinkela_wire_3435),
        .dout(new_Jinkela_wire_3436)
    );

    bfr new_Jinkela_buffer_4625 (
        .din(new_Jinkela_wire_5505),
        .dout(new_Jinkela_wire_5506)
    );

    bfr new_Jinkela_buffer_2883 (
        .din(new_Jinkela_wire_3306),
        .dout(new_Jinkela_wire_3307)
    );

    bfr new_Jinkela_buffer_4564 (
        .din(new_Jinkela_wire_5436),
        .dout(new_Jinkela_wire_5437)
    );

    bfr new_Jinkela_buffer_2942 (
        .din(new_Jinkela_wire_3369),
        .dout(new_Jinkela_wire_3370)
    );

    bfr new_Jinkela_buffer_4585 (
        .din(new_Jinkela_wire_5463),
        .dout(new_Jinkela_wire_5464)
    );

    bfr new_Jinkela_buffer_2884 (
        .din(new_Jinkela_wire_3307),
        .dout(new_Jinkela_wire_3308)
    );

    bfr new_Jinkela_buffer_4565 (
        .din(new_Jinkela_wire_5437),
        .dout(new_Jinkela_wire_5438)
    );

    bfr new_Jinkela_buffer_3006 (
        .din(new_Jinkela_wire_3433),
        .dout(new_Jinkela_wire_3434)
    );

    bfr new_Jinkela_buffer_4673 (
        .din(n_1198_),
        .dout(new_Jinkela_wire_5554)
    );

    bfr new_Jinkela_buffer_2885 (
        .din(new_Jinkela_wire_3308),
        .dout(new_Jinkela_wire_3309)
    );

    bfr new_Jinkela_buffer_4566 (
        .din(new_Jinkela_wire_5438),
        .dout(new_Jinkela_wire_5439)
    );

    bfr new_Jinkela_buffer_2943 (
        .din(new_Jinkela_wire_3370),
        .dout(new_Jinkela_wire_3371)
    );

    bfr new_Jinkela_buffer_4586 (
        .din(new_Jinkela_wire_5464),
        .dout(new_Jinkela_wire_5465)
    );

    bfr new_Jinkela_buffer_2886 (
        .din(new_Jinkela_wire_3309),
        .dout(new_Jinkela_wire_3310)
    );

    bfr new_Jinkela_buffer_4567 (
        .din(new_Jinkela_wire_5439),
        .dout(new_Jinkela_wire_5440)
    );

    bfr new_Jinkela_buffer_3015 (
        .din(N274),
        .dout(new_Jinkela_wire_3443)
    );

    bfr new_Jinkela_buffer_3080 (
        .din(N100),
        .dout(new_Jinkela_wire_3510)
    );

    bfr new_Jinkela_buffer_4674 (
        .din(n_0855_),
        .dout(new_Jinkela_wire_5555)
    );

    bfr new_Jinkela_buffer_2887 (
        .din(new_Jinkela_wire_3310),
        .dout(new_Jinkela_wire_3311)
    );

    bfr new_Jinkela_buffer_4568 (
        .din(new_Jinkela_wire_5440),
        .dout(new_Jinkela_wire_5441)
    );

    bfr new_Jinkela_buffer_2944 (
        .din(new_Jinkela_wire_3371),
        .dout(new_Jinkela_wire_3372)
    );

    bfr new_Jinkela_buffer_4587 (
        .din(new_Jinkela_wire_5465),
        .dout(new_Jinkela_wire_5466)
    );

    bfr new_Jinkela_buffer_2888 (
        .din(new_Jinkela_wire_3311),
        .dout(new_Jinkela_wire_3312)
    );

    bfr new_Jinkela_buffer_4569 (
        .din(new_Jinkela_wire_5441),
        .dout(new_Jinkela_wire_5442)
    );

    bfr new_Jinkela_buffer_3009 (
        .din(new_Jinkela_wire_3436),
        .dout(new_Jinkela_wire_3437)
    );

    bfr new_Jinkela_buffer_4626 (
        .din(new_Jinkela_wire_5506),
        .dout(new_Jinkela_wire_5507)
    );

    bfr new_Jinkela_buffer_2889 (
        .din(new_Jinkela_wire_3312),
        .dout(new_Jinkela_wire_3313)
    );

    bfr new_Jinkela_buffer_4570 (
        .din(new_Jinkela_wire_5442),
        .dout(new_Jinkela_wire_5443)
    );

    bfr new_Jinkela_buffer_2945 (
        .din(new_Jinkela_wire_3372),
        .dout(new_Jinkela_wire_3373)
    );

    bfr new_Jinkela_buffer_4588 (
        .din(new_Jinkela_wire_5466),
        .dout(new_Jinkela_wire_5467)
    );

    bfr new_Jinkela_buffer_2890 (
        .din(new_Jinkela_wire_3313),
        .dout(new_Jinkela_wire_3314)
    );

    bfr new_Jinkela_buffer_4571 (
        .din(new_Jinkela_wire_5443),
        .dout(new_Jinkela_wire_5444)
    );

    bfr new_Jinkela_buffer_3012 (
        .din(new_Jinkela_wire_3439),
        .dout(new_Jinkela_wire_3440)
    );

    bfr new_Jinkela_buffer_2891 (
        .din(new_Jinkela_wire_3314),
        .dout(new_Jinkela_wire_3315)
    );

    bfr new_Jinkela_buffer_413 (
        .din(new_Jinkela_wire_449),
        .dout(new_Jinkela_wire_450)
    );

    bfr new_Jinkela_buffer_4675 (
        .din(n_0966_),
        .dout(new_Jinkela_wire_5556)
    );

    bfr new_Jinkela_buffer_4572 (
        .din(new_Jinkela_wire_5444),
        .dout(new_Jinkela_wire_5445)
    );

    bfr new_Jinkela_buffer_2946 (
        .din(new_Jinkela_wire_3373),
        .dout(new_Jinkela_wire_3374)
    );

    bfr new_Jinkela_buffer_4589 (
        .din(new_Jinkela_wire_5467),
        .dout(new_Jinkela_wire_5468)
    );

    bfr new_Jinkela_buffer_2892 (
        .din(new_Jinkela_wire_3315),
        .dout(new_Jinkela_wire_3316)
    );

    bfr new_Jinkela_buffer_4573 (
        .din(new_Jinkela_wire_5445),
        .dout(new_Jinkela_wire_5446)
    );

    bfr new_Jinkela_buffer_3010 (
        .din(new_Jinkela_wire_3437),
        .dout(new_Jinkela_wire_3438)
    );

    bfr new_Jinkela_buffer_4676 (
        .din(n_0517_),
        .dout(new_Jinkela_wire_5559)
    );

    bfr new_Jinkela_buffer_4627 (
        .din(new_Jinkela_wire_5507),
        .dout(new_Jinkela_wire_5508)
    );

    bfr new_Jinkela_buffer_2893 (
        .din(new_Jinkela_wire_3316),
        .dout(new_Jinkela_wire_3317)
    );

    bfr new_Jinkela_buffer_4574 (
        .din(new_Jinkela_wire_5446),
        .dout(new_Jinkela_wire_5447)
    );

    bfr new_Jinkela_buffer_5425 (
        .din(new_Jinkela_wire_6504),
        .dout(new_Jinkela_wire_6505)
    );

    bfr new_Jinkela_buffer_5398 (
        .din(new_Jinkela_wire_6477),
        .dout(new_Jinkela_wire_6478)
    );

    bfr new_Jinkela_buffer_7712 (
        .din(new_Jinkela_wire_9703),
        .dout(new_Jinkela_wire_9704)
    );

    spl2 new_Jinkela_splitter_800 (
        .a(n_0680_),
        .b(new_Jinkela_wire_9732),
        .c(new_Jinkela_wire_9733)
    );

    bfr new_Jinkela_buffer_7658 (
        .din(new_Jinkela_wire_9632),
        .dout(new_Jinkela_wire_9633)
    );

    bfr new_Jinkela_buffer_5399 (
        .din(new_Jinkela_wire_6478),
        .dout(new_Jinkela_wire_6479)
    );

    bfr new_Jinkela_buffer_7679 (
        .din(new_Jinkela_wire_9665),
        .dout(new_Jinkela_wire_9666)
    );

    bfr new_Jinkela_buffer_5444 (
        .din(new_Jinkela_wire_6541),
        .dout(new_Jinkela_wire_6542)
    );

    bfr new_Jinkela_buffer_7659 (
        .din(new_Jinkela_wire_9633),
        .dout(new_Jinkela_wire_9634)
    );

    bfr new_Jinkela_buffer_5426 (
        .din(new_Jinkela_wire_6505),
        .dout(new_Jinkela_wire_6506)
    );

    bfr new_Jinkela_buffer_5400 (
        .din(new_Jinkela_wire_6479),
        .dout(new_Jinkela_wire_6480)
    );

    spl2 new_Jinkela_splitter_806 (
        .a(n_1139_),
        .b(new_Jinkela_wire_9755),
        .c(new_Jinkela_wire_9756)
    );

    bfr new_Jinkela_buffer_7670 (
        .din(new_Jinkela_wire_9654),
        .dout(new_Jinkela_wire_9655)
    );

    bfr new_Jinkela_buffer_7660 (
        .din(new_Jinkela_wire_9634),
        .dout(new_Jinkela_wire_9635)
    );

    bfr new_Jinkela_buffer_5451 (
        .din(new_net_2572),
        .dout(new_Jinkela_wire_6549)
    );

    bfr new_Jinkela_buffer_5401 (
        .din(new_Jinkela_wire_6480),
        .dout(new_Jinkela_wire_6481)
    );

    spl4L new_Jinkela_splitter_799 (
        .a(new_Jinkela_wire_9705),
        .d(new_Jinkela_wire_9706),
        .b(new_Jinkela_wire_9707),
        .e(new_Jinkela_wire_9708),
        .c(new_Jinkela_wire_9709)
    );

    bfr new_Jinkela_buffer_7661 (
        .din(new_Jinkela_wire_9635),
        .dout(new_Jinkela_wire_9636)
    );

    bfr new_Jinkela_buffer_5427 (
        .din(new_Jinkela_wire_6506),
        .dout(new_Jinkela_wire_6507)
    );

    bfr new_Jinkela_buffer_5402 (
        .din(new_Jinkela_wire_6481),
        .dout(new_Jinkela_wire_6482)
    );

    bfr new_Jinkela_buffer_7671 (
        .din(new_Jinkela_wire_9655),
        .dout(new_Jinkela_wire_9656)
    );

    bfr new_Jinkela_buffer_7662 (
        .din(new_Jinkela_wire_9636),
        .dout(new_Jinkela_wire_9637)
    );

    spl4L new_Jinkela_splitter_426 (
        .a(n_0145_),
        .d(new_Jinkela_wire_6555),
        .b(new_Jinkela_wire_6556),
        .e(new_Jinkela_wire_6557),
        .c(new_Jinkela_wire_6558)
    );

    bfr new_Jinkela_buffer_5403 (
        .din(new_Jinkela_wire_6482),
        .dout(new_Jinkela_wire_6483)
    );

    bfr new_Jinkela_buffer_5465 (
        .din(n_0174_),
        .dout(new_Jinkela_wire_6567)
    );

    bfr new_Jinkela_buffer_7663 (
        .din(new_Jinkela_wire_9637),
        .dout(new_Jinkela_wire_9638)
    );

    bfr new_Jinkela_buffer_5428 (
        .din(new_Jinkela_wire_6507),
        .dout(new_Jinkela_wire_6508)
    );

    bfr new_Jinkela_buffer_5404 (
        .din(new_Jinkela_wire_6483),
        .dout(new_Jinkela_wire_6484)
    );

    spl2 new_Jinkela_splitter_795 (
        .a(new_Jinkela_wire_9656),
        .b(new_Jinkela_wire_9657),
        .c(new_Jinkela_wire_9658)
    );

    spl2 new_Jinkela_splitter_791 (
        .a(new_Jinkela_wire_9638),
        .b(new_Jinkela_wire_9639),
        .c(new_Jinkela_wire_9640)
    );

    bfr new_Jinkela_buffer_5445 (
        .din(new_Jinkela_wire_6542),
        .dout(new_Jinkela_wire_6543)
    );

    bfr new_Jinkela_buffer_7714 (
        .din(new_Jinkela_wire_9710),
        .dout(new_Jinkela_wire_9711)
    );

    bfr new_Jinkela_buffer_5429 (
        .din(new_Jinkela_wire_6508),
        .dout(new_Jinkela_wire_6509)
    );

    bfr new_Jinkela_buffer_7672 (
        .din(new_Jinkela_wire_9658),
        .dout(new_Jinkela_wire_9659)
    );

    bfr new_Jinkela_buffer_5452 (
        .din(new_Jinkela_wire_6549),
        .dout(new_Jinkela_wire_6550)
    );

    bfr new_Jinkela_buffer_7715 (
        .din(new_Jinkela_wire_9711),
        .dout(new_Jinkela_wire_9712)
    );

    bfr new_Jinkela_buffer_5430 (
        .din(new_Jinkela_wire_6509),
        .dout(new_Jinkela_wire_6510)
    );

    bfr new_Jinkela_buffer_360 (
        .din(new_Jinkela_wire_391),
        .dout(new_Jinkela_wire_392)
    );

    bfr new_Jinkela_buffer_7673 (
        .din(new_Jinkela_wire_9659),
        .dout(new_Jinkela_wire_9660)
    );

    bfr new_Jinkela_buffer_5446 (
        .din(new_Jinkela_wire_6543),
        .dout(new_Jinkela_wire_6544)
    );

    bfr new_Jinkela_buffer_5431 (
        .din(new_Jinkela_wire_6510),
        .dout(new_Jinkela_wire_6511)
    );

    bfr new_Jinkela_buffer_7674 (
        .din(new_Jinkela_wire_9660),
        .dout(new_Jinkela_wire_9661)
    );

    bfr new_Jinkela_buffer_5457 (
        .din(new_Jinkela_wire_6558),
        .dout(new_Jinkela_wire_6559)
    );

    bfr new_Jinkela_buffer_7716 (
        .din(new_Jinkela_wire_9712),
        .dout(new_Jinkela_wire_9713)
    );

    bfr new_Jinkela_buffer_5432 (
        .din(new_Jinkela_wire_6511),
        .dout(new_Jinkela_wire_6512)
    );

    bfr new_Jinkela_buffer_7675 (
        .din(new_Jinkela_wire_9661),
        .dout(new_Jinkela_wire_9662)
    );

    bfr new_Jinkela_buffer_5447 (
        .din(new_Jinkela_wire_6544),
        .dout(new_Jinkela_wire_6545)
    );

    bfr new_Jinkela_buffer_7735 (
        .din(new_Jinkela_wire_9733),
        .dout(new_Jinkela_wire_9734)
    );

    bfr new_Jinkela_buffer_5453 (
        .din(new_Jinkela_wire_6550),
        .dout(new_Jinkela_wire_6551)
    );

    bfr new_Jinkela_buffer_7676 (
        .din(new_Jinkela_wire_9662),
        .dout(new_Jinkela_wire_9663)
    );

    bfr new_Jinkela_buffer_5448 (
        .din(new_Jinkela_wire_6545),
        .dout(new_Jinkela_wire_6546)
    );

    bfr new_Jinkela_buffer_7717 (
        .din(new_Jinkela_wire_9713),
        .dout(new_Jinkela_wire_9714)
    );

    bfr new_Jinkela_buffer_5466 (
        .din(new_Jinkela_wire_6567),
        .dout(new_Jinkela_wire_6568)
    );

    bfr new_Jinkela_buffer_7677 (
        .din(new_Jinkela_wire_9663),
        .dout(new_Jinkela_wire_9664)
    );

    bfr new_Jinkela_buffer_5449 (
        .din(new_Jinkela_wire_6546),
        .dout(new_Jinkela_wire_6547)
    );

    bfr new_Jinkela_buffer_7742 (
        .din(n_0435_),
        .dout(new_Jinkela_wire_9749)
    );

    spl3L new_Jinkela_splitter_804 (
        .a(n_0927_),
        .d(new_Jinkela_wire_9750),
        .b(new_Jinkela_wire_9751),
        .c(new_Jinkela_wire_9752)
    );

    bfr new_Jinkela_buffer_5454 (
        .din(new_Jinkela_wire_6551),
        .dout(new_Jinkela_wire_6552)
    );

    bfr new_Jinkela_buffer_361 (
        .din(new_Jinkela_wire_392),
        .dout(new_Jinkela_wire_393)
    );

    bfr new_Jinkela_buffer_7678 (
        .din(new_Jinkela_wire_9664),
        .dout(new_Jinkela_wire_9665)
    );

    bfr new_Jinkela_buffer_5450 (
        .din(new_Jinkela_wire_6547),
        .dout(new_Jinkela_wire_6548)
    );

    bfr new_Jinkela_buffer_7718 (
        .din(new_Jinkela_wire_9714),
        .dout(new_Jinkela_wire_9715)
    );

    spl3L new_Jinkela_splitter_427 (
        .a(n_0039_),
        .d(new_Jinkela_wire_6604),
        .b(new_Jinkela_wire_6605),
        .c(new_Jinkela_wire_6606)
    );

    bfr new_Jinkela_buffer_7680 (
        .din(new_Jinkela_wire_9666),
        .dout(new_Jinkela_wire_9667)
    );

    bfr new_Jinkela_buffer_5455 (
        .din(new_Jinkela_wire_6552),
        .dout(new_Jinkela_wire_6553)
    );

    bfr new_Jinkela_buffer_7736 (
        .din(new_Jinkela_wire_9734),
        .dout(new_Jinkela_wire_9735)
    );

    bfr new_Jinkela_buffer_5535 (
        .din(n_0431_),
        .dout(new_Jinkela_wire_6640)
    );

    bfr new_Jinkela_buffer_5458 (
        .din(new_Jinkela_wire_6559),
        .dout(new_Jinkela_wire_6560)
    );

    spl2 new_Jinkela_splitter_807 (
        .a(n_0773_),
        .b(new_Jinkela_wire_9757),
        .c(new_Jinkela_wire_9758)
    );

    bfr new_Jinkela_buffer_5456 (
        .din(new_Jinkela_wire_6553),
        .dout(new_Jinkela_wire_6554)
    );

    bfr new_Jinkela_buffer_7719 (
        .din(new_Jinkela_wire_9715),
        .dout(new_Jinkela_wire_9716)
    );

    bfr new_Jinkela_buffer_7681 (
        .din(new_Jinkela_wire_9667),
        .dout(new_Jinkela_wire_9668)
    );

    bfr new_Jinkela_buffer_5459 (
        .din(new_Jinkela_wire_6560),
        .dout(new_Jinkela_wire_6561)
    );

    spl4L new_Jinkela_splitter_803 (
        .a(n_0673_),
        .d(new_Jinkela_wire_9745),
        .b(new_Jinkela_wire_9746),
        .e(new_Jinkela_wire_9747),
        .c(new_Jinkela_wire_9748)
    );

    bfr new_Jinkela_buffer_7682 (
        .din(new_Jinkela_wire_9668),
        .dout(new_Jinkela_wire_9669)
    );

    bfr new_Jinkela_buffer_5467 (
        .din(new_Jinkela_wire_6568),
        .dout(new_Jinkela_wire_6569)
    );

    bfr new_Jinkela_buffer_5460 (
        .din(new_Jinkela_wire_6561),
        .dout(new_Jinkela_wire_6562)
    );

    bfr new_Jinkela_buffer_7720 (
        .din(new_Jinkela_wire_9716),
        .dout(new_Jinkela_wire_9717)
    );

    bfr new_Jinkela_buffer_362 (
        .din(new_Jinkela_wire_393),
        .dout(new_Jinkela_wire_394)
    );

    bfr new_Jinkela_buffer_7683 (
        .din(new_Jinkela_wire_9669),
        .dout(new_Jinkela_wire_9670)
    );

    bfr new_Jinkela_buffer_5502 (
        .din(new_Jinkela_wire_6606),
        .dout(new_Jinkela_wire_6607)
    );

    bfr new_Jinkela_buffer_5461 (
        .din(new_Jinkela_wire_6562),
        .dout(new_Jinkela_wire_6563)
    );

    bfr new_Jinkela_buffer_7737 (
        .din(new_Jinkela_wire_9735),
        .dout(new_Jinkela_wire_9736)
    );

    spl2 new_Jinkela_splitter_429 (
        .a(n_1185_),
        .b(new_Jinkela_wire_6672),
        .c(new_Jinkela_wire_6673)
    );

    bfr new_Jinkela_buffer_7684 (
        .din(new_Jinkela_wire_9670),
        .dout(new_Jinkela_wire_9671)
    );

    bfr new_Jinkela_buffer_5468 (
        .din(new_Jinkela_wire_6569),
        .dout(new_Jinkela_wire_6570)
    );

    bfr new_Jinkela_buffer_5462 (
        .din(new_Jinkela_wire_6563),
        .dout(new_Jinkela_wire_6564)
    );

    bfr new_Jinkela_buffer_7721 (
        .din(new_Jinkela_wire_9717),
        .dout(new_Jinkela_wire_9718)
    );

    bfr new_Jinkela_buffer_7685 (
        .din(new_Jinkela_wire_9671),
        .dout(new_Jinkela_wire_9672)
    );

    bfr new_Jinkela_buffer_1158 (
        .din(new_Jinkela_wire_1469),
        .dout(new_Jinkela_wire_1470)
    );

    or_bb n_2241_ (
        .a(n_0126_),
        .b(n_0125_),
        .c(new_net_2497)
    );

    bfr new_Jinkela_buffer_1190 (
        .din(new_Jinkela_wire_1506),
        .dout(new_Jinkela_wire_1507)
    );

    and_bi n_2242_ (
        .a(new_Jinkela_wire_5144),
        .b(new_Jinkela_wire_7066),
        .c(n_0127_)
    );

    bfr new_Jinkela_buffer_478 (
        .din(new_Jinkela_wire_516),
        .dout(new_Jinkela_wire_517)
    );

    bfr new_Jinkela_buffer_1159 (
        .din(new_Jinkela_wire_1470),
        .dout(new_Jinkela_wire_1471)
    );

    or_bi n_2243_ (
        .a(n_0127_),
        .b(new_Jinkela_wire_6058),
        .c(n_0128_)
    );

    bfr new_Jinkela_buffer_1238 (
        .din(new_Jinkela_wire_1558),
        .dout(new_Jinkela_wire_1559)
    );

    and_bi n_2244_ (
        .a(new_Jinkela_wire_5279),
        .b(new_Jinkela_wire_9088),
        .c(n_0129_)
    );

    bfr new_Jinkela_buffer_1191 (
        .din(new_Jinkela_wire_1507),
        .dout(new_Jinkela_wire_1508)
    );

    and_bi n_2245_ (
        .a(new_Jinkela_wire_9087),
        .b(new_Jinkela_wire_5278),
        .c(n_0130_)
    );

    bfr new_Jinkela_buffer_1360 (
        .din(new_Jinkela_wire_1685),
        .dout(new_Jinkela_wire_1686)
    );

    or_bb n_2246_ (
        .a(n_0130_),
        .b(n_0129_),
        .c(new_net_2537)
    );

    bfr new_Jinkela_buffer_1192 (
        .din(new_Jinkela_wire_1508),
        .dout(new_Jinkela_wire_1509)
    );

    and_ii n_2247_ (
        .a(new_Jinkela_wire_4012),
        .b(new_Jinkela_wire_6484),
        .c(n_0131_)
    );

    bfr new_Jinkela_buffer_1239 (
        .din(new_Jinkela_wire_1559),
        .dout(new_Jinkela_wire_1560)
    );

    and_bi n_2248_ (
        .a(new_Jinkela_wire_5592),
        .b(new_Jinkela_wire_5803),
        .c(n_0132_)
    );

    bfr new_Jinkela_buffer_1193 (
        .din(new_Jinkela_wire_1509),
        .dout(new_Jinkela_wire_1510)
    );

    and_bi n_2249_ (
        .a(new_Jinkela_wire_5804),
        .b(new_Jinkela_wire_5591),
        .c(n_0133_)
    );

    bfr new_Jinkela_buffer_1298 (
        .din(new_Jinkela_wire_1620),
        .dout(new_Jinkela_wire_1621)
    );

    and_ii n_2250_ (
        .a(n_0133_),
        .b(n_0132_),
        .c(new_net_2572)
    );

    bfr new_Jinkela_buffer_1194 (
        .din(new_Jinkela_wire_1510),
        .dout(new_Jinkela_wire_1511)
    );

    or_bb n_2251_ (
        .a(new_Jinkela_wire_3610),
        .b(new_Jinkela_wire_8199),
        .c(n_0134_)
    );

    bfr new_Jinkela_buffer_1240 (
        .din(new_Jinkela_wire_1560),
        .dout(new_Jinkela_wire_1561)
    );

    or_bb n_2252_ (
        .a(new_Jinkela_wire_10229),
        .b(new_Jinkela_wire_10154),
        .c(n_0135_)
    );

    bfr new_Jinkela_buffer_416 (
        .din(new_Jinkela_wire_452),
        .dout(new_Jinkela_wire_453)
    );

    bfr new_Jinkela_buffer_1195 (
        .din(new_Jinkela_wire_1511),
        .dout(new_Jinkela_wire_1512)
    );

    or_bb n_2253_ (
        .a(n_0135_),
        .b(n_0134_),
        .c(n_0136_)
    );

    bfr new_Jinkela_buffer_1369 (
        .din(N79),
        .dout(new_Jinkela_wire_1695)
    );

    or_bb n_2254_ (
        .a(new_Jinkela_wire_4427),
        .b(new_Jinkela_wire_9984),
        .c(n_0137_)
    );

    bfr new_Jinkela_buffer_1196 (
        .din(new_Jinkela_wire_1512),
        .dout(new_Jinkela_wire_1513)
    );

    or_bb n_2255_ (
        .a(new_Jinkela_wire_8578),
        .b(new_Jinkela_wire_10295),
        .c(n_0138_)
    );

    bfr new_Jinkela_buffer_1241 (
        .din(new_Jinkela_wire_1561),
        .dout(new_Jinkela_wire_1562)
    );

    or_bb n_2256_ (
        .a(n_0138_),
        .b(n_0137_),
        .c(new_net_2560)
    );

    bfr new_Jinkela_buffer_1197 (
        .din(new_Jinkela_wire_1513),
        .dout(new_Jinkela_wire_1514)
    );

    and_bi n_2257_ (
        .a(new_Jinkela_wire_9931),
        .b(new_Jinkela_wire_9397),
        .c(n_0139_)
    );

    spl3L new_Jinkela_splitter_101 (
        .a(new_Jinkela_wire_1621),
        .d(new_Jinkela_wire_1622),
        .b(new_Jinkela_wire_1623),
        .c(new_Jinkela_wire_1624)
    );

    and_bi n_2258_ (
        .a(new_Jinkela_wire_6129),
        .b(new_Jinkela_wire_9433),
        .c(n_0140_)
    );

    bfr new_Jinkela_buffer_1198 (
        .din(new_Jinkela_wire_1514),
        .dout(new_Jinkela_wire_1515)
    );

    and_bi n_2259_ (
        .a(new_Jinkela_wire_9432),
        .b(new_Jinkela_wire_6128),
        .c(n_0141_)
    );

    bfr new_Jinkela_buffer_1242 (
        .din(new_Jinkela_wire_1562),
        .dout(new_Jinkela_wire_1563)
    );

    and_ii n_2260_ (
        .a(new_Jinkela_wire_9581),
        .b(new_Jinkela_wire_10032),
        .c(new_net_2525)
    );

    bfr new_Jinkela_buffer_1199 (
        .din(new_Jinkela_wire_1515),
        .dout(new_Jinkela_wire_1516)
    );

    or_bb n_2261_ (
        .a(new_Jinkela_wire_9428),
        .b(new_Jinkela_wire_3693),
        .c(n_0142_)
    );

    bfr new_Jinkela_buffer_1363 (
        .din(new_Jinkela_wire_1688),
        .dout(new_Jinkela_wire_1689)
    );

    and_ii n_2262_ (
        .a(new_Jinkela_wire_5161),
        .b(new_Jinkela_wire_7321),
        .c(n_0143_)
    );

    bfr new_Jinkela_buffer_1200 (
        .din(new_Jinkela_wire_1516),
        .dout(new_Jinkela_wire_1517)
    );

    and_bb n_2263_ (
        .a(new_Jinkela_wire_5162),
        .b(new_Jinkela_wire_7320),
        .c(n_0144_)
    );

    bfr new_Jinkela_buffer_1243 (
        .din(new_Jinkela_wire_1563),
        .dout(new_Jinkela_wire_1564)
    );

    and_ii n_2264_ (
        .a(n_0144_),
        .b(n_0143_),
        .c(n_0145_)
    );

    bfr new_Jinkela_buffer_1201 (
        .din(new_Jinkela_wire_1517),
        .dout(new_Jinkela_wire_1518)
    );

    and_bi n_2265_ (
        .a(n_0142_),
        .b(new_Jinkela_wire_6566),
        .c(n_0146_)
    );

    bfr new_Jinkela_buffer_1299 (
        .din(new_Jinkela_wire_1624),
        .dout(new_Jinkela_wire_1625)
    );

    and_bi n_2266_ (
        .a(new_Jinkela_wire_8512),
        .b(n_0146_),
        .c(new_net_2543)
    );

    bfr new_Jinkela_buffer_1202 (
        .din(new_Jinkela_wire_1518),
        .dout(new_Jinkela_wire_1519)
    );

    and_bb n_2267_ (
        .a(new_Jinkela_wire_5984),
        .b(new_Jinkela_wire_7838),
        .c(n_0147_)
    );

    bfr new_Jinkela_buffer_1244 (
        .din(new_Jinkela_wire_1564),
        .dout(new_Jinkela_wire_1565)
    );

    and_bi n_2268_ (
        .a(new_Jinkela_wire_4501),
        .b(new_Jinkela_wire_9427),
        .c(n_0148_)
    );

    bfr new_Jinkela_buffer_1203 (
        .din(new_Jinkela_wire_1519),
        .dout(new_Jinkela_wire_1520)
    );

    and_bi n_2269_ (
        .a(new_Jinkela_wire_3609),
        .b(n_0148_),
        .c(n_0149_)
    );

    bfr new_Jinkela_buffer_1366 (
        .din(new_Jinkela_wire_1691),
        .dout(new_Jinkela_wire_1692)
    );

    or_ii n_2270_ (
        .a(new_Jinkela_wire_5568),
        .b(new_Jinkela_wire_8648),
        .c(n_0150_)
    );

    bfr new_Jinkela_buffer_1204 (
        .din(new_Jinkela_wire_1520),
        .dout(new_Jinkela_wire_1521)
    );

    or_bb n_2271_ (
        .a(new_Jinkela_wire_5567),
        .b(new_Jinkela_wire_8649),
        .c(n_0151_)
    );

    bfr new_Jinkela_buffer_1245 (
        .din(new_Jinkela_wire_1565),
        .dout(new_Jinkela_wire_1566)
    );

    or_ii n_2272_ (
        .a(n_0151_),
        .b(n_0150_),
        .c(new_net_2511)
    );

    bfr new_Jinkela_buffer_1205 (
        .din(new_Jinkela_wire_1521),
        .dout(new_Jinkela_wire_1522)
    );

    and_ii n_2273_ (
        .a(new_Jinkela_wire_8758),
        .b(new_Jinkela_wire_4080),
        .c(n_0152_)
    );

    bfr new_Jinkela_buffer_1300 (
        .din(new_Jinkela_wire_1625),
        .dout(new_Jinkela_wire_1626)
    );

    inv n_2274_ (
        .din(new_Jinkela_wire_8944),
        .dout(n_0153_)
    );

    bfr new_Jinkela_buffer_1206 (
        .din(new_Jinkela_wire_1522),
        .dout(new_Jinkela_wire_1523)
    );

    and_bi n_2275_ (
        .a(new_Jinkela_wire_10030),
        .b(new_Jinkela_wire_6922),
        .c(n_0154_)
    );

    bfr new_Jinkela_buffer_1246 (
        .din(new_Jinkela_wire_1566),
        .dout(new_Jinkela_wire_1567)
    );

    or_bi n_2276_ (
        .a(n_0154_),
        .b(new_Jinkela_wire_5391),
        .c(n_0155_)
    );

    bfr new_Jinkela_buffer_1207 (
        .din(new_Jinkela_wire_1523),
        .dout(new_Jinkela_wire_1524)
    );

    and_bi n_2277_ (
        .a(new_Jinkela_wire_7544),
        .b(new_Jinkela_wire_6007),
        .c(n_0156_)
    );

    bfr new_Jinkela_buffer_1364 (
        .din(new_Jinkela_wire_1689),
        .dout(new_Jinkela_wire_1690)
    );

    and_bi n_2278_ (
        .a(new_Jinkela_wire_6006),
        .b(new_Jinkela_wire_7543),
        .c(n_0157_)
    );

    bfr new_Jinkela_buffer_1208 (
        .din(new_Jinkela_wire_1524),
        .dout(new_Jinkela_wire_1525)
    );

    or_bb n_2279_ (
        .a(n_0157_),
        .b(n_0156_),
        .c(new_net_2523)
    );

    bfr new_Jinkela_buffer_1247 (
        .din(new_Jinkela_wire_1567),
        .dout(new_Jinkela_wire_1568)
    );

    and_bi n_2280_ (
        .a(new_Jinkela_wire_9954),
        .b(new_Jinkela_wire_10031),
        .c(n_0158_)
    );

    bfr new_Jinkela_buffer_1209 (
        .din(new_Jinkela_wire_1525),
        .dout(new_Jinkela_wire_1526)
    );

    and_bi n_2281_ (
        .a(new_Jinkela_wire_7996),
        .b(new_Jinkela_wire_6926),
        .c(n_0159_)
    );

    bfr new_Jinkela_buffer_1301 (
        .din(new_Jinkela_wire_1626),
        .dout(new_Jinkela_wire_1627)
    );

    and_bi n_2282_ (
        .a(new_Jinkela_wire_6925),
        .b(new_Jinkela_wire_7995),
        .c(n_0160_)
    );

    bfr new_Jinkela_buffer_7627 (
        .din(new_Jinkela_wire_9568),
        .dout(new_Jinkela_wire_9569)
    );

    bfr new_Jinkela_buffer_8220 (
        .din(new_Jinkela_wire_10323),
        .dout(new_Jinkela_wire_10324)
    );

    and_ii n_1527_ (
        .a(n_0794_),
        .b(n_0793_),
        .c(n_0795_)
    );

    bfr new_Jinkela_buffer_7637 (
        .din(new_Jinkela_wire_9606),
        .dout(new_Jinkela_wire_9607)
    );

    bfr new_Jinkela_buffer_8187 (
        .din(new_Jinkela_wire_10288),
        .dout(new_Jinkela_wire_10289)
    );

    or_bi n_1528_ (
        .a(new_Jinkela_wire_9844),
        .b(new_Jinkela_wire_5589),
        .c(n_0796_)
    );

    bfr new_Jinkela_buffer_367 (
        .din(new_Jinkela_wire_398),
        .dout(new_Jinkela_wire_399)
    );

    bfr new_Jinkela_buffer_7631 (
        .din(new_Jinkela_wire_9589),
        .dout(new_Jinkela_wire_9590)
    );

    spl2 new_Jinkela_splitter_852 (
        .a(n_1316_),
        .b(new_Jinkela_wire_10390),
        .c(new_Jinkela_wire_10391)
    );

    and_bi n_1529_ (
        .a(new_Jinkela_wire_9843),
        .b(new_Jinkela_wire_5588),
        .c(n_0797_)
    );

    bfr new_Jinkela_buffer_8253 (
        .din(new_Jinkela_wire_10356),
        .dout(new_Jinkela_wire_10357)
    );

    bfr new_Jinkela_buffer_8188 (
        .din(new_Jinkela_wire_10289),
        .dout(new_Jinkela_wire_10290)
    );

    and_bi n_1530_ (
        .a(n_0796_),
        .b(n_0797_),
        .c(n_0798_)
    );

    spl2 new_Jinkela_splitter_784 (
        .a(new_Jinkela_wire_9590),
        .b(new_Jinkela_wire_9591),
        .c(new_Jinkela_wire_9592)
    );

    bfr new_Jinkela_buffer_8221 (
        .din(new_Jinkela_wire_10324),
        .dout(new_Jinkela_wire_10325)
    );

    and_ii n_1531_ (
        .a(new_Jinkela_wire_3932),
        .b(new_Jinkela_wire_4963),
        .c(n_0799_)
    );

    bfr new_Jinkela_buffer_7632 (
        .din(new_Jinkela_wire_9592),
        .dout(new_Jinkela_wire_9593)
    );

    bfr new_Jinkela_buffer_8189 (
        .din(new_Jinkela_wire_10290),
        .dout(new_Jinkela_wire_10291)
    );

    or_bb n_1532_ (
        .a(n_0799_),
        .b(new_Jinkela_wire_7933),
        .c(n_0800_)
    );

    bfr new_Jinkela_buffer_7636 (
        .din(n_0581_),
        .dout(new_Jinkela_wire_9606)
    );

    or_bb n_1533_ (
        .a(n_0800_),
        .b(new_Jinkela_wire_6428),
        .c(n_0801_)
    );

    bfr new_Jinkela_buffer_7640 (
        .din(n_0337_),
        .dout(new_Jinkela_wire_9610)
    );

    bfr new_Jinkela_buffer_8190 (
        .din(new_Jinkela_wire_10291),
        .dout(new_Jinkela_wire_10292)
    );

    and_bb n_1534_ (
        .a(new_Jinkela_wire_1089),
        .b(new_Jinkela_wire_1316),
        .c(n_0802_)
    );

    spl3L new_Jinkela_splitter_789 (
        .a(n_0775_),
        .d(new_Jinkela_wire_9617),
        .b(new_Jinkela_wire_9618),
        .c(new_Jinkela_wire_9619)
    );

    bfr new_Jinkela_buffer_7633 (
        .din(new_Jinkela_wire_9593),
        .dout(new_Jinkela_wire_9594)
    );

    bfr new_Jinkela_buffer_8222 (
        .din(new_Jinkela_wire_10325),
        .dout(new_Jinkela_wire_10326)
    );

    and_bi n_1535_ (
        .a(new_Jinkela_wire_879),
        .b(new_Jinkela_wire_1389),
        .c(n_0803_)
    );

    bfr new_Jinkela_buffer_7647 (
        .din(n_0810_),
        .dout(new_Jinkela_wire_9620)
    );

    bfr new_Jinkela_buffer_8191 (
        .din(new_Jinkela_wire_10292),
        .dout(new_Jinkela_wire_10293)
    );

    and_ii n_1536_ (
        .a(new_Jinkela_wire_7275),
        .b(new_Jinkela_wire_10101),
        .c(n_0804_)
    );

    bfr new_Jinkela_buffer_7638 (
        .din(new_Jinkela_wire_9607),
        .dout(new_Jinkela_wire_9608)
    );

    bfr new_Jinkela_buffer_7634 (
        .din(new_Jinkela_wire_9594),
        .dout(new_Jinkela_wire_9595)
    );

    bfr new_Jinkela_buffer_8261 (
        .din(new_Jinkela_wire_10373),
        .dout(new_Jinkela_wire_10374)
    );

    and_bb n_1537_ (
        .a(new_Jinkela_wire_438),
        .b(new_Jinkela_wire_1366),
        .c(n_0805_)
    );

    bfr new_Jinkela_buffer_8254 (
        .din(new_Jinkela_wire_10357),
        .dout(new_Jinkela_wire_10358)
    );

    bfr new_Jinkela_buffer_8223 (
        .din(new_Jinkela_wire_10326),
        .dout(new_Jinkela_wire_10327)
    );

    and_bi n_1538_ (
        .a(new_Jinkela_wire_8362),
        .b(new_Jinkela_wire_4630),
        .c(n_0806_)
    );

    bfr new_Jinkela_buffer_7641 (
        .din(new_Jinkela_wire_9610),
        .dout(new_Jinkela_wire_9611)
    );

    spl2 new_Jinkela_splitter_785 (
        .a(new_Jinkela_wire_9595),
        .b(new_Jinkela_wire_9596),
        .c(new_Jinkela_wire_9597)
    );

    and_bi n_1539_ (
        .a(new_Jinkela_wire_9020),
        .b(new_Jinkela_wire_7306),
        .c(n_0807_)
    );

    bfr new_Jinkela_buffer_8224 (
        .din(new_Jinkela_wire_10327),
        .dout(new_Jinkela_wire_10328)
    );

    and_bi n_1540_ (
        .a(new_Jinkela_wire_7305),
        .b(new_Jinkela_wire_9021),
        .c(n_0808_)
    );

    and_ii n_1541_ (
        .a(n_0808_),
        .b(n_0807_),
        .c(n_0809_)
    );

    bfr new_Jinkela_buffer_7639 (
        .din(new_Jinkela_wire_9608),
        .dout(new_Jinkela_wire_9609)
    );

    bfr new_Jinkela_buffer_8255 (
        .din(new_Jinkela_wire_10358),
        .dout(new_Jinkela_wire_10359)
    );

    bfr new_Jinkela_buffer_7648 (
        .din(n_0354_),
        .dout(new_Jinkela_wire_9621)
    );

    bfr new_Jinkela_buffer_8225 (
        .din(new_Jinkela_wire_10328),
        .dout(new_Jinkela_wire_10329)
    );

    and_bb n_1542_ (
        .a(new_Jinkela_wire_875),
        .b(new_Jinkela_wire_1326),
        .c(n_0810_)
    );

    bfr new_Jinkela_buffer_7642 (
        .din(new_Jinkela_wire_9611),
        .dout(new_Jinkela_wire_9612)
    );

    and_bi n_1543_ (
        .a(new_Jinkela_wire_3513),
        .b(new_Jinkela_wire_1292),
        .c(n_0811_)
    );

    bfr new_Jinkela_buffer_7664 (
        .din(n_1254_),
        .dout(new_Jinkela_wire_9641)
    );

    spl3L new_Jinkela_splitter_851 (
        .a(n_0720_),
        .d(new_Jinkela_wire_10387),
        .b(new_Jinkela_wire_10388),
        .c(new_Jinkela_wire_10389)
    );

    bfr new_Jinkela_buffer_8226 (
        .din(new_Jinkela_wire_10329),
        .dout(new_Jinkela_wire_10330)
    );

    and_ii n_1544_ (
        .a(new_Jinkela_wire_7082),
        .b(new_Jinkela_wire_9620),
        .c(n_0812_)
    );

    bfr new_Jinkela_buffer_7643 (
        .din(new_Jinkela_wire_9612),
        .dout(new_Jinkela_wire_9613)
    );

    bfr new_Jinkela_buffer_8262 (
        .din(new_Jinkela_wire_10374),
        .dout(new_Jinkela_wire_10375)
    );

    and_bi n_1545_ (
        .a(new_Jinkela_wire_7452),
        .b(new_Jinkela_wire_3938),
        .c(n_0813_)
    );

    bfr new_Jinkela_buffer_7665 (
        .din(n_0633_),
        .dout(new_Jinkela_wire_9644)
    );

    bfr new_Jinkela_buffer_8227 (
        .din(new_Jinkela_wire_10330),
        .dout(new_Jinkela_wire_10331)
    );

    and_bi n_1546_ (
        .a(new_Jinkela_wire_3936),
        .b(new_Jinkela_wire_7450),
        .c(n_0814_)
    );

    bfr new_Jinkela_buffer_7644 (
        .din(new_Jinkela_wire_9613),
        .dout(new_Jinkela_wire_9614)
    );

    spl2 new_Jinkela_splitter_854 (
        .a(n_0984_),
        .b(new_Jinkela_wire_10417),
        .c(new_Jinkela_wire_10418)
    );

    and_ii n_1547_ (
        .a(n_0814_),
        .b(n_0813_),
        .c(n_0815_)
    );

    spl4L new_Jinkela_splitter_855 (
        .a(n_1260_),
        .d(new_Jinkela_wire_10419),
        .b(new_Jinkela_wire_10420),
        .e(new_Jinkela_wire_10421),
        .c(new_Jinkela_wire_10422)
    );

    bfr new_Jinkela_buffer_7652 (
        .din(new_Jinkela_wire_9626),
        .dout(new_Jinkela_wire_9627)
    );

    bfr new_Jinkela_buffer_8228 (
        .din(new_Jinkela_wire_10331),
        .dout(new_Jinkela_wire_10332)
    );

    and_bi n_1548_ (
        .a(new_Jinkela_wire_4540),
        .b(new_Jinkela_wire_6191),
        .c(n_0816_)
    );

    bfr new_Jinkela_buffer_7645 (
        .din(new_Jinkela_wire_9614),
        .dout(new_Jinkela_wire_9615)
    );

    bfr new_Jinkela_buffer_8263 (
        .din(new_Jinkela_wire_10375),
        .dout(new_Jinkela_wire_10376)
    );

    and_bi n_1549_ (
        .a(new_Jinkela_wire_6190),
        .b(new_Jinkela_wire_4539),
        .c(n_0817_)
    );

    bfr new_Jinkela_buffer_7649 (
        .din(new_Jinkela_wire_9621),
        .dout(new_Jinkela_wire_9622)
    );

    bfr new_Jinkela_buffer_8229 (
        .din(new_Jinkela_wire_10332),
        .dout(new_Jinkela_wire_10333)
    );

    or_bb n_1550_ (
        .a(n_0817_),
        .b(n_0816_),
        .c(n_0818_)
    );

    bfr new_Jinkela_buffer_7646 (
        .din(new_Jinkela_wire_9615),
        .dout(new_Jinkela_wire_9616)
    );

    bfr new_Jinkela_buffer_8268 (
        .din(new_Jinkela_wire_10391),
        .dout(new_Jinkela_wire_10392)
    );

    and_bi n_1551_ (
        .a(new_Jinkela_wire_9748),
        .b(new_Jinkela_wire_9025),
        .c(n_0819_)
    );

    spl2 new_Jinkela_splitter_792 (
        .a(n_1258_),
        .b(new_Jinkela_wire_9642),
        .c(new_Jinkela_wire_9643)
    );

    bfr new_Jinkela_buffer_7668 (
        .din(n_1166_),
        .dout(new_Jinkela_wire_9649)
    );

    bfr new_Jinkela_buffer_8230 (
        .din(new_Jinkela_wire_10333),
        .dout(new_Jinkela_wire_10334)
    );

    and_bi n_1552_ (
        .a(new_Jinkela_wire_9023),
        .b(new_Jinkela_wire_9745),
        .c(n_0820_)
    );

    spl2 new_Jinkela_splitter_790 (
        .a(new_Jinkela_wire_9622),
        .b(new_Jinkela_wire_9623),
        .c(new_Jinkela_wire_9624)
    );

    bfr new_Jinkela_buffer_8264 (
        .din(new_Jinkela_wire_10376),
        .dout(new_Jinkela_wire_10377)
    );

    or_bb n_1553_ (
        .a(n_0820_),
        .b(n_0819_),
        .c(n_0821_)
    );

    bfr new_Jinkela_buffer_7650 (
        .din(new_Jinkela_wire_9624),
        .dout(new_Jinkela_wire_9625)
    );

    bfr new_Jinkela_buffer_8231 (
        .din(new_Jinkela_wire_10334),
        .dout(new_Jinkela_wire_10335)
    );

    or_ii n_1554_ (
        .a(new_Jinkela_wire_2735),
        .b(new_Jinkela_wire_1315),
        .c(n_0822_)
    );

    bfr new_Jinkela_buffer_7667 (
        .din(n_0225_),
        .dout(new_Jinkela_wire_9648)
    );

    and_bi n_1555_ (
        .a(new_Jinkela_wire_2478),
        .b(new_Jinkela_wire_1255),
        .c(n_0823_)
    );

    bfr new_Jinkela_buffer_7666 (
        .din(new_Jinkela_wire_9644),
        .dout(new_Jinkela_wire_9645)
    );

    bfr new_Jinkela_buffer_8305 (
        .din(n_0412_),
        .dout(new_Jinkela_wire_10443)
    );

    bfr new_Jinkela_buffer_8232 (
        .din(new_Jinkela_wire_10335),
        .dout(new_Jinkela_wire_10336)
    );

    and_bi n_1556_ (
        .a(new_Jinkela_wire_5249),
        .b(new_Jinkela_wire_10361),
        .c(n_0824_)
    );

    bfr new_Jinkela_buffer_7651 (
        .din(new_Jinkela_wire_9625),
        .dout(new_Jinkela_wire_9626)
    );

    or_ii n_1557_ (
        .a(new_Jinkela_wire_2662),
        .b(new_Jinkela_wire_1251),
        .c(n_0825_)
    );

    bfr new_Jinkela_buffer_8233 (
        .din(new_Jinkela_wire_10336),
        .dout(new_Jinkela_wire_10337)
    );

    and_bi n_1558_ (
        .a(new_Jinkela_wire_3438),
        .b(new_Jinkela_wire_1354),
        .c(n_0826_)
    );

    spl2 new_Jinkela_splitter_856 (
        .a(n_0028_),
        .b(new_Jinkela_wire_10423),
        .c(new_Jinkela_wire_10424)
    );

    and_bi n_1559_ (
        .a(new_Jinkela_wire_5368),
        .b(new_Jinkela_wire_9393),
        .c(n_0827_)
    );

    spl4L new_Jinkela_splitter_794 (
        .a(n_0116_),
        .d(new_Jinkela_wire_9650),
        .b(new_Jinkela_wire_9651),
        .e(new_Jinkela_wire_9652),
        .c(new_Jinkela_wire_9653)
    );

    bfr new_Jinkela_buffer_8269 (
        .din(new_Jinkela_wire_10392),
        .dout(new_Jinkela_wire_10393)
    );

    spl2 new_Jinkela_splitter_793 (
        .a(new_Jinkela_wire_9645),
        .b(new_Jinkela_wire_9646),
        .c(new_Jinkela_wire_9647)
    );

    bfr new_Jinkela_buffer_8234 (
        .din(new_Jinkela_wire_10337),
        .dout(new_Jinkela_wire_10338)
    );

    and_bi n_1560_ (
        .a(new_Jinkela_wire_9248),
        .b(new_Jinkela_wire_6841),
        .c(n_0828_)
    );

    bfr new_Jinkela_buffer_7653 (
        .din(new_Jinkela_wire_9627),
        .dout(new_Jinkela_wire_9628)
    );

    and_bi n_1561_ (
        .a(new_Jinkela_wire_6839),
        .b(new_Jinkela_wire_9247),
        .c(n_0829_)
    );

    bfr new_Jinkela_buffer_8235 (
        .din(new_Jinkela_wire_10338),
        .dout(new_Jinkela_wire_10339)
    );

    and_ii n_1562_ (
        .a(n_0829_),
        .b(n_0828_),
        .c(n_0830_)
    );

    bfr new_Jinkela_buffer_7654 (
        .din(new_Jinkela_wire_9628),
        .dout(new_Jinkela_wire_9629)
    );

    spl2 new_Jinkela_splitter_858 (
        .a(n_0047_),
        .b(new_Jinkela_wire_10433),
        .c(new_Jinkela_wire_10434)
    );

    and_bb n_1563_ (
        .a(new_Jinkela_wire_1613),
        .b(new_Jinkela_wire_1305),
        .c(n_0831_)
    );

    bfr new_Jinkela_buffer_8270 (
        .din(new_Jinkela_wire_10393),
        .dout(new_Jinkela_wire_10394)
    );

    spl2 new_Jinkela_splitter_798 (
        .a(n_1367_),
        .b(new_Jinkela_wire_9703),
        .c(new_Jinkela_wire_9705)
    );

    bfr new_Jinkela_buffer_8236 (
        .din(new_Jinkela_wire_10339),
        .dout(new_Jinkela_wire_10340)
    );

    and_bi n_1564_ (
        .a(new_Jinkela_wire_584),
        .b(new_Jinkela_wire_1181),
        .c(n_0832_)
    );

    bfr new_Jinkela_buffer_7655 (
        .din(new_Jinkela_wire_9629),
        .dout(new_Jinkela_wire_9630)
    );

    and_ii n_1565_ (
        .a(new_Jinkela_wire_5068),
        .b(new_Jinkela_wire_6323),
        .c(n_0833_)
    );

    bfr new_Jinkela_buffer_7713 (
        .din(n_0465_),
        .dout(new_Jinkela_wire_9710)
    );

    bfr new_Jinkela_buffer_8296 (
        .din(n_0381_),
        .dout(new_Jinkela_wire_10432)
    );

    and_bi n_1566_ (
        .a(new_Jinkela_wire_5875),
        .b(new_Jinkela_wire_7264),
        .c(n_0834_)
    );

    bfr new_Jinkela_buffer_7656 (
        .din(new_Jinkela_wire_9630),
        .dout(new_Jinkela_wire_9631)
    );

    bfr new_Jinkela_buffer_8271 (
        .din(new_Jinkela_wire_10394),
        .dout(new_Jinkela_wire_10395)
    );

    and_bi n_1567_ (
        .a(new_Jinkela_wire_7267),
        .b(new_Jinkela_wire_5874),
        .c(n_0835_)
    );

    bfr new_Jinkela_buffer_7669 (
        .din(new_Jinkela_wire_9653),
        .dout(new_Jinkela_wire_9654)
    );

    bfr new_Jinkela_buffer_8291 (
        .din(new_Jinkela_wire_10424),
        .dout(new_Jinkela_wire_10425)
    );

    and_ii n_1568_ (
        .a(n_0835_),
        .b(n_0834_),
        .c(n_0836_)
    );

    bfr new_Jinkela_buffer_7657 (
        .din(new_Jinkela_wire_9631),
        .dout(new_Jinkela_wire_9632)
    );

    bfr new_Jinkela_buffer_8272 (
        .din(new_Jinkela_wire_10395),
        .dout(new_Jinkela_wire_10396)
    );

    bfr new_Jinkela_buffer_813 (
        .din(new_Jinkela_wire_873),
        .dout(new_Jinkela_wire_874)
    );

    bfr new_Jinkela_buffer_4590 (
        .din(new_Jinkela_wire_5468),
        .dout(new_Jinkela_wire_5469)
    );

    bfr new_Jinkela_buffer_695 (
        .din(new_Jinkela_wire_747),
        .dout(new_Jinkela_wire_748)
    );

    bfr new_Jinkela_buffer_7067 (
        .din(new_Jinkela_wire_8731),
        .dout(new_Jinkela_wire_8732)
    );

    bfr new_Jinkela_buffer_4575 (
        .din(new_Jinkela_wire_5447),
        .dout(new_Jinkela_wire_5448)
    );

    bfr new_Jinkela_buffer_749 (
        .din(new_Jinkela_wire_809),
        .dout(new_Jinkela_wire_810)
    );

    bfr new_Jinkela_buffer_7126 (
        .din(new_Jinkela_wire_8814),
        .dout(new_Jinkela_wire_8815)
    );

    spl3L new_Jinkela_splitter_678 (
        .a(n_1349_),
        .d(new_Jinkela_wire_8843),
        .b(new_Jinkela_wire_8844),
        .c(new_Jinkela_wire_8845)
    );

    bfr new_Jinkela_buffer_696 (
        .din(new_Jinkela_wire_748),
        .dout(new_Jinkela_wire_749)
    );

    bfr new_Jinkela_buffer_7068 (
        .din(new_Jinkela_wire_8732),
        .dout(new_Jinkela_wire_8733)
    );

    bfr new_Jinkela_buffer_4591 (
        .din(new_Jinkela_wire_5469),
        .dout(new_Jinkela_wire_5470)
    );

    bfr new_Jinkela_buffer_816 (
        .din(new_Jinkela_wire_876),
        .dout(new_Jinkela_wire_877)
    );

    bfr new_Jinkela_buffer_7086 (
        .din(new_Jinkela_wire_8769),
        .dout(new_Jinkela_wire_8770)
    );

    bfr new_Jinkela_buffer_697 (
        .din(new_Jinkela_wire_749),
        .dout(new_Jinkela_wire_750)
    );

    bfr new_Jinkela_buffer_4628 (
        .din(new_Jinkela_wire_5508),
        .dout(new_Jinkela_wire_5509)
    );

    bfr new_Jinkela_buffer_7069 (
        .din(new_Jinkela_wire_8733),
        .dout(new_Jinkela_wire_8734)
    );

    bfr new_Jinkela_buffer_4592 (
        .din(new_Jinkela_wire_5470),
        .dout(new_Jinkela_wire_5471)
    );

    bfr new_Jinkela_buffer_750 (
        .din(new_Jinkela_wire_810),
        .dout(new_Jinkela_wire_811)
    );

    spl2 new_Jinkela_splitter_677 (
        .a(n_1057_),
        .b(new_Jinkela_wire_8821),
        .c(new_Jinkela_wire_8822)
    );

    bfr new_Jinkela_buffer_698 (
        .din(new_Jinkela_wire_750),
        .dout(new_Jinkela_wire_751)
    );

    spl3L new_Jinkela_splitter_334 (
        .a(n_0700_),
        .d(new_Jinkela_wire_5560),
        .b(new_Jinkela_wire_5561),
        .c(new_Jinkela_wire_5562)
    );

    bfr new_Jinkela_buffer_7070 (
        .din(new_Jinkela_wire_8734),
        .dout(new_Jinkela_wire_8735)
    );

    bfr new_Jinkela_buffer_4593 (
        .din(new_Jinkela_wire_5471),
        .dout(new_Jinkela_wire_5472)
    );

    bfr new_Jinkela_buffer_814 (
        .din(new_Jinkela_wire_874),
        .dout(new_Jinkela_wire_875)
    );

    bfr new_Jinkela_buffer_7087 (
        .din(new_Jinkela_wire_8770),
        .dout(new_Jinkela_wire_8771)
    );

    spl2 new_Jinkela_splitter_333 (
        .a(new_Jinkela_wire_5556),
        .b(new_Jinkela_wire_5557),
        .c(new_Jinkela_wire_5558)
    );

    bfr new_Jinkela_buffer_699 (
        .din(new_Jinkela_wire_751),
        .dout(new_Jinkela_wire_752)
    );

    bfr new_Jinkela_buffer_4629 (
        .din(new_Jinkela_wire_5509),
        .dout(new_Jinkela_wire_5510)
    );

    bfr new_Jinkela_buffer_7071 (
        .din(new_Jinkela_wire_8735),
        .dout(new_Jinkela_wire_8736)
    );

    bfr new_Jinkela_buffer_4594 (
        .din(new_Jinkela_wire_5472),
        .dout(new_Jinkela_wire_5473)
    );

    bfr new_Jinkela_buffer_751 (
        .din(new_Jinkela_wire_811),
        .dout(new_Jinkela_wire_812)
    );

    bfr new_Jinkela_buffer_7128 (
        .din(n_1245_),
        .dout(new_Jinkela_wire_8823)
    );

    bfr new_Jinkela_buffer_700 (
        .din(new_Jinkela_wire_752),
        .dout(new_Jinkela_wire_753)
    );

    bfr new_Jinkela_buffer_7072 (
        .din(new_Jinkela_wire_8736),
        .dout(new_Jinkela_wire_8737)
    );

    bfr new_Jinkela_buffer_4595 (
        .din(new_Jinkela_wire_5473),
        .dout(new_Jinkela_wire_5474)
    );

    bfr new_Jinkela_buffer_7088 (
        .din(new_Jinkela_wire_8771),
        .dout(new_Jinkela_wire_8772)
    );

    spl3L new_Jinkela_splitter_337 (
        .a(n_0104_),
        .d(new_Jinkela_wire_5569),
        .b(new_Jinkela_wire_5570),
        .c(new_Jinkela_wire_5571)
    );

    bfr new_Jinkela_buffer_7073 (
        .din(new_Jinkela_wire_8737),
        .dout(new_Jinkela_wire_8738)
    );

    bfr new_Jinkela_buffer_701 (
        .din(new_Jinkela_wire_753),
        .dout(new_Jinkela_wire_754)
    );

    bfr new_Jinkela_buffer_4630 (
        .din(new_Jinkela_wire_5510),
        .dout(new_Jinkela_wire_5511)
    );

    bfr new_Jinkela_buffer_4596 (
        .din(new_Jinkela_wire_5474),
        .dout(new_Jinkela_wire_5475)
    );

    spl2 new_Jinkela_splitter_675 (
        .a(new_Jinkela_wire_8815),
        .b(new_Jinkela_wire_8816),
        .c(new_Jinkela_wire_8817)
    );

    bfr new_Jinkela_buffer_752 (
        .din(new_Jinkela_wire_812),
        .dout(new_Jinkela_wire_813)
    );

    bfr new_Jinkela_buffer_7074 (
        .din(new_Jinkela_wire_8738),
        .dout(new_Jinkela_wire_8739)
    );

    bfr new_Jinkela_buffer_702 (
        .din(new_Jinkela_wire_754),
        .dout(new_Jinkela_wire_755)
    );

    bfr new_Jinkela_buffer_4597 (
        .din(new_Jinkela_wire_5475),
        .dout(new_Jinkela_wire_5476)
    );

    bfr new_Jinkela_buffer_7089 (
        .din(new_Jinkela_wire_8772),
        .dout(new_Jinkela_wire_8773)
    );

    bfr new_Jinkela_buffer_817 (
        .din(new_Jinkela_wire_877),
        .dout(new_Jinkela_wire_878)
    );

    spl2 new_Jinkela_splitter_336 (
        .a(n_0149_),
        .b(new_Jinkela_wire_5567),
        .c(new_Jinkela_wire_5568)
    );

    bfr new_Jinkela_buffer_7075 (
        .din(new_Jinkela_wire_8739),
        .dout(new_Jinkela_wire_8740)
    );

    bfr new_Jinkela_buffer_703 (
        .din(new_Jinkela_wire_755),
        .dout(new_Jinkela_wire_756)
    );

    bfr new_Jinkela_buffer_4631 (
        .din(new_Jinkela_wire_5511),
        .dout(new_Jinkela_wire_5512)
    );

    bfr new_Jinkela_buffer_4598 (
        .din(new_Jinkela_wire_5476),
        .dout(new_Jinkela_wire_5477)
    );

    bfr new_Jinkela_buffer_753 (
        .din(new_Jinkela_wire_813),
        .dout(new_Jinkela_wire_814)
    );

    spl2 new_Jinkela_splitter_676 (
        .a(new_Jinkela_wire_8817),
        .b(new_Jinkela_wire_8818),
        .c(new_Jinkela_wire_8819)
    );

    bfr new_Jinkela_buffer_7076 (
        .din(new_Jinkela_wire_8740),
        .dout(new_Jinkela_wire_8741)
    );

    bfr new_Jinkela_buffer_704 (
        .din(new_Jinkela_wire_756),
        .dout(new_Jinkela_wire_757)
    );

    spl2 new_Jinkela_splitter_339 (
        .a(n_0906_),
        .b(new_Jinkela_wire_5575),
        .c(new_Jinkela_wire_5576)
    );

    bfr new_Jinkela_buffer_4599 (
        .din(new_Jinkela_wire_5477),
        .dout(new_Jinkela_wire_5478)
    );

    bfr new_Jinkela_buffer_7090 (
        .din(new_Jinkela_wire_8773),
        .dout(new_Jinkela_wire_8774)
    );

    bfr new_Jinkela_buffer_947 (
        .din(new_Jinkela_wire_1019),
        .dout(new_Jinkela_wire_1020)
    );

    bfr new_Jinkela_buffer_1011 (
        .din(N232),
        .dout(new_Jinkela_wire_1086)
    );

    bfr new_Jinkela_buffer_4677 (
        .din(new_Jinkela_wire_5564),
        .dout(new_Jinkela_wire_5565)
    );

    bfr new_Jinkela_buffer_7077 (
        .din(new_Jinkela_wire_8741),
        .dout(new_Jinkela_wire_8742)
    );

    bfr new_Jinkela_buffer_705 (
        .din(new_Jinkela_wire_757),
        .dout(new_Jinkela_wire_758)
    );

    bfr new_Jinkela_buffer_4632 (
        .din(new_Jinkela_wire_5512),
        .dout(new_Jinkela_wire_5513)
    );

    bfr new_Jinkela_buffer_4600 (
        .din(new_Jinkela_wire_5478),
        .dout(new_Jinkela_wire_5479)
    );

    bfr new_Jinkela_buffer_754 (
        .din(new_Jinkela_wire_814),
        .dout(new_Jinkela_wire_815)
    );

    bfr new_Jinkela_buffer_7078 (
        .din(new_Jinkela_wire_8742),
        .dout(new_Jinkela_wire_8743)
    );

    bfr new_Jinkela_buffer_818 (
        .din(new_Jinkela_wire_878),
        .dout(new_Jinkela_wire_879)
    );

    spl2 new_Jinkela_splitter_335 (
        .a(new_Jinkela_wire_5562),
        .b(new_Jinkela_wire_5563),
        .c(new_Jinkela_wire_5564)
    );

    bfr new_Jinkela_buffer_4601 (
        .din(new_Jinkela_wire_5479),
        .dout(new_Jinkela_wire_5480)
    );

    bfr new_Jinkela_buffer_7091 (
        .din(new_Jinkela_wire_8774),
        .dout(new_Jinkela_wire_8775)
    );

    bfr new_Jinkela_buffer_755 (
        .din(new_Jinkela_wire_815),
        .dout(new_Jinkela_wire_816)
    );

    bfr new_Jinkela_buffer_7079 (
        .din(new_Jinkela_wire_8743),
        .dout(new_Jinkela_wire_8744)
    );

    bfr new_Jinkela_buffer_4633 (
        .din(new_Jinkela_wire_5513),
        .dout(new_Jinkela_wire_5514)
    );

    bfr new_Jinkela_buffer_4602 (
        .din(new_Jinkela_wire_5480),
        .dout(new_Jinkela_wire_5481)
    );

    bfr new_Jinkela_buffer_7129 (
        .din(n_0068_),
        .dout(new_Jinkela_wire_8824)
    );

    bfr new_Jinkela_buffer_756 (
        .din(new_Jinkela_wire_816),
        .dout(new_Jinkela_wire_817)
    );

    bfr new_Jinkela_buffer_7080 (
        .din(new_Jinkela_wire_8744),
        .dout(new_Jinkela_wire_8745)
    );

    bfr new_Jinkela_buffer_821 (
        .din(new_Jinkela_wire_881),
        .dout(new_Jinkela_wire_882)
    );

    bfr new_Jinkela_buffer_4603 (
        .din(new_Jinkela_wire_5481),
        .dout(new_Jinkela_wire_5482)
    );

    bfr new_Jinkela_buffer_7092 (
        .din(new_Jinkela_wire_8775),
        .dout(new_Jinkela_wire_8776)
    );

    bfr new_Jinkela_buffer_757 (
        .din(new_Jinkela_wire_817),
        .dout(new_Jinkela_wire_818)
    );

    bfr new_Jinkela_buffer_7081 (
        .din(new_Jinkela_wire_8745),
        .dout(new_Jinkela_wire_8746)
    );

    bfr new_Jinkela_buffer_4634 (
        .din(new_Jinkela_wire_5514),
        .dout(new_Jinkela_wire_5515)
    );

    bfr new_Jinkela_buffer_820 (
        .din(new_Jinkela_wire_880),
        .dout(new_Jinkela_wire_881)
    );

    bfr new_Jinkela_buffer_4604 (
        .din(new_Jinkela_wire_5482),
        .dout(new_Jinkela_wire_5483)
    );

    bfr new_Jinkela_buffer_7151 (
        .din(n_0529_),
        .dout(new_Jinkela_wire_8853)
    );

    bfr new_Jinkela_buffer_758 (
        .din(new_Jinkela_wire_818),
        .dout(new_Jinkela_wire_819)
    );

    bfr new_Jinkela_buffer_7148 (
        .din(n_0597_),
        .dout(new_Jinkela_wire_8848)
    );

    bfr new_Jinkela_buffer_7093 (
        .din(new_Jinkela_wire_8776),
        .dout(new_Jinkela_wire_8777)
    );

    spl2 new_Jinkela_splitter_27 (
        .a(new_Jinkela_wire_882),
        .b(new_Jinkela_wire_883),
        .c(new_Jinkela_wire_884)
    );

    bfr new_Jinkela_buffer_4605 (
        .din(new_Jinkela_wire_5483),
        .dout(new_Jinkela_wire_5484)
    );

    bfr new_Jinkela_buffer_7130 (
        .din(new_Jinkela_wire_8824),
        .dout(new_Jinkela_wire_8825)
    );

    bfr new_Jinkela_buffer_759 (
        .din(new_Jinkela_wire_819),
        .dout(new_Jinkela_wire_820)
    );

    bfr new_Jinkela_buffer_4679 (
        .din(n_0609_),
        .dout(new_Jinkela_wire_5572)
    );

    bfr new_Jinkela_buffer_7094 (
        .din(new_Jinkela_wire_8777),
        .dout(new_Jinkela_wire_8778)
    );

    bfr new_Jinkela_buffer_822 (
        .din(new_Jinkela_wire_884),
        .dout(new_Jinkela_wire_885)
    );

    bfr new_Jinkela_buffer_4635 (
        .din(new_Jinkela_wire_5515),
        .dout(new_Jinkela_wire_5516)
    );

    bfr new_Jinkela_buffer_4606 (
        .din(new_Jinkela_wire_5484),
        .dout(new_Jinkela_wire_5485)
    );

    bfr new_Jinkela_buffer_7131 (
        .din(new_Jinkela_wire_8825),
        .dout(new_Jinkela_wire_8826)
    );

    bfr new_Jinkela_buffer_760 (
        .din(new_Jinkela_wire_820),
        .dout(new_Jinkela_wire_821)
    );

    bfr new_Jinkela_buffer_7095 (
        .din(new_Jinkela_wire_8778),
        .dout(new_Jinkela_wire_8779)
    );

    bfr new_Jinkela_buffer_4607 (
        .din(new_Jinkela_wire_5485),
        .dout(new_Jinkela_wire_5486)
    );

    bfr new_Jinkela_buffer_761 (
        .din(new_Jinkela_wire_821),
        .dout(new_Jinkela_wire_822)
    );

    spl2 new_Jinkela_splitter_338 (
        .a(n_0869_),
        .b(new_Jinkela_wire_5573),
        .c(new_Jinkela_wire_5574)
    );

    bfr new_Jinkela_buffer_7096 (
        .din(new_Jinkela_wire_8779),
        .dout(new_Jinkela_wire_8780)
    );

    bfr new_Jinkela_buffer_4636 (
        .din(new_Jinkela_wire_5516),
        .dout(new_Jinkela_wire_5517)
    );

    bfr new_Jinkela_buffer_884 (
        .din(new_Jinkela_wire_949),
        .dout(new_Jinkela_wire_950)
    );

    bfr new_Jinkela_buffer_4608 (
        .din(new_Jinkela_wire_5486),
        .dout(new_Jinkela_wire_5487)
    );

    bfr new_Jinkela_buffer_7132 (
        .din(new_Jinkela_wire_8826),
        .dout(new_Jinkela_wire_8827)
    );

    bfr new_Jinkela_buffer_762 (
        .din(new_Jinkela_wire_822),
        .dout(new_Jinkela_wire_823)
    );

    bfr new_Jinkela_buffer_7097 (
        .din(new_Jinkela_wire_8780),
        .dout(new_Jinkela_wire_8781)
    );

    bfr new_Jinkela_buffer_885 (
        .din(new_Jinkela_wire_950),
        .dout(new_Jinkela_wire_951)
    );

    bfr new_Jinkela_buffer_4678 (
        .din(new_Jinkela_wire_5565),
        .dout(new_Jinkela_wire_5566)
    );

    spl2 new_Jinkela_splitter_31 (
        .a(N364),
        .b(new_Jinkela_wire_1018),
        .c(new_Jinkela_wire_1019)
    );

    bfr new_Jinkela_buffer_4609 (
        .din(new_Jinkela_wire_5487),
        .dout(new_Jinkela_wire_5488)
    );

    spl2 new_Jinkela_splitter_679 (
        .a(new_Jinkela_wire_8845),
        .b(new_Jinkela_wire_8846),
        .c(new_Jinkela_wire_8847)
    );

    bfr new_Jinkela_buffer_763 (
        .din(new_Jinkela_wire_823),
        .dout(new_Jinkela_wire_824)
    );

    spl2 new_Jinkela_splitter_680 (
        .a(n_0302_),
        .b(new_Jinkela_wire_8850),
        .c(new_Jinkela_wire_8851)
    );

    bfr new_Jinkela_buffer_7098 (
        .din(new_Jinkela_wire_8781),
        .dout(new_Jinkela_wire_8782)
    );

    bfr new_Jinkela_buffer_823 (
        .din(new_Jinkela_wire_885),
        .dout(new_Jinkela_wire_886)
    );

    bfr new_Jinkela_buffer_4637 (
        .din(new_Jinkela_wire_5517),
        .dout(new_Jinkela_wire_5518)
    );

    bfr new_Jinkela_buffer_4610 (
        .din(new_Jinkela_wire_5488),
        .dout(new_Jinkela_wire_5489)
    );

    bfr new_Jinkela_buffer_7133 (
        .din(new_Jinkela_wire_8827),
        .dout(new_Jinkela_wire_8828)
    );

    bfr new_Jinkela_buffer_1137 (
        .din(new_Jinkela_wire_1448),
        .dout(new_Jinkela_wire_1449)
    );

    bfr new_Jinkela_buffer_6246 (
        .din(new_Jinkela_wire_7619),
        .dout(new_Jinkela_wire_7620)
    );

    spl2 new_Jinkela_splitter_100 (
        .a(new_Jinkela_wire_1616),
        .b(new_Jinkela_wire_1617),
        .c(new_Jinkela_wire_1618)
    );

    bfr new_Jinkela_buffer_6291 (
        .din(new_Jinkela_wire_7668),
        .dout(new_Jinkela_wire_7669)
    );

    bfr new_Jinkela_buffer_1138 (
        .din(new_Jinkela_wire_1449),
        .dout(new_Jinkela_wire_1450)
    );

    bfr new_Jinkela_buffer_6247 (
        .din(new_Jinkela_wire_7620),
        .dout(new_Jinkela_wire_7621)
    );

    bfr new_Jinkela_buffer_1180 (
        .din(new_Jinkela_wire_1496),
        .dout(new_Jinkela_wire_1497)
    );

    bfr new_Jinkela_buffer_6351 (
        .din(new_Jinkela_wire_7736),
        .dout(new_Jinkela_wire_7737)
    );

    bfr new_Jinkela_buffer_1139 (
        .din(new_Jinkela_wire_1450),
        .dout(new_Jinkela_wire_1451)
    );

    bfr new_Jinkela_buffer_6248 (
        .din(new_Jinkela_wire_7621),
        .dout(new_Jinkela_wire_7622)
    );

    bfr new_Jinkela_buffer_1233 (
        .din(new_Jinkela_wire_1553),
        .dout(new_Jinkela_wire_1554)
    );

    bfr new_Jinkela_buffer_6292 (
        .din(new_Jinkela_wire_7669),
        .dout(new_Jinkela_wire_7670)
    );

    bfr new_Jinkela_buffer_1140 (
        .din(new_Jinkela_wire_1451),
        .dout(new_Jinkela_wire_1452)
    );

    bfr new_Jinkela_buffer_6249 (
        .din(new_Jinkela_wire_7622),
        .dout(new_Jinkela_wire_7623)
    );

    bfr new_Jinkela_buffer_1181 (
        .din(new_Jinkela_wire_1497),
        .dout(new_Jinkela_wire_1498)
    );

    bfr new_Jinkela_buffer_6313 (
        .din(new_Jinkela_wire_7694),
        .dout(new_Jinkela_wire_7695)
    );

    bfr new_Jinkela_buffer_1141 (
        .din(new_Jinkela_wire_1452),
        .dout(new_Jinkela_wire_1453)
    );

    bfr new_Jinkela_buffer_6250 (
        .din(new_Jinkela_wire_7623),
        .dout(new_Jinkela_wire_7624)
    );

    bfr new_Jinkela_buffer_1296 (
        .din(new_Jinkela_wire_1618),
        .dout(new_Jinkela_wire_1619)
    );

    bfr new_Jinkela_buffer_6293 (
        .din(new_Jinkela_wire_7670),
        .dout(new_Jinkela_wire_7671)
    );

    bfr new_Jinkela_buffer_1142 (
        .din(new_Jinkela_wire_1453),
        .dout(new_Jinkela_wire_1454)
    );

    bfr new_Jinkela_buffer_6251 (
        .din(new_Jinkela_wire_7624),
        .dout(new_Jinkela_wire_7625)
    );

    bfr new_Jinkela_buffer_1182 (
        .din(new_Jinkela_wire_1498),
        .dout(new_Jinkela_wire_1499)
    );

    bfr new_Jinkela_buffer_6348 (
        .din(new_Jinkela_wire_7733),
        .dout(new_Jinkela_wire_7734)
    );

    bfr new_Jinkela_buffer_1143 (
        .din(new_Jinkela_wire_1454),
        .dout(new_Jinkela_wire_1455)
    );

    bfr new_Jinkela_buffer_6252 (
        .din(new_Jinkela_wire_7625),
        .dout(new_Jinkela_wire_7626)
    );

    bfr new_Jinkela_buffer_1234 (
        .din(new_Jinkela_wire_1554),
        .dout(new_Jinkela_wire_1555)
    );

    bfr new_Jinkela_buffer_6294 (
        .din(new_Jinkela_wire_7671),
        .dout(new_Jinkela_wire_7672)
    );

    bfr new_Jinkela_buffer_1144 (
        .din(new_Jinkela_wire_1455),
        .dout(new_Jinkela_wire_1456)
    );

    bfr new_Jinkela_buffer_6253 (
        .din(new_Jinkela_wire_7626),
        .dout(new_Jinkela_wire_7627)
    );

    bfr new_Jinkela_buffer_1183 (
        .din(new_Jinkela_wire_1499),
        .dout(new_Jinkela_wire_1500)
    );

    bfr new_Jinkela_buffer_6314 (
        .din(new_Jinkela_wire_7695),
        .dout(new_Jinkela_wire_7696)
    );

    bfr new_Jinkela_buffer_1145 (
        .din(new_Jinkela_wire_1456),
        .dout(new_Jinkela_wire_1457)
    );

    bfr new_Jinkela_buffer_6254 (
        .din(new_Jinkela_wire_7627),
        .dout(new_Jinkela_wire_7628)
    );

    bfr new_Jinkela_buffer_1365 (
        .din(N29),
        .dout(new_Jinkela_wire_1691)
    );

    bfr new_Jinkela_buffer_6295 (
        .din(new_Jinkela_wire_7672),
        .dout(new_Jinkela_wire_7673)
    );

    bfr new_Jinkela_buffer_1146 (
        .din(new_Jinkela_wire_1457),
        .dout(new_Jinkela_wire_1458)
    );

    bfr new_Jinkela_buffer_6255 (
        .din(new_Jinkela_wire_7628),
        .dout(new_Jinkela_wire_7629)
    );

    bfr new_Jinkela_buffer_1184 (
        .din(new_Jinkela_wire_1500),
        .dout(new_Jinkela_wire_1501)
    );

    bfr new_Jinkela_buffer_6353 (
        .din(n_0459_),
        .dout(new_Jinkela_wire_7741)
    );

    spl3L new_Jinkela_splitter_548 (
        .a(n_1134_),
        .d(new_Jinkela_wire_7744),
        .b(new_Jinkela_wire_7745),
        .c(new_Jinkela_wire_7746)
    );

    bfr new_Jinkela_buffer_1147 (
        .din(new_Jinkela_wire_1458),
        .dout(new_Jinkela_wire_1459)
    );

    bfr new_Jinkela_buffer_6256 (
        .din(new_Jinkela_wire_7629),
        .dout(new_Jinkela_wire_7630)
    );

    bfr new_Jinkela_buffer_1235 (
        .din(new_Jinkela_wire_1555),
        .dout(new_Jinkela_wire_1556)
    );

    bfr new_Jinkela_buffer_6296 (
        .din(new_Jinkela_wire_7673),
        .dout(new_Jinkela_wire_7674)
    );

    bfr new_Jinkela_buffer_1148 (
        .din(new_Jinkela_wire_1459),
        .dout(new_Jinkela_wire_1460)
    );

    bfr new_Jinkela_buffer_6257 (
        .din(new_Jinkela_wire_7630),
        .dout(new_Jinkela_wire_7631)
    );

    bfr new_Jinkela_buffer_1185 (
        .din(new_Jinkela_wire_1501),
        .dout(new_Jinkela_wire_1502)
    );

    bfr new_Jinkela_buffer_6315 (
        .din(new_Jinkela_wire_7696),
        .dout(new_Jinkela_wire_7697)
    );

    bfr new_Jinkela_buffer_1149 (
        .din(new_Jinkela_wire_1460),
        .dout(new_Jinkela_wire_1461)
    );

    bfr new_Jinkela_buffer_6258 (
        .din(new_Jinkela_wire_7631),
        .dout(new_Jinkela_wire_7632)
    );

    bfr new_Jinkela_buffer_1359 (
        .din(new_Jinkela_wire_1684),
        .dout(new_Jinkela_wire_1685)
    );

    bfr new_Jinkela_buffer_6297 (
        .din(new_Jinkela_wire_7674),
        .dout(new_Jinkela_wire_7675)
    );

    bfr new_Jinkela_buffer_1150 (
        .din(new_Jinkela_wire_1461),
        .dout(new_Jinkela_wire_1462)
    );

    bfr new_Jinkela_buffer_6259 (
        .din(new_Jinkela_wire_7632),
        .dout(new_Jinkela_wire_7633)
    );

    bfr new_Jinkela_buffer_1186 (
        .din(new_Jinkela_wire_1502),
        .dout(new_Jinkela_wire_1503)
    );

    bfr new_Jinkela_buffer_6349 (
        .din(new_Jinkela_wire_7734),
        .dout(new_Jinkela_wire_7735)
    );

    bfr new_Jinkela_buffer_1151 (
        .din(new_Jinkela_wire_1462),
        .dout(new_Jinkela_wire_1463)
    );

    bfr new_Jinkela_buffer_6260 (
        .din(new_Jinkela_wire_7633),
        .dout(new_Jinkela_wire_7634)
    );

    bfr new_Jinkela_buffer_1236 (
        .din(new_Jinkela_wire_1556),
        .dout(new_Jinkela_wire_1557)
    );

    bfr new_Jinkela_buffer_6298 (
        .din(new_Jinkela_wire_7675),
        .dout(new_Jinkela_wire_7676)
    );

    bfr new_Jinkela_buffer_1152 (
        .din(new_Jinkela_wire_1463),
        .dout(new_Jinkela_wire_1464)
    );

    bfr new_Jinkela_buffer_6261 (
        .din(new_Jinkela_wire_7634),
        .dout(new_Jinkela_wire_7635)
    );

    bfr new_Jinkela_buffer_1187 (
        .din(new_Jinkela_wire_1503),
        .dout(new_Jinkela_wire_1504)
    );

    bfr new_Jinkela_buffer_6316 (
        .din(new_Jinkela_wire_7697),
        .dout(new_Jinkela_wire_7698)
    );

    bfr new_Jinkela_buffer_1153 (
        .din(new_Jinkela_wire_1464),
        .dout(new_Jinkela_wire_1465)
    );

    bfr new_Jinkela_buffer_6262 (
        .din(new_Jinkela_wire_7635),
        .dout(new_Jinkela_wire_7636)
    );

    bfr new_Jinkela_buffer_1362 (
        .din(new_Jinkela_wire_1687),
        .dout(new_Jinkela_wire_1688)
    );

    bfr new_Jinkela_buffer_6299 (
        .din(new_Jinkela_wire_7676),
        .dout(new_Jinkela_wire_7677)
    );

    bfr new_Jinkela_buffer_1154 (
        .din(new_Jinkela_wire_1465),
        .dout(new_Jinkela_wire_1466)
    );

    bfr new_Jinkela_buffer_6263 (
        .din(new_Jinkela_wire_7636),
        .dout(new_Jinkela_wire_7637)
    );

    bfr new_Jinkela_buffer_1188 (
        .din(new_Jinkela_wire_1504),
        .dout(new_Jinkela_wire_1505)
    );

    bfr new_Jinkela_buffer_6352 (
        .din(new_Jinkela_wire_7737),
        .dout(new_Jinkela_wire_7738)
    );

    bfr new_Jinkela_buffer_1155 (
        .din(new_Jinkela_wire_1466),
        .dout(new_Jinkela_wire_1467)
    );

    bfr new_Jinkela_buffer_6264 (
        .din(new_Jinkela_wire_7637),
        .dout(new_Jinkela_wire_7638)
    );

    bfr new_Jinkela_buffer_1237 (
        .din(new_Jinkela_wire_1557),
        .dout(new_Jinkela_wire_1558)
    );

    bfr new_Jinkela_buffer_6300 (
        .din(new_Jinkela_wire_7677),
        .dout(new_Jinkela_wire_7678)
    );

    bfr new_Jinkela_buffer_1156 (
        .din(new_Jinkela_wire_1467),
        .dout(new_Jinkela_wire_1468)
    );

    bfr new_Jinkela_buffer_6265 (
        .din(new_Jinkela_wire_7638),
        .dout(new_Jinkela_wire_7639)
    );

    bfr new_Jinkela_buffer_1189 (
        .din(new_Jinkela_wire_1505),
        .dout(new_Jinkela_wire_1506)
    );

    bfr new_Jinkela_buffer_6317 (
        .din(new_Jinkela_wire_7698),
        .dout(new_Jinkela_wire_7699)
    );

    bfr new_Jinkela_buffer_1157 (
        .din(new_Jinkela_wire_1468),
        .dout(new_Jinkela_wire_1469)
    );

    bfr new_Jinkela_buffer_6266 (
        .din(new_Jinkela_wire_7639),
        .dout(new_Jinkela_wire_7640)
    );

    bfr new_Jinkela_buffer_1297 (
        .din(new_Jinkela_wire_1619),
        .dout(new_Jinkela_wire_1620)
    );

    bfr new_Jinkela_buffer_6301 (
        .din(new_Jinkela_wire_7678),
        .dout(new_Jinkela_wire_7679)
    );

    bfr new_Jinkela_buffer_2947 (
        .din(new_Jinkela_wire_3374),
        .dout(new_Jinkela_wire_3375)
    );

    bfr new_Jinkela_buffer_1116 (
        .din(new_Jinkela_wire_1427),
        .dout(new_Jinkela_wire_1428)
    );

    bfr new_Jinkela_buffer_2894 (
        .din(new_Jinkela_wire_3317),
        .dout(new_Jinkela_wire_3318)
    );

    bfr new_Jinkela_buffer_1169 (
        .din(new_Jinkela_wire_1485),
        .dout(new_Jinkela_wire_1486)
    );

    bfr new_Jinkela_buffer_3796 (
        .din(new_Jinkela_wire_4418),
        .dout(new_Jinkela_wire_4419)
    );

    bfr new_Jinkela_buffer_3751 (
        .din(new_Jinkela_wire_4371),
        .dout(new_Jinkela_wire_4372)
    );

    bfr new_Jinkela_buffer_1117 (
        .din(new_Jinkela_wire_1428),
        .dout(new_Jinkela_wire_1429)
    );

    bfr new_Jinkela_buffer_2895 (
        .din(new_Jinkela_wire_3318),
        .dout(new_Jinkela_wire_3319)
    );

    bfr new_Jinkela_buffer_1361 (
        .din(N202),
        .dout(new_Jinkela_wire_1687)
    );

    bfr new_Jinkela_buffer_3752 (
        .din(new_Jinkela_wire_4372),
        .dout(new_Jinkela_wire_4373)
    );

    bfr new_Jinkela_buffer_2948 (
        .din(new_Jinkela_wire_3375),
        .dout(new_Jinkela_wire_3376)
    );

    bfr new_Jinkela_buffer_1118 (
        .din(new_Jinkela_wire_1429),
        .dout(new_Jinkela_wire_1430)
    );

    bfr new_Jinkela_buffer_3852 (
        .din(n_0147_),
        .dout(new_Jinkela_wire_4486)
    );

    bfr new_Jinkela_buffer_2896 (
        .din(new_Jinkela_wire_3319),
        .dout(new_Jinkela_wire_3320)
    );

    bfr new_Jinkela_buffer_1170 (
        .din(new_Jinkela_wire_1486),
        .dout(new_Jinkela_wire_1487)
    );

    bfr new_Jinkela_buffer_3797 (
        .din(new_Jinkela_wire_4419),
        .dout(new_Jinkela_wire_4420)
    );

    bfr new_Jinkela_buffer_3753 (
        .din(new_Jinkela_wire_4373),
        .dout(new_Jinkela_wire_4374)
    );

    bfr new_Jinkela_buffer_3013 (
        .din(new_Jinkela_wire_3440),
        .dout(new_Jinkela_wire_3441)
    );

    bfr new_Jinkela_buffer_1119 (
        .din(new_Jinkela_wire_1430),
        .dout(new_Jinkela_wire_1431)
    );

    bfr new_Jinkela_buffer_2897 (
        .din(new_Jinkela_wire_3320),
        .dout(new_Jinkela_wire_3321)
    );

    bfr new_Jinkela_buffer_1228 (
        .din(new_Jinkela_wire_1548),
        .dout(new_Jinkela_wire_1549)
    );

    bfr new_Jinkela_buffer_3811 (
        .din(new_Jinkela_wire_4444),
        .dout(new_Jinkela_wire_4445)
    );

    bfr new_Jinkela_buffer_3754 (
        .din(new_Jinkela_wire_4374),
        .dout(new_Jinkela_wire_4375)
    );

    bfr new_Jinkela_buffer_2949 (
        .din(new_Jinkela_wire_3376),
        .dout(new_Jinkela_wire_3377)
    );

    bfr new_Jinkela_buffer_1120 (
        .din(new_Jinkela_wire_1431),
        .dout(new_Jinkela_wire_1432)
    );

    bfr new_Jinkela_buffer_3809 (
        .din(new_Jinkela_wire_4442),
        .dout(new_Jinkela_wire_4443)
    );

    bfr new_Jinkela_buffer_2898 (
        .din(new_Jinkela_wire_3321),
        .dout(new_Jinkela_wire_3322)
    );

    bfr new_Jinkela_buffer_1171 (
        .din(new_Jinkela_wire_1487),
        .dout(new_Jinkela_wire_1488)
    );

    bfr new_Jinkela_buffer_3798 (
        .din(new_Jinkela_wire_4420),
        .dout(new_Jinkela_wire_4421)
    );

    bfr new_Jinkela_buffer_3755 (
        .din(new_Jinkela_wire_4375),
        .dout(new_Jinkela_wire_4376)
    );

    bfr new_Jinkela_buffer_3084 (
        .din(N222),
        .dout(new_Jinkela_wire_3514)
    );

    bfr new_Jinkela_buffer_1121 (
        .din(new_Jinkela_wire_1432),
        .dout(new_Jinkela_wire_1433)
    );

    bfr new_Jinkela_buffer_3016 (
        .din(new_Jinkela_wire_3443),
        .dout(new_Jinkela_wire_3444)
    );

    bfr new_Jinkela_buffer_2899 (
        .din(new_Jinkela_wire_3322),
        .dout(new_Jinkela_wire_3323)
    );

    bfr new_Jinkela_buffer_1292 (
        .din(new_Jinkela_wire_1612),
        .dout(new_Jinkela_wire_1613)
    );

    bfr new_Jinkela_buffer_3866 (
        .din(n_0430_),
        .dout(new_Jinkela_wire_4502)
    );

    bfr new_Jinkela_buffer_3756 (
        .din(new_Jinkela_wire_4376),
        .dout(new_Jinkela_wire_4377)
    );

    bfr new_Jinkela_buffer_2950 (
        .din(new_Jinkela_wire_3377),
        .dout(new_Jinkela_wire_3378)
    );

    bfr new_Jinkela_buffer_1122 (
        .din(new_Jinkela_wire_1433),
        .dout(new_Jinkela_wire_1434)
    );

    bfr new_Jinkela_buffer_2900 (
        .din(new_Jinkela_wire_3323),
        .dout(new_Jinkela_wire_3324)
    );

    bfr new_Jinkela_buffer_1172 (
        .din(new_Jinkela_wire_1488),
        .dout(new_Jinkela_wire_1489)
    );

    bfr new_Jinkela_buffer_3799 (
        .din(new_Jinkela_wire_4421),
        .dout(new_Jinkela_wire_4422)
    );

    bfr new_Jinkela_buffer_3757 (
        .din(new_Jinkela_wire_4377),
        .dout(new_Jinkela_wire_4378)
    );

    bfr new_Jinkela_buffer_3014 (
        .din(new_Jinkela_wire_3441),
        .dout(new_Jinkela_wire_3442)
    );

    bfr new_Jinkela_buffer_1123 (
        .din(new_Jinkela_wire_1434),
        .dout(new_Jinkela_wire_1435)
    );

    bfr new_Jinkela_buffer_2901 (
        .din(new_Jinkela_wire_3324),
        .dout(new_Jinkela_wire_3325)
    );

    bfr new_Jinkela_buffer_1229 (
        .din(new_Jinkela_wire_1549),
        .dout(new_Jinkela_wire_1550)
    );

    bfr new_Jinkela_buffer_3758 (
        .din(new_Jinkela_wire_4378),
        .dout(new_Jinkela_wire_4379)
    );

    bfr new_Jinkela_buffer_2951 (
        .din(new_Jinkela_wire_3378),
        .dout(new_Jinkela_wire_3379)
    );

    bfr new_Jinkela_buffer_1124 (
        .din(new_Jinkela_wire_1435),
        .dout(new_Jinkela_wire_1436)
    );

    bfr new_Jinkela_buffer_2902 (
        .din(new_Jinkela_wire_3325),
        .dout(new_Jinkela_wire_3326)
    );

    bfr new_Jinkela_buffer_1173 (
        .din(new_Jinkela_wire_1489),
        .dout(new_Jinkela_wire_1490)
    );

    bfr new_Jinkela_buffer_3800 (
        .din(new_Jinkela_wire_4422),
        .dout(new_Jinkela_wire_4423)
    );

    bfr new_Jinkela_buffer_3759 (
        .din(new_Jinkela_wire_4379),
        .dout(new_Jinkela_wire_4380)
    );

    bfr new_Jinkela_buffer_1125 (
        .din(new_Jinkela_wire_1436),
        .dout(new_Jinkela_wire_1437)
    );

    spl2 new_Jinkela_splitter_230 (
        .a(n_1108_),
        .b(new_Jinkela_wire_4503),
        .c(new_Jinkela_wire_4504)
    );

    bfr new_Jinkela_buffer_2903 (
        .din(new_Jinkela_wire_3326),
        .dout(new_Jinkela_wire_3327)
    );

    bfr new_Jinkela_buffer_3760 (
        .din(new_Jinkela_wire_4380),
        .dout(new_Jinkela_wire_4381)
    );

    bfr new_Jinkela_buffer_2952 (
        .din(new_Jinkela_wire_3379),
        .dout(new_Jinkela_wire_3380)
    );

    bfr new_Jinkela_buffer_1126 (
        .din(new_Jinkela_wire_1437),
        .dout(new_Jinkela_wire_1438)
    );

    bfr new_Jinkela_buffer_2904 (
        .din(new_Jinkela_wire_3327),
        .dout(new_Jinkela_wire_3328)
    );

    bfr new_Jinkela_buffer_1174 (
        .din(new_Jinkela_wire_1490),
        .dout(new_Jinkela_wire_1491)
    );

    bfr new_Jinkela_buffer_3801 (
        .din(new_Jinkela_wire_4423),
        .dout(new_Jinkela_wire_4424)
    );

    bfr new_Jinkela_buffer_3761 (
        .din(new_Jinkela_wire_4381),
        .dout(new_Jinkela_wire_4382)
    );

    bfr new_Jinkela_buffer_3081 (
        .din(new_Jinkela_wire_3510),
        .dout(new_Jinkela_wire_3511)
    );

    bfr new_Jinkela_buffer_1127 (
        .din(new_Jinkela_wire_1438),
        .dout(new_Jinkela_wire_1439)
    );

    bfr new_Jinkela_buffer_3017 (
        .din(new_Jinkela_wire_3444),
        .dout(new_Jinkela_wire_3445)
    );

    bfr new_Jinkela_buffer_1230 (
        .din(new_Jinkela_wire_1550),
        .dout(new_Jinkela_wire_1551)
    );

    bfr new_Jinkela_buffer_2905 (
        .din(new_Jinkela_wire_3328),
        .dout(new_Jinkela_wire_3329)
    );

    bfr new_Jinkela_buffer_3812 (
        .din(new_Jinkela_wire_4445),
        .dout(new_Jinkela_wire_4446)
    );

    bfr new_Jinkela_buffer_3762 (
        .din(new_Jinkela_wire_4382),
        .dout(new_Jinkela_wire_4383)
    );

    bfr new_Jinkela_buffer_1128 (
        .din(new_Jinkela_wire_1439),
        .dout(new_Jinkela_wire_1440)
    );

    bfr new_Jinkela_buffer_2953 (
        .din(new_Jinkela_wire_3380),
        .dout(new_Jinkela_wire_3381)
    );

    bfr new_Jinkela_buffer_1175 (
        .din(new_Jinkela_wire_1491),
        .dout(new_Jinkela_wire_1492)
    );

    bfr new_Jinkela_buffer_2906 (
        .din(new_Jinkela_wire_3329),
        .dout(new_Jinkela_wire_3330)
    );

    bfr new_Jinkela_buffer_3802 (
        .din(new_Jinkela_wire_4424),
        .dout(new_Jinkela_wire_4425)
    );

    bfr new_Jinkela_buffer_3763 (
        .din(new_Jinkela_wire_4383),
        .dout(new_Jinkela_wire_4384)
    );

    bfr new_Jinkela_buffer_1129 (
        .din(new_Jinkela_wire_1440),
        .dout(new_Jinkela_wire_1441)
    );

    bfr new_Jinkela_buffer_1295 (
        .din(new_Jinkela_wire_1615),
        .dout(new_Jinkela_wire_1616)
    );

    bfr new_Jinkela_buffer_2907 (
        .din(new_Jinkela_wire_3330),
        .dout(new_Jinkela_wire_3331)
    );

    spl2 new_Jinkela_splitter_229 (
        .a(new_Jinkela_wire_4486),
        .b(new_Jinkela_wire_4487),
        .c(new_Jinkela_wire_4488)
    );

    bfr new_Jinkela_buffer_1358 (
        .din(new_Jinkela_wire_1683),
        .dout(new_Jinkela_wire_1684)
    );

    bfr new_Jinkela_buffer_3764 (
        .din(new_Jinkela_wire_4384),
        .dout(new_Jinkela_wire_4385)
    );

    bfr new_Jinkela_buffer_1130 (
        .din(new_Jinkela_wire_1441),
        .dout(new_Jinkela_wire_1442)
    );

    bfr new_Jinkela_buffer_2954 (
        .din(new_Jinkela_wire_3381),
        .dout(new_Jinkela_wire_3382)
    );

    bfr new_Jinkela_buffer_1176 (
        .din(new_Jinkela_wire_1492),
        .dout(new_Jinkela_wire_1493)
    );

    bfr new_Jinkela_buffer_2908 (
        .din(new_Jinkela_wire_3331),
        .dout(new_Jinkela_wire_3332)
    );

    bfr new_Jinkela_buffer_3803 (
        .din(new_Jinkela_wire_4425),
        .dout(new_Jinkela_wire_4426)
    );

    bfr new_Jinkela_buffer_3765 (
        .din(new_Jinkela_wire_4385),
        .dout(new_Jinkela_wire_4386)
    );

    bfr new_Jinkela_buffer_1131 (
        .din(new_Jinkela_wire_1442),
        .dout(new_Jinkela_wire_1443)
    );

    spl4L new_Jinkela_splitter_147 (
        .a(N382),
        .d(new_Jinkela_wire_3518),
        .b(new_Jinkela_wire_3519),
        .e(new_Jinkela_wire_3520),
        .c(new_Jinkela_wire_3521)
    );

    spl2 new_Jinkela_splitter_146 (
        .a(new_Jinkela_wire_3445),
        .b(new_Jinkela_wire_3446),
        .c(new_Jinkela_wire_3447)
    );

    bfr new_Jinkela_buffer_1231 (
        .din(new_Jinkela_wire_1551),
        .dout(new_Jinkela_wire_1552)
    );

    bfr new_Jinkela_buffer_2909 (
        .din(new_Jinkela_wire_3332),
        .dout(new_Jinkela_wire_3333)
    );

    bfr new_Jinkela_buffer_3813 (
        .din(new_Jinkela_wire_4446),
        .dout(new_Jinkela_wire_4447)
    );

    bfr new_Jinkela_buffer_3766 (
        .din(new_Jinkela_wire_4386),
        .dout(new_Jinkela_wire_4387)
    );

    bfr new_Jinkela_buffer_1132 (
        .din(new_Jinkela_wire_1443),
        .dout(new_Jinkela_wire_1444)
    );

    bfr new_Jinkela_buffer_2955 (
        .din(new_Jinkela_wire_3382),
        .dout(new_Jinkela_wire_3383)
    );

    bfr new_Jinkela_buffer_1177 (
        .din(new_Jinkela_wire_1493),
        .dout(new_Jinkela_wire_1494)
    );

    bfr new_Jinkela_buffer_2910 (
        .din(new_Jinkela_wire_3333),
        .dout(new_Jinkela_wire_3334)
    );

    bfr new_Jinkela_buffer_3804 (
        .din(new_Jinkela_wire_4426),
        .dout(new_Jinkela_wire_4427)
    );

    bfr new_Jinkela_buffer_3767 (
        .din(new_Jinkela_wire_4387),
        .dout(new_Jinkela_wire_4388)
    );

    bfr new_Jinkela_buffer_1133 (
        .din(new_Jinkela_wire_1444),
        .dout(new_Jinkela_wire_1445)
    );

    bfr new_Jinkela_buffer_3018 (
        .din(new_Jinkela_wire_3447),
        .dout(new_Jinkela_wire_3448)
    );

    bfr new_Jinkela_buffer_1294 (
        .din(new_Jinkela_wire_1614),
        .dout(new_Jinkela_wire_1615)
    );

    bfr new_Jinkela_buffer_2911 (
        .din(new_Jinkela_wire_3334),
        .dout(new_Jinkela_wire_3335)
    );

    bfr new_Jinkela_buffer_3768 (
        .din(new_Jinkela_wire_4388),
        .dout(new_Jinkela_wire_4389)
    );

    bfr new_Jinkela_buffer_1134 (
        .din(new_Jinkela_wire_1445),
        .dout(new_Jinkela_wire_1446)
    );

    bfr new_Jinkela_buffer_2956 (
        .din(new_Jinkela_wire_3383),
        .dout(new_Jinkela_wire_3384)
    );

    bfr new_Jinkela_buffer_3853 (
        .din(new_Jinkela_wire_4488),
        .dout(new_Jinkela_wire_4489)
    );

    bfr new_Jinkela_buffer_1178 (
        .din(new_Jinkela_wire_1494),
        .dout(new_Jinkela_wire_1495)
    );

    bfr new_Jinkela_buffer_2912 (
        .din(new_Jinkela_wire_3335),
        .dout(new_Jinkela_wire_3336)
    );

    bfr new_Jinkela_buffer_3814 (
        .din(new_Jinkela_wire_4447),
        .dout(new_Jinkela_wire_4448)
    );

    bfr new_Jinkela_buffer_3769 (
        .din(new_Jinkela_wire_4389),
        .dout(new_Jinkela_wire_4390)
    );

    bfr new_Jinkela_buffer_1135 (
        .din(new_Jinkela_wire_1446),
        .dout(new_Jinkela_wire_1447)
    );

    bfr new_Jinkela_buffer_3090 (
        .din(N238),
        .dout(new_Jinkela_wire_3524)
    );

    bfr new_Jinkela_buffer_1232 (
        .din(new_Jinkela_wire_1552),
        .dout(new_Jinkela_wire_1553)
    );

    bfr new_Jinkela_buffer_2913 (
        .din(new_Jinkela_wire_3336),
        .dout(new_Jinkela_wire_3337)
    );

    bfr new_Jinkela_buffer_3770 (
        .din(new_Jinkela_wire_4390),
        .dout(new_Jinkela_wire_4391)
    );

    bfr new_Jinkela_buffer_1136 (
        .din(new_Jinkela_wire_1447),
        .dout(new_Jinkela_wire_1448)
    );

    bfr new_Jinkela_buffer_2957 (
        .din(new_Jinkela_wire_3384),
        .dout(new_Jinkela_wire_3385)
    );

    bfr new_Jinkela_buffer_3867 (
        .din(n_0734_),
        .dout(new_Jinkela_wire_4505)
    );

    bfr new_Jinkela_buffer_1179 (
        .din(new_Jinkela_wire_1495),
        .dout(new_Jinkela_wire_1496)
    );

    bfr new_Jinkela_buffer_2914 (
        .din(new_Jinkela_wire_3337),
        .dout(new_Jinkela_wire_3338)
    );

    bfr new_Jinkela_buffer_3815 (
        .din(new_Jinkela_wire_4448),
        .dout(new_Jinkela_wire_4449)
    );

    spl2 new_Jinkela_splitter_224 (
        .a(new_Jinkela_wire_4391),
        .b(new_Jinkela_wire_4392),
        .c(new_Jinkela_wire_4393)
    );

    bfr new_Jinkela_buffer_7592 (
        .din(new_Jinkela_wire_9513),
        .dout(new_Jinkela_wire_9514)
    );

    spl2 new_Jinkela_splitter_775 (
        .a(n_0436_),
        .b(new_Jinkela_wire_9551),
        .c(new_Jinkela_wire_9552)
    );

    bfr new_Jinkela_buffer_7593 (
        .din(new_Jinkela_wire_9514),
        .dout(new_Jinkela_wire_9515)
    );

    bfr new_Jinkela_buffer_7605 (
        .din(new_Jinkela_wire_9526),
        .dout(new_Jinkela_wire_9527)
    );

    bfr new_Jinkela_buffer_7594 (
        .din(new_Jinkela_wire_9515),
        .dout(new_Jinkela_wire_9516)
    );

    bfr new_Jinkela_buffer_7595 (
        .din(new_Jinkela_wire_9516),
        .dout(new_Jinkela_wire_9517)
    );

    bfr new_Jinkela_buffer_7606 (
        .din(new_Jinkela_wire_9527),
        .dout(new_Jinkela_wire_9528)
    );

    bfr new_Jinkela_buffer_7596 (
        .din(new_Jinkela_wire_9517),
        .dout(new_Jinkela_wire_9518)
    );

    spl2 new_Jinkela_splitter_774 (
        .a(n_0756_),
        .b(new_Jinkela_wire_9549),
        .c(new_Jinkela_wire_9550)
    );

    bfr new_Jinkela_buffer_7607 (
        .din(new_Jinkela_wire_9528),
        .dout(new_Jinkela_wire_9529)
    );

    spl2 new_Jinkela_splitter_773 (
        .a(new_Jinkela_wire_9545),
        .b(new_Jinkela_wire_9546),
        .c(new_Jinkela_wire_9547)
    );

    bfr new_Jinkela_buffer_7615 (
        .din(n_0749_),
        .dout(new_Jinkela_wire_9553)
    );

    bfr new_Jinkela_buffer_7608 (
        .din(new_Jinkela_wire_9529),
        .dout(new_Jinkela_wire_9530)
    );

    bfr new_Jinkela_buffer_7609 (
        .din(new_Jinkela_wire_9530),
        .dout(new_Jinkela_wire_9531)
    );

    spl2 new_Jinkela_splitter_777 (
        .a(n_1337_),
        .b(new_Jinkela_wire_9556),
        .c(new_Jinkela_wire_9557)
    );

    bfr new_Jinkela_buffer_7610 (
        .din(new_Jinkela_wire_9531),
        .dout(new_Jinkela_wire_9532)
    );

    spl2 new_Jinkela_splitter_776 (
        .a(n_0744_),
        .b(new_Jinkela_wire_9554),
        .c(new_Jinkela_wire_9555)
    );

    spl2 new_Jinkela_splitter_778 (
        .a(n_0706_),
        .b(new_Jinkela_wire_9570),
        .c(new_Jinkela_wire_9571)
    );

    bfr new_Jinkela_buffer_7616 (
        .din(new_Jinkela_wire_9557),
        .dout(new_Jinkela_wire_9558)
    );

    spl2 new_Jinkela_splitter_779 (
        .a(n_0070_),
        .b(new_Jinkela_wire_9572),
        .c(new_Jinkela_wire_9576)
    );

    bfr new_Jinkela_buffer_7635 (
        .din(n_0278_),
        .dout(new_Jinkela_wire_9598)
    );

    bfr new_Jinkela_buffer_7617 (
        .din(new_Jinkela_wire_9558),
        .dout(new_Jinkela_wire_9559)
    );

    bfr new_Jinkela_buffer_7618 (
        .din(new_Jinkela_wire_9559),
        .dout(new_Jinkela_wire_9560)
    );

    spl3L new_Jinkela_splitter_782 (
        .a(n_0024_),
        .d(new_Jinkela_wire_9582),
        .b(new_Jinkela_wire_9583),
        .c(new_Jinkela_wire_9584)
    );

    spl2 new_Jinkela_splitter_786 (
        .a(n_0485_),
        .b(new_Jinkela_wire_9599),
        .c(new_Jinkela_wire_9600)
    );

    bfr new_Jinkela_buffer_7619 (
        .din(new_Jinkela_wire_9560),
        .dout(new_Jinkela_wire_9561)
    );

    bfr new_Jinkela_buffer_7628 (
        .din(n_0141_),
        .dout(new_Jinkela_wire_9581)
    );

    spl4L new_Jinkela_splitter_781 (
        .a(new_Jinkela_wire_9576),
        .d(new_Jinkela_wire_9577),
        .b(new_Jinkela_wire_9578),
        .e(new_Jinkela_wire_9579),
        .c(new_Jinkela_wire_9580)
    );

    bfr new_Jinkela_buffer_7620 (
        .din(new_Jinkela_wire_9561),
        .dout(new_Jinkela_wire_9562)
    );

    spl3L new_Jinkela_splitter_783 (
        .a(n_0707_),
        .d(new_Jinkela_wire_9585),
        .b(new_Jinkela_wire_9586),
        .c(new_Jinkela_wire_9587)
    );

    bfr new_Jinkela_buffer_7621 (
        .din(new_Jinkela_wire_9562),
        .dout(new_Jinkela_wire_9563)
    );

    spl3L new_Jinkela_splitter_780 (
        .a(new_Jinkela_wire_9572),
        .d(new_Jinkela_wire_9573),
        .b(new_Jinkela_wire_9574),
        .c(new_Jinkela_wire_9575)
    );

    bfr new_Jinkela_buffer_7622 (
        .din(new_Jinkela_wire_9563),
        .dout(new_Jinkela_wire_9564)
    );

    spl3L new_Jinkela_splitter_787 (
        .a(n_1127_),
        .d(new_Jinkela_wire_9601),
        .b(new_Jinkela_wire_9602),
        .c(new_Jinkela_wire_9603)
    );

    spl2 new_Jinkela_splitter_788 (
        .a(n_0500_),
        .b(new_Jinkela_wire_9604),
        .c(new_Jinkela_wire_9605)
    );

    bfr new_Jinkela_buffer_7623 (
        .din(new_Jinkela_wire_9564),
        .dout(new_Jinkela_wire_9565)
    );

    bfr new_Jinkela_buffer_7629 (
        .din(new_Jinkela_wire_9587),
        .dout(new_Jinkela_wire_9588)
    );

    bfr new_Jinkela_buffer_7624 (
        .din(new_Jinkela_wire_9565),
        .dout(new_Jinkela_wire_9566)
    );

    bfr new_Jinkela_buffer_7625 (
        .din(new_Jinkela_wire_9566),
        .dout(new_Jinkela_wire_9567)
    );

    bfr new_Jinkela_buffer_7626 (
        .din(new_Jinkela_wire_9567),
        .dout(new_Jinkela_wire_9568)
    );

    bfr new_Jinkela_buffer_7630 (
        .din(new_Jinkela_wire_9588),
        .dout(new_Jinkela_wire_9589)
    );

    bfr new_Jinkela_buffer_7099 (
        .din(new_Jinkela_wire_8782),
        .dout(new_Jinkela_wire_8783)
    );

    bfr new_Jinkela_buffer_8297 (
        .din(new_Jinkela_wire_10434),
        .dout(new_Jinkela_wire_10435)
    );

    bfr new_Jinkela_buffer_4611 (
        .din(new_Jinkela_wire_5489),
        .dout(new_Jinkela_wire_5490)
    );

    bfr new_Jinkela_buffer_8273 (
        .din(new_Jinkela_wire_10396),
        .dout(new_Jinkela_wire_10397)
    );

    bfr new_Jinkela_buffer_7150 (
        .din(new_Jinkela_wire_8851),
        .dout(new_Jinkela_wire_8852)
    );

    bfr new_Jinkela_buffer_7100 (
        .din(new_Jinkela_wire_8783),
        .dout(new_Jinkela_wire_8784)
    );

    bfr new_Jinkela_buffer_8292 (
        .din(new_Jinkela_wire_10425),
        .dout(new_Jinkela_wire_10426)
    );

    bfr new_Jinkela_buffer_4638 (
        .din(new_Jinkela_wire_5518),
        .dout(new_Jinkela_wire_5519)
    );

    bfr new_Jinkela_buffer_4612 (
        .din(new_Jinkela_wire_5490),
        .dout(new_Jinkela_wire_5491)
    );

    bfr new_Jinkela_buffer_7134 (
        .din(new_Jinkela_wire_8828),
        .dout(new_Jinkela_wire_8829)
    );

    bfr new_Jinkela_buffer_8274 (
        .din(new_Jinkela_wire_10397),
        .dout(new_Jinkela_wire_10398)
    );

    bfr new_Jinkela_buffer_7101 (
        .din(new_Jinkela_wire_8784),
        .dout(new_Jinkela_wire_8785)
    );

    bfr new_Jinkela_buffer_8308 (
        .din(new_net_2493),
        .dout(new_Jinkela_wire_10448)
    );

    bfr new_Jinkela_buffer_4613 (
        .din(new_Jinkela_wire_5491),
        .dout(new_Jinkela_wire_5492)
    );

    bfr new_Jinkela_buffer_7149 (
        .din(new_Jinkela_wire_8848),
        .dout(new_Jinkela_wire_8849)
    );

    bfr new_Jinkela_buffer_8275 (
        .din(new_Jinkela_wire_10398),
        .dout(new_Jinkela_wire_10399)
    );

    spl2 new_Jinkela_splitter_340 (
        .a(n_1329_),
        .b(new_Jinkela_wire_5577),
        .c(new_Jinkela_wire_5578)
    );

    bfr new_Jinkela_buffer_7102 (
        .din(new_Jinkela_wire_8785),
        .dout(new_Jinkela_wire_8786)
    );

    bfr new_Jinkela_buffer_8293 (
        .din(new_Jinkela_wire_10426),
        .dout(new_Jinkela_wire_10427)
    );

    bfr new_Jinkela_buffer_4639 (
        .din(new_Jinkela_wire_5519),
        .dout(new_Jinkela_wire_5520)
    );

    bfr new_Jinkela_buffer_4614 (
        .din(new_Jinkela_wire_5492),
        .dout(new_Jinkela_wire_5493)
    );

    bfr new_Jinkela_buffer_7135 (
        .din(new_Jinkela_wire_8829),
        .dout(new_Jinkela_wire_8830)
    );

    bfr new_Jinkela_buffer_8276 (
        .din(new_Jinkela_wire_10399),
        .dout(new_Jinkela_wire_10400)
    );

    bfr new_Jinkela_buffer_7103 (
        .din(new_Jinkela_wire_8786),
        .dout(new_Jinkela_wire_8787)
    );

    bfr new_Jinkela_buffer_4615 (
        .din(new_Jinkela_wire_5493),
        .dout(new_Jinkela_wire_5494)
    );

    bfr new_Jinkela_buffer_8277 (
        .din(new_Jinkela_wire_10400),
        .dout(new_Jinkela_wire_10401)
    );

    bfr new_Jinkela_buffer_7104 (
        .din(new_Jinkela_wire_8787),
        .dout(new_Jinkela_wire_8788)
    );

    spl2 new_Jinkela_splitter_857 (
        .a(new_Jinkela_wire_10427),
        .b(new_Jinkela_wire_10428),
        .c(new_Jinkela_wire_10429)
    );

    bfr new_Jinkela_buffer_4640 (
        .din(new_Jinkela_wire_5520),
        .dout(new_Jinkela_wire_5521)
    );

    bfr new_Jinkela_buffer_4616 (
        .din(new_Jinkela_wire_5494),
        .dout(new_Jinkela_wire_5495)
    );

    bfr new_Jinkela_buffer_7136 (
        .din(new_Jinkela_wire_8830),
        .dout(new_Jinkela_wire_8831)
    );

    bfr new_Jinkela_buffer_8278 (
        .din(new_Jinkela_wire_10401),
        .dout(new_Jinkela_wire_10402)
    );

    bfr new_Jinkela_buffer_7105 (
        .din(new_Jinkela_wire_8788),
        .dout(new_Jinkela_wire_8789)
    );

    bfr new_Jinkela_buffer_8294 (
        .din(new_Jinkela_wire_10429),
        .dout(new_Jinkela_wire_10430)
    );

    spl2 new_Jinkela_splitter_341 (
        .a(n_0795_),
        .b(new_Jinkela_wire_5588),
        .c(new_Jinkela_wire_5589)
    );

    bfr new_Jinkela_buffer_4617 (
        .din(new_Jinkela_wire_5495),
        .dout(new_Jinkela_wire_5496)
    );

    spl2 new_Jinkela_splitter_681 (
        .a(n_1129_),
        .b(new_Jinkela_wire_8868),
        .c(new_Jinkela_wire_8869)
    );

    bfr new_Jinkela_buffer_8279 (
        .din(new_Jinkela_wire_10402),
        .dout(new_Jinkela_wire_10403)
    );

    spl2 new_Jinkela_splitter_682 (
        .a(n_1305_),
        .b(new_Jinkela_wire_8870),
        .c(new_Jinkela_wire_8871)
    );

    bfr new_Jinkela_buffer_4680 (
        .din(new_Jinkela_wire_5578),
        .dout(new_Jinkela_wire_5579)
    );

    bfr new_Jinkela_buffer_7106 (
        .din(new_Jinkela_wire_8789),
        .dout(new_Jinkela_wire_8790)
    );

    bfr new_Jinkela_buffer_8345 (
        .din(n_0286_),
        .dout(new_Jinkela_wire_10485)
    );

    bfr new_Jinkela_buffer_4641 (
        .din(new_Jinkela_wire_5521),
        .dout(new_Jinkela_wire_5522)
    );

    bfr new_Jinkela_buffer_8298 (
        .din(new_Jinkela_wire_10435),
        .dout(new_Jinkela_wire_10436)
    );

    bfr new_Jinkela_buffer_4618 (
        .din(new_Jinkela_wire_5496),
        .dout(new_Jinkela_wire_5497)
    );

    bfr new_Jinkela_buffer_7137 (
        .din(new_Jinkela_wire_8831),
        .dout(new_Jinkela_wire_8832)
    );

    bfr new_Jinkela_buffer_8280 (
        .din(new_Jinkela_wire_10403),
        .dout(new_Jinkela_wire_10404)
    );

    bfr new_Jinkela_buffer_7107 (
        .din(new_Jinkela_wire_8790),
        .dout(new_Jinkela_wire_8791)
    );

    bfr new_Jinkela_buffer_4689 (
        .din(new_net_2554),
        .dout(new_Jinkela_wire_5590)
    );

    bfr new_Jinkela_buffer_8306 (
        .din(new_Jinkela_wire_10443),
        .dout(new_Jinkela_wire_10444)
    );

    bfr new_Jinkela_buffer_4619 (
        .din(new_Jinkela_wire_5497),
        .dout(new_Jinkela_wire_5498)
    );

    bfr new_Jinkela_buffer_7152 (
        .din(new_Jinkela_wire_8853),
        .dout(new_Jinkela_wire_8854)
    );

    bfr new_Jinkela_buffer_8281 (
        .din(new_Jinkela_wire_10404),
        .dout(new_Jinkela_wire_10405)
    );

    spl2 new_Jinkela_splitter_346 (
        .a(n_0274_),
        .b(new_Jinkela_wire_5637),
        .c(new_Jinkela_wire_5638)
    );

    bfr new_Jinkela_buffer_7108 (
        .din(new_Jinkela_wire_8791),
        .dout(new_Jinkela_wire_8792)
    );

    bfr new_Jinkela_buffer_8295 (
        .din(new_Jinkela_wire_10430),
        .dout(new_Jinkela_wire_10431)
    );

    bfr new_Jinkela_buffer_4642 (
        .din(new_Jinkela_wire_5522),
        .dout(new_Jinkela_wire_5523)
    );

    bfr new_Jinkela_buffer_4620 (
        .din(new_Jinkela_wire_5498),
        .dout(new_Jinkela_wire_5499)
    );

    bfr new_Jinkela_buffer_7138 (
        .din(new_Jinkela_wire_8832),
        .dout(new_Jinkela_wire_8833)
    );

    bfr new_Jinkela_buffer_8282 (
        .din(new_Jinkela_wire_10405),
        .dout(new_Jinkela_wire_10406)
    );

    bfr new_Jinkela_buffer_7109 (
        .din(new_Jinkela_wire_8792),
        .dout(new_Jinkela_wire_8793)
    );

    bfr new_Jinkela_buffer_8299 (
        .din(new_Jinkela_wire_10436),
        .dout(new_Jinkela_wire_10437)
    );

    bfr new_Jinkela_buffer_4681 (
        .din(new_Jinkela_wire_5579),
        .dout(new_Jinkela_wire_5580)
    );

    bfr new_Jinkela_buffer_8283 (
        .din(new_Jinkela_wire_10406),
        .dout(new_Jinkela_wire_10407)
    );

    bfr new_Jinkela_buffer_4643 (
        .din(new_Jinkela_wire_5523),
        .dout(new_Jinkela_wire_5524)
    );

    bfr new_Jinkela_buffer_7110 (
        .din(new_Jinkela_wire_8793),
        .dout(new_Jinkela_wire_8794)
    );

    spl3L new_Jinkela_splitter_343 (
        .a(n_0367_),
        .d(new_Jinkela_wire_5593),
        .b(new_Jinkela_wire_5594),
        .c(new_Jinkela_wire_5595)
    );

    bfr new_Jinkela_buffer_7139 (
        .din(new_Jinkela_wire_8833),
        .dout(new_Jinkela_wire_8834)
    );

    bfr new_Jinkela_buffer_8284 (
        .din(new_Jinkela_wire_10407),
        .dout(new_Jinkela_wire_10408)
    );

    bfr new_Jinkela_buffer_4644 (
        .din(new_Jinkela_wire_5524),
        .dout(new_Jinkela_wire_5525)
    );

    bfr new_Jinkela_buffer_7111 (
        .din(new_Jinkela_wire_8794),
        .dout(new_Jinkela_wire_8795)
    );

    bfr new_Jinkela_buffer_8309 (
        .din(new_Jinkela_wire_10448),
        .dout(new_Jinkela_wire_10449)
    );

    spl2 new_Jinkela_splitter_342 (
        .a(n_0131_),
        .b(new_Jinkela_wire_5591),
        .c(new_Jinkela_wire_5592)
    );

    bfr new_Jinkela_buffer_8300 (
        .din(new_Jinkela_wire_10437),
        .dout(new_Jinkela_wire_10438)
    );

    bfr new_Jinkela_buffer_4682 (
        .din(new_Jinkela_wire_5580),
        .dout(new_Jinkela_wire_5581)
    );

    bfr new_Jinkela_buffer_7153 (
        .din(new_Jinkela_wire_8854),
        .dout(new_Jinkela_wire_8855)
    );

    bfr new_Jinkela_buffer_8285 (
        .din(new_Jinkela_wire_10408),
        .dout(new_Jinkela_wire_10409)
    );

    bfr new_Jinkela_buffer_4645 (
        .din(new_Jinkela_wire_5525),
        .dout(new_Jinkela_wire_5526)
    );

    bfr new_Jinkela_buffer_7112 (
        .din(new_Jinkela_wire_8795),
        .dout(new_Jinkela_wire_8796)
    );

    bfr new_Jinkela_buffer_8307 (
        .din(new_Jinkela_wire_10444),
        .dout(new_Jinkela_wire_10445)
    );

    bfr new_Jinkela_buffer_7140 (
        .din(new_Jinkela_wire_8834),
        .dout(new_Jinkela_wire_8835)
    );

    bfr new_Jinkela_buffer_8286 (
        .din(new_Jinkela_wire_10409),
        .dout(new_Jinkela_wire_10410)
    );

    bfr new_Jinkela_buffer_4646 (
        .din(new_Jinkela_wire_5526),
        .dout(new_Jinkela_wire_5527)
    );

    bfr new_Jinkela_buffer_7113 (
        .din(new_Jinkela_wire_8796),
        .dout(new_Jinkela_wire_8797)
    );

    bfr new_Jinkela_buffer_8301 (
        .din(new_Jinkela_wire_10438),
        .dout(new_Jinkela_wire_10439)
    );

    bfr new_Jinkela_buffer_4683 (
        .din(new_Jinkela_wire_5581),
        .dout(new_Jinkela_wire_5582)
    );

    bfr new_Jinkela_buffer_8287 (
        .din(new_Jinkela_wire_10410),
        .dout(new_Jinkela_wire_10411)
    );

    bfr new_Jinkela_buffer_4647 (
        .din(new_Jinkela_wire_5527),
        .dout(new_Jinkela_wire_5528)
    );

    bfr new_Jinkela_buffer_7168 (
        .din(n_1232_),
        .dout(new_Jinkela_wire_8874)
    );

    bfr new_Jinkela_buffer_7114 (
        .din(new_Jinkela_wire_8797),
        .dout(new_Jinkela_wire_8798)
    );

    spl2 new_Jinkela_splitter_345 (
        .a(n_0073_),
        .b(new_Jinkela_wire_5635),
        .c(new_Jinkela_wire_5636)
    );

    bfr new_Jinkela_buffer_7141 (
        .din(new_Jinkela_wire_8835),
        .dout(new_Jinkela_wire_8836)
    );

    bfr new_Jinkela_buffer_8288 (
        .din(new_Jinkela_wire_10411),
        .dout(new_Jinkela_wire_10412)
    );

    bfr new_Jinkela_buffer_4648 (
        .din(new_Jinkela_wire_5528),
        .dout(new_Jinkela_wire_5529)
    );

    bfr new_Jinkela_buffer_7115 (
        .din(new_Jinkela_wire_8798),
        .dout(new_Jinkela_wire_8799)
    );

    bfr new_Jinkela_buffer_8346 (
        .din(new_net_2505),
        .dout(new_Jinkela_wire_10486)
    );

    bfr new_Jinkela_buffer_8302 (
        .din(new_Jinkela_wire_10439),
        .dout(new_Jinkela_wire_10440)
    );

    bfr new_Jinkela_buffer_4684 (
        .din(new_Jinkela_wire_5582),
        .dout(new_Jinkela_wire_5583)
    );

    bfr new_Jinkela_buffer_7154 (
        .din(new_Jinkela_wire_8855),
        .dout(new_Jinkela_wire_8856)
    );

    bfr new_Jinkela_buffer_8289 (
        .din(new_Jinkela_wire_10412),
        .dout(new_Jinkela_wire_10413)
    );

    bfr new_Jinkela_buffer_4649 (
        .din(new_Jinkela_wire_5529),
        .dout(new_Jinkela_wire_5530)
    );

    bfr new_Jinkela_buffer_7116 (
        .din(new_Jinkela_wire_8799),
        .dout(new_Jinkela_wire_8800)
    );

    spl2 new_Jinkela_splitter_859 (
        .a(new_Jinkela_wire_10445),
        .b(new_Jinkela_wire_10446),
        .c(new_Jinkela_wire_10447)
    );

    spl4L new_Jinkela_splitter_347 (
        .a(n_1253_),
        .d(new_Jinkela_wire_5639),
        .b(new_Jinkela_wire_5640),
        .e(new_Jinkela_wire_5641),
        .c(new_Jinkela_wire_5642)
    );

    bfr new_Jinkela_buffer_7142 (
        .din(new_Jinkela_wire_8836),
        .dout(new_Jinkela_wire_8837)
    );

    bfr new_Jinkela_buffer_8290 (
        .din(new_Jinkela_wire_10413),
        .dout(new_Jinkela_wire_10414)
    );

    bfr new_Jinkela_buffer_4650 (
        .din(new_Jinkela_wire_5530),
        .dout(new_Jinkela_wire_5531)
    );

    bfr new_Jinkela_buffer_7117 (
        .din(new_Jinkela_wire_8800),
        .dout(new_Jinkela_wire_8801)
    );

    bfr new_Jinkela_buffer_4690 (
        .din(new_Jinkela_wire_5595),
        .dout(new_Jinkela_wire_5596)
    );

    bfr new_Jinkela_buffer_8303 (
        .din(new_Jinkela_wire_10440),
        .dout(new_Jinkela_wire_10441)
    );

    bfr new_Jinkela_buffer_4685 (
        .din(new_Jinkela_wire_5583),
        .dout(new_Jinkela_wire_5584)
    );

    bfr new_Jinkela_buffer_7166 (
        .din(new_Jinkela_wire_8871),
        .dout(new_Jinkela_wire_8872)
    );

    spl2 new_Jinkela_splitter_853 (
        .a(new_Jinkela_wire_10414),
        .b(new_Jinkela_wire_10415),
        .c(new_Jinkela_wire_10416)
    );

    bfr new_Jinkela_buffer_4651 (
        .din(new_Jinkela_wire_5531),
        .dout(new_Jinkela_wire_5532)
    );

    bfr new_Jinkela_buffer_7118 (
        .din(new_Jinkela_wire_8801),
        .dout(new_Jinkela_wire_8802)
    );

    spl2 new_Jinkela_splitter_860 (
        .a(n_1368_),
        .b(new_Jinkela_wire_10502),
        .c(new_Jinkela_wire_10503)
    );

    bfr new_Jinkela_buffer_8304 (
        .din(new_Jinkela_wire_10441),
        .dout(new_Jinkela_wire_10442)
    );

    bfr new_Jinkela_buffer_7143 (
        .din(new_Jinkela_wire_8837),
        .dout(new_Jinkela_wire_8838)
    );

    bfr new_Jinkela_buffer_4652 (
        .din(new_Jinkela_wire_5532),
        .dout(new_Jinkela_wire_5533)
    );

    bfr new_Jinkela_buffer_7119 (
        .din(new_Jinkela_wire_8802),
        .dout(new_Jinkela_wire_8803)
    );

    bfr new_Jinkela_buffer_4686 (
        .din(new_Jinkela_wire_5584),
        .dout(new_Jinkela_wire_5585)
    );

    bfr new_Jinkela_buffer_7155 (
        .din(new_Jinkela_wire_8856),
        .dout(new_Jinkela_wire_8857)
    );

    bfr new_Jinkela_buffer_8310 (
        .din(new_Jinkela_wire_10449),
        .dout(new_Jinkela_wire_10450)
    );

    spl2 new_Jinkela_splitter_767 (
        .a(new_Jinkela_wire_9482),
        .b(new_Jinkela_wire_9483),
        .c(new_Jinkela_wire_9484)
    );

    spl2 new_Jinkela_splitter_430 (
        .a(n_1298_),
        .b(new_Jinkela_wire_6674),
        .c(new_Jinkela_wire_6675)
    );

    bfr new_Jinkela_buffer_5463 (
        .din(new_Jinkela_wire_6564),
        .dout(new_Jinkela_wire_6565)
    );

    spl4L new_Jinkela_splitter_232 (
        .a(n_0690_),
        .d(new_Jinkela_wire_4508),
        .b(new_Jinkela_wire_4509),
        .e(new_Jinkela_wire_4510),
        .c(new_Jinkela_wire_4511)
    );

    bfr new_Jinkela_buffer_7576 (
        .din(n_0021_),
        .dout(new_Jinkela_wire_9498)
    );

    bfr new_Jinkela_buffer_7567 (
        .din(new_Jinkela_wire_9486),
        .dout(new_Jinkela_wire_9487)
    );

    bfr new_Jinkela_buffer_3816 (
        .din(new_Jinkela_wire_4449),
        .dout(new_Jinkela_wire_4450)
    );

    bfr new_Jinkela_buffer_5469 (
        .din(new_Jinkela_wire_6570),
        .dout(new_Jinkela_wire_6571)
    );

    bfr new_Jinkela_buffer_5464 (
        .din(new_Jinkela_wire_6565),
        .dout(new_Jinkela_wire_6566)
    );

    spl2 new_Jinkela_splitter_768 (
        .a(n_1246_),
        .b(new_Jinkela_wire_9496),
        .c(new_Jinkela_wire_9497)
    );

    bfr new_Jinkela_buffer_3854 (
        .din(new_Jinkela_wire_4489),
        .dout(new_Jinkela_wire_4490)
    );

    bfr new_Jinkela_buffer_5503 (
        .din(new_Jinkela_wire_6607),
        .dout(new_Jinkela_wire_6608)
    );

    bfr new_Jinkela_buffer_3817 (
        .din(new_Jinkela_wire_4450),
        .dout(new_Jinkela_wire_4451)
    );

    bfr new_Jinkela_buffer_7568 (
        .din(new_Jinkela_wire_9487),
        .dout(new_Jinkela_wire_9488)
    );

    bfr new_Jinkela_buffer_5470 (
        .din(new_Jinkela_wire_6571),
        .dout(new_Jinkela_wire_6572)
    );

    bfr new_Jinkela_buffer_5536 (
        .din(new_Jinkela_wire_6640),
        .dout(new_Jinkela_wire_6641)
    );

    bfr new_Jinkela_buffer_3818 (
        .din(new_Jinkela_wire_4451),
        .dout(new_Jinkela_wire_4452)
    );

    bfr new_Jinkela_buffer_7569 (
        .din(new_Jinkela_wire_9488),
        .dout(new_Jinkela_wire_9489)
    );

    bfr new_Jinkela_buffer_5471 (
        .din(new_Jinkela_wire_6572),
        .dout(new_Jinkela_wire_6573)
    );

    spl2 new_Jinkela_splitter_231 (
        .a(n_1211_),
        .b(new_Jinkela_wire_4506),
        .c(new_Jinkela_wire_4507)
    );

    bfr new_Jinkela_buffer_3855 (
        .din(new_Jinkela_wire_4490),
        .dout(new_Jinkela_wire_4491)
    );

    bfr new_Jinkela_buffer_7577 (
        .din(new_net_2578),
        .dout(new_Jinkela_wire_9499)
    );

    bfr new_Jinkela_buffer_5504 (
        .din(new_Jinkela_wire_6608),
        .dout(new_Jinkela_wire_6609)
    );

    bfr new_Jinkela_buffer_3819 (
        .din(new_Jinkela_wire_4452),
        .dout(new_Jinkela_wire_4453)
    );

    bfr new_Jinkela_buffer_7570 (
        .din(new_Jinkela_wire_9489),
        .dout(new_Jinkela_wire_9490)
    );

    bfr new_Jinkela_buffer_5472 (
        .din(new_Jinkela_wire_6573),
        .dout(new_Jinkela_wire_6574)
    );

    spl2 new_Jinkela_splitter_236 (
        .a(n_0002_),
        .b(new_Jinkela_wire_4523),
        .c(new_Jinkela_wire_4524)
    );

    bfr new_Jinkela_buffer_7578 (
        .din(new_Jinkela_wire_9499),
        .dout(new_Jinkela_wire_9500)
    );

    spl2 new_Jinkela_splitter_432 (
        .a(n_0279_),
        .b(new_Jinkela_wire_6708),
        .c(new_Jinkela_wire_6709)
    );

    bfr new_Jinkela_buffer_3820 (
        .din(new_Jinkela_wire_4453),
        .dout(new_Jinkela_wire_4454)
    );

    bfr new_Jinkela_buffer_7571 (
        .din(new_Jinkela_wire_9490),
        .dout(new_Jinkela_wire_9491)
    );

    bfr new_Jinkela_buffer_5473 (
        .din(new_Jinkela_wire_6574),
        .dout(new_Jinkela_wire_6575)
    );

    bfr new_Jinkela_buffer_3856 (
        .din(new_Jinkela_wire_4491),
        .dout(new_Jinkela_wire_4492)
    );

    spl2 new_Jinkela_splitter_769 (
        .a(n_0246_),
        .b(new_Jinkela_wire_9533),
        .c(new_Jinkela_wire_9534)
    );

    bfr new_Jinkela_buffer_5505 (
        .din(new_Jinkela_wire_6609),
        .dout(new_Jinkela_wire_6610)
    );

    bfr new_Jinkela_buffer_3821 (
        .din(new_Jinkela_wire_4454),
        .dout(new_Jinkela_wire_4455)
    );

    bfr new_Jinkela_buffer_7572 (
        .din(new_Jinkela_wire_9491),
        .dout(new_Jinkela_wire_9492)
    );

    spl3L new_Jinkela_splitter_770 (
        .a(n_0993_),
        .d(new_Jinkela_wire_9536),
        .b(new_Jinkela_wire_9537),
        .c(new_Jinkela_wire_9538)
    );

    bfr new_Jinkela_buffer_7579 (
        .din(new_Jinkela_wire_9500),
        .dout(new_Jinkela_wire_9501)
    );

    bfr new_Jinkela_buffer_5474 (
        .din(new_Jinkela_wire_6575),
        .dout(new_Jinkela_wire_6576)
    );

    bfr new_Jinkela_buffer_5537 (
        .din(new_Jinkela_wire_6641),
        .dout(new_Jinkela_wire_6642)
    );

    bfr new_Jinkela_buffer_3822 (
        .din(new_Jinkela_wire_4455),
        .dout(new_Jinkela_wire_4456)
    );

    bfr new_Jinkela_buffer_7573 (
        .din(new_Jinkela_wire_9492),
        .dout(new_Jinkela_wire_9493)
    );

    bfr new_Jinkela_buffer_5475 (
        .din(new_Jinkela_wire_6576),
        .dout(new_Jinkela_wire_6577)
    );

    spl3L new_Jinkela_splitter_233 (
        .a(n_1030_),
        .d(new_Jinkela_wire_4515),
        .b(new_Jinkela_wire_4516),
        .c(new_Jinkela_wire_4517)
    );

    bfr new_Jinkela_buffer_3857 (
        .din(new_Jinkela_wire_4492),
        .dout(new_Jinkela_wire_4493)
    );

    bfr new_Jinkela_buffer_7598 (
        .din(new_Jinkela_wire_9519),
        .dout(new_Jinkela_wire_9520)
    );

    bfr new_Jinkela_buffer_5506 (
        .din(new_Jinkela_wire_6610),
        .dout(new_Jinkela_wire_6611)
    );

    bfr new_Jinkela_buffer_3823 (
        .din(new_Jinkela_wire_4456),
        .dout(new_Jinkela_wire_4457)
    );

    bfr new_Jinkela_buffer_7574 (
        .din(new_Jinkela_wire_9493),
        .dout(new_Jinkela_wire_9494)
    );

    bfr new_Jinkela_buffer_5476 (
        .din(new_Jinkela_wire_6577),
        .dout(new_Jinkela_wire_6578)
    );

    bfr new_Jinkela_buffer_3869 (
        .din(new_Jinkela_wire_4512),
        .dout(new_Jinkela_wire_4513)
    );

    bfr new_Jinkela_buffer_7580 (
        .din(new_Jinkela_wire_9501),
        .dout(new_Jinkela_wire_9502)
    );

    bfr new_Jinkela_buffer_7575 (
        .din(new_Jinkela_wire_9494),
        .dout(new_Jinkela_wire_9495)
    );

    bfr new_Jinkela_buffer_3824 (
        .din(new_Jinkela_wire_4457),
        .dout(new_Jinkela_wire_4458)
    );

    bfr new_Jinkela_buffer_5477 (
        .din(new_Jinkela_wire_6578),
        .dout(new_Jinkela_wire_6579)
    );

    bfr new_Jinkela_buffer_3871 (
        .din(n_0677_),
        .dout(new_Jinkela_wire_4520)
    );

    bfr new_Jinkela_buffer_3858 (
        .din(new_Jinkela_wire_4493),
        .dout(new_Jinkela_wire_4494)
    );

    bfr new_Jinkela_buffer_7611 (
        .din(new_Jinkela_wire_9534),
        .dout(new_Jinkela_wire_9535)
    );

    spl2 new_Jinkela_splitter_431 (
        .a(n_0315_),
        .b(new_Jinkela_wire_6706),
        .c(new_Jinkela_wire_6707)
    );

    bfr new_Jinkela_buffer_5507 (
        .din(new_Jinkela_wire_6611),
        .dout(new_Jinkela_wire_6612)
    );

    bfr new_Jinkela_buffer_3825 (
        .din(new_Jinkela_wire_4458),
        .dout(new_Jinkela_wire_4459)
    );

    bfr new_Jinkela_buffer_7581 (
        .din(new_Jinkela_wire_9502),
        .dout(new_Jinkela_wire_9503)
    );

    bfr new_Jinkela_buffer_5478 (
        .din(new_Jinkela_wire_6579),
        .dout(new_Jinkela_wire_6580)
    );

    bfr new_Jinkela_buffer_3868 (
        .din(new_Jinkela_wire_4511),
        .dout(new_Jinkela_wire_4512)
    );

    bfr new_Jinkela_buffer_7599 (
        .din(new_Jinkela_wire_9520),
        .dout(new_Jinkela_wire_9521)
    );

    bfr new_Jinkela_buffer_5538 (
        .din(new_Jinkela_wire_6642),
        .dout(new_Jinkela_wire_6643)
    );

    bfr new_Jinkela_buffer_3826 (
        .din(new_Jinkela_wire_4459),
        .dout(new_Jinkela_wire_4460)
    );

    bfr new_Jinkela_buffer_7582 (
        .din(new_Jinkela_wire_9503),
        .dout(new_Jinkela_wire_9504)
    );

    bfr new_Jinkela_buffer_5479 (
        .din(new_Jinkela_wire_6580),
        .dout(new_Jinkela_wire_6581)
    );

    bfr new_Jinkela_buffer_3859 (
        .din(new_Jinkela_wire_4494),
        .dout(new_Jinkela_wire_4495)
    );

    bfr new_Jinkela_buffer_5508 (
        .din(new_Jinkela_wire_6612),
        .dout(new_Jinkela_wire_6613)
    );

    bfr new_Jinkela_buffer_3827 (
        .din(new_Jinkela_wire_4460),
        .dout(new_Jinkela_wire_4461)
    );

    bfr new_Jinkela_buffer_7583 (
        .din(new_Jinkela_wire_9504),
        .dout(new_Jinkela_wire_9505)
    );

    bfr new_Jinkela_buffer_7600 (
        .din(new_Jinkela_wire_9521),
        .dout(new_Jinkela_wire_9522)
    );

    bfr new_Jinkela_buffer_5480 (
        .din(new_Jinkela_wire_6581),
        .dout(new_Jinkela_wire_6582)
    );

    bfr new_Jinkela_buffer_5565 (
        .din(new_Jinkela_wire_6675),
        .dout(new_Jinkela_wire_6676)
    );

    bfr new_Jinkela_buffer_3828 (
        .din(new_Jinkela_wire_4461),
        .dout(new_Jinkela_wire_4462)
    );

    bfr new_Jinkela_buffer_7584 (
        .din(new_Jinkela_wire_9505),
        .dout(new_Jinkela_wire_9506)
    );

    bfr new_Jinkela_buffer_5481 (
        .din(new_Jinkela_wire_6582),
        .dout(new_Jinkela_wire_6583)
    );

    bfr new_Jinkela_buffer_3860 (
        .din(new_Jinkela_wire_4495),
        .dout(new_Jinkela_wire_4496)
    );

    bfr new_Jinkela_buffer_7612 (
        .din(n_0288_),
        .dout(new_Jinkela_wire_9541)
    );

    bfr new_Jinkela_buffer_5509 (
        .din(new_Jinkela_wire_6613),
        .dout(new_Jinkela_wire_6614)
    );

    bfr new_Jinkela_buffer_3829 (
        .din(new_Jinkela_wire_4462),
        .dout(new_Jinkela_wire_4463)
    );

    bfr new_Jinkela_buffer_7585 (
        .din(new_Jinkela_wire_9506),
        .dout(new_Jinkela_wire_9507)
    );

    spl2 new_Jinkela_splitter_771 (
        .a(new_Jinkela_wire_9538),
        .b(new_Jinkela_wire_9539),
        .c(new_Jinkela_wire_9540)
    );

    bfr new_Jinkela_buffer_5482 (
        .din(new_Jinkela_wire_6583),
        .dout(new_Jinkela_wire_6584)
    );

    bfr new_Jinkela_buffer_3873 (
        .din(n_0270_),
        .dout(new_Jinkela_wire_4526)
    );

    bfr new_Jinkela_buffer_7601 (
        .din(new_Jinkela_wire_9522),
        .dout(new_Jinkela_wire_9523)
    );

    bfr new_Jinkela_buffer_5539 (
        .din(new_Jinkela_wire_6643),
        .dout(new_Jinkela_wire_6644)
    );

    bfr new_Jinkela_buffer_3830 (
        .din(new_Jinkela_wire_4463),
        .dout(new_Jinkela_wire_4464)
    );

    bfr new_Jinkela_buffer_7586 (
        .din(new_Jinkela_wire_9507),
        .dout(new_Jinkela_wire_9508)
    );

    bfr new_Jinkela_buffer_5483 (
        .din(new_Jinkela_wire_6584),
        .dout(new_Jinkela_wire_6585)
    );

    spl2 new_Jinkela_splitter_234 (
        .a(new_Jinkela_wire_4517),
        .b(new_Jinkela_wire_4518),
        .c(new_Jinkela_wire_4519)
    );

    bfr new_Jinkela_buffer_3861 (
        .din(new_Jinkela_wire_4496),
        .dout(new_Jinkela_wire_4497)
    );

    bfr new_Jinkela_buffer_5510 (
        .din(new_Jinkela_wire_6614),
        .dout(new_Jinkela_wire_6615)
    );

    bfr new_Jinkela_buffer_3831 (
        .din(new_Jinkela_wire_4464),
        .dout(new_Jinkela_wire_4465)
    );

    bfr new_Jinkela_buffer_7587 (
        .din(new_Jinkela_wire_9508),
        .dout(new_Jinkela_wire_9509)
    );

    bfr new_Jinkela_buffer_7613 (
        .din(new_Jinkela_wire_9541),
        .dout(new_Jinkela_wire_9542)
    );

    bfr new_Jinkela_buffer_5484 (
        .din(new_Jinkela_wire_6585),
        .dout(new_Jinkela_wire_6586)
    );

    bfr new_Jinkela_buffer_3870 (
        .din(new_Jinkela_wire_4513),
        .dout(new_Jinkela_wire_4514)
    );

    bfr new_Jinkela_buffer_7602 (
        .din(new_Jinkela_wire_9523),
        .dout(new_Jinkela_wire_9524)
    );

    bfr new_Jinkela_buffer_5595 (
        .din(new_net_2515),
        .dout(new_Jinkela_wire_6710)
    );

    bfr new_Jinkela_buffer_3832 (
        .din(new_Jinkela_wire_4465),
        .dout(new_Jinkela_wire_4466)
    );

    bfr new_Jinkela_buffer_7588 (
        .din(new_Jinkela_wire_9509),
        .dout(new_Jinkela_wire_9510)
    );

    bfr new_Jinkela_buffer_5485 (
        .din(new_Jinkela_wire_6586),
        .dout(new_Jinkela_wire_6587)
    );

    bfr new_Jinkela_buffer_3862 (
        .din(new_Jinkela_wire_4497),
        .dout(new_Jinkela_wire_4498)
    );

    bfr new_Jinkela_buffer_5511 (
        .din(new_Jinkela_wire_6615),
        .dout(new_Jinkela_wire_6616)
    );

    bfr new_Jinkela_buffer_3833 (
        .din(new_Jinkela_wire_4466),
        .dout(new_Jinkela_wire_4467)
    );

    bfr new_Jinkela_buffer_7589 (
        .din(new_Jinkela_wire_9510),
        .dout(new_Jinkela_wire_9511)
    );

    bfr new_Jinkela_buffer_5486 (
        .din(new_Jinkela_wire_6587),
        .dout(new_Jinkela_wire_6588)
    );

    spl2 new_Jinkela_splitter_235 (
        .a(n_0886_),
        .b(new_Jinkela_wire_4521),
        .c(new_Jinkela_wire_4522)
    );

    bfr new_Jinkela_buffer_7603 (
        .din(new_Jinkela_wire_9524),
        .dout(new_Jinkela_wire_9525)
    );

    bfr new_Jinkela_buffer_5540 (
        .din(new_Jinkela_wire_6644),
        .dout(new_Jinkela_wire_6645)
    );

    bfr new_Jinkela_buffer_3834 (
        .din(new_Jinkela_wire_4467),
        .dout(new_Jinkela_wire_4468)
    );

    bfr new_Jinkela_buffer_7590 (
        .din(new_Jinkela_wire_9511),
        .dout(new_Jinkela_wire_9512)
    );

    bfr new_Jinkela_buffer_5487 (
        .din(new_Jinkela_wire_6588),
        .dout(new_Jinkela_wire_6589)
    );

    bfr new_Jinkela_buffer_3863 (
        .din(new_Jinkela_wire_4498),
        .dout(new_Jinkela_wire_4499)
    );

    bfr new_Jinkela_buffer_7614 (
        .din(n_1252_),
        .dout(new_Jinkela_wire_9548)
    );

    bfr new_Jinkela_buffer_5512 (
        .din(new_Jinkela_wire_6616),
        .dout(new_Jinkela_wire_6617)
    );

    bfr new_Jinkela_buffer_3835 (
        .din(new_Jinkela_wire_4468),
        .dout(new_Jinkela_wire_4469)
    );

    bfr new_Jinkela_buffer_7591 (
        .din(new_Jinkela_wire_9512),
        .dout(new_Jinkela_wire_9513)
    );

    spl3L new_Jinkela_splitter_772 (
        .a(n_1078_),
        .d(new_Jinkela_wire_9543),
        .b(new_Jinkela_wire_9544),
        .c(new_Jinkela_wire_9545)
    );

    bfr new_Jinkela_buffer_7604 (
        .din(new_Jinkela_wire_9525),
        .dout(new_Jinkela_wire_9526)
    );

    bfr new_Jinkela_buffer_5488 (
        .din(new_Jinkela_wire_6589),
        .dout(new_Jinkela_wire_6590)
    );

    and_ii n_1569_ (
        .a(new_Jinkela_wire_7458),
        .b(new_Jinkela_wire_9303),
        .c(n_0837_)
    );

    or_bb n_2283_ (
        .a(n_0160_),
        .b(n_0159_),
        .c(new_net_2547)
    );

    bfr new_Jinkela_buffer_6267 (
        .din(new_Jinkela_wire_7640),
        .dout(new_Jinkela_wire_7641)
    );

    and_bb n_1570_ (
        .a(new_Jinkela_wire_7457),
        .b(new_Jinkela_wire_9302),
        .c(n_0838_)
    );

    and_bb n_2284_ (
        .a(new_Jinkela_wire_0),
        .b(new_Jinkela_wire_1699),
        .c(new_net_2499)
    );

    spl2 new_Jinkela_splitter_547 (
        .a(new_Jinkela_wire_7741),
        .b(new_Jinkela_wire_7742),
        .c(new_Jinkela_wire_7743)
    );

    or_bb n_1571_ (
        .a(n_0838_),
        .b(n_0837_),
        .c(n_0839_)
    );

    inv n_2285_ (
        .din(new_Jinkela_wire_350),
        .dout(n_0161_)
    );

    bfr new_Jinkela_buffer_6268 (
        .din(new_Jinkela_wire_7641),
        .dout(new_Jinkela_wire_7642)
    );

    and_ii n_1572_ (
        .a(new_Jinkela_wire_8191),
        .b(new_Jinkela_wire_7240),
        .c(n_0840_)
    );

    and_bb n_2286_ (
        .a(new_Jinkela_wire_3519),
        .b(new_Jinkela_wire_2976),
        .c(n_0162_)
    );

    bfr new_Jinkela_buffer_6302 (
        .din(new_Jinkela_wire_7679),
        .dout(new_Jinkela_wire_7680)
    );

    and_bb n_1573_ (
        .a(new_Jinkela_wire_8190),
        .b(new_Jinkela_wire_7239),
        .c(n_0841_)
    );

    or_ii n_2287_ (
        .a(new_Jinkela_wire_6949),
        .b(new_Jinkela_wire_5252),
        .c(n_0163_)
    );

    bfr new_Jinkela_buffer_6269 (
        .din(new_Jinkela_wire_7642),
        .dout(new_Jinkela_wire_7643)
    );

    and_ii n_1574_ (
        .a(n_0841_),
        .b(n_0840_),
        .c(n_0842_)
    );

    and_bb n_2288_ (
        .a(new_Jinkela_wire_6947),
        .b(new_Jinkela_wire_1909),
        .c(n_0164_)
    );

    bfr new_Jinkela_buffer_6318 (
        .din(new_Jinkela_wire_7699),
        .dout(new_Jinkela_wire_7700)
    );

    or_bi n_1575_ (
        .a(new_Jinkela_wire_3859),
        .b(new_Jinkela_wire_8997),
        .c(n_0843_)
    );

    and_bi n_2289_ (
        .a(new_Jinkela_wire_355),
        .b(n_0164_),
        .c(n_0165_)
    );

    bfr new_Jinkela_buffer_6270 (
        .din(new_Jinkela_wire_7643),
        .dout(new_Jinkela_wire_7644)
    );

    and_bi n_1576_ (
        .a(new_Jinkela_wire_3858),
        .b(new_Jinkela_wire_8996),
        .c(n_0844_)
    );

    and_bb n_2290_ (
        .a(new_Jinkela_wire_3518),
        .b(new_Jinkela_wire_1904),
        .c(n_0166_)
    );

    bfr new_Jinkela_buffer_6303 (
        .din(new_Jinkela_wire_7680),
        .dout(new_Jinkela_wire_7681)
    );

    and_bi n_1577_ (
        .a(n_0843_),
        .b(n_0844_),
        .c(n_0845_)
    );

    and_bi n_2291_ (
        .a(new_Jinkela_wire_4855),
        .b(new_Jinkela_wire_5251),
        .c(n_0167_)
    );

    bfr new_Jinkela_buffer_6271 (
        .din(new_Jinkela_wire_7644),
        .dout(new_Jinkela_wire_7645)
    );

    and_bb n_1578_ (
        .a(new_Jinkela_wire_783),
        .b(new_Jinkela_wire_1379),
        .c(n_0846_)
    );

    and_bi n_2292_ (
        .a(new_Jinkela_wire_5250),
        .b(new_Jinkela_wire_4854),
        .c(n_0168_)
    );

    spl2 new_Jinkela_splitter_546 (
        .a(new_Jinkela_wire_7738),
        .b(new_Jinkela_wire_7739),
        .c(new_Jinkela_wire_7740)
    );

    and_bi n_1579_ (
        .a(new_Jinkela_wire_1093),
        .b(new_Jinkela_wire_1322),
        .c(n_0847_)
    );

    and_ii n_2293_ (
        .a(new_Jinkela_wire_4680),
        .b(new_Jinkela_wire_8104),
        .c(n_0169_)
    );

    bfr new_Jinkela_buffer_6272 (
        .din(new_Jinkela_wire_7645),
        .dout(new_Jinkela_wire_7646)
    );

    or_bb n_1580_ (
        .a(new_Jinkela_wire_8999),
        .b(new_Jinkela_wire_8820),
        .c(n_0848_)
    );

    and_bi n_2294_ (
        .a(new_Jinkela_wire_10367),
        .b(new_Jinkela_wire_8478),
        .c(n_0170_)
    );

    bfr new_Jinkela_buffer_6319 (
        .din(new_Jinkela_wire_7700),
        .dout(new_Jinkela_wire_7701)
    );

    and_bb n_1581_ (
        .a(new_Jinkela_wire_1830),
        .b(new_Jinkela_wire_1184),
        .c(n_0849_)
    );

    and_ii n_2295_ (
        .a(n_0170_),
        .b(new_Jinkela_wire_3872),
        .c(n_0171_)
    );

    bfr new_Jinkela_buffer_6273 (
        .din(new_Jinkela_wire_7646),
        .dout(new_Jinkela_wire_7647)
    );

    and_bi n_1582_ (
        .a(new_Jinkela_wire_2458),
        .b(new_Jinkela_wire_1372),
        .c(n_0850_)
    );

    or_ii n_2296_ (
        .a(new_Jinkela_wire_5676),
        .b(new_Jinkela_wire_9651),
        .c(n_0172_)
    );

    bfr new_Jinkela_buffer_6354 (
        .din(new_Jinkela_wire_7750),
        .dout(new_Jinkela_wire_7751)
    );

    and_ii n_1583_ (
        .a(new_Jinkela_wire_6518),
        .b(new_Jinkela_wire_4172),
        .c(n_0851_)
    );

    and_ii n_2297_ (
        .a(new_Jinkela_wire_4193),
        .b(new_Jinkela_wire_6196),
        .c(n_0173_)
    );

    bfr new_Jinkela_buffer_6274 (
        .din(new_Jinkela_wire_7647),
        .dout(new_Jinkela_wire_7648)
    );

    or_bb n_1584_ (
        .a(new_Jinkela_wire_4647),
        .b(new_Jinkela_wire_10139),
        .c(n_0852_)
    );

    and_bi n_2298_ (
        .a(new_Jinkela_wire_5976),
        .b(n_0173_),
        .c(n_0174_)
    );

    bfr new_Jinkela_buffer_6320 (
        .din(new_Jinkela_wire_7701),
        .dout(new_Jinkela_wire_7702)
    );

    and_bb n_1585_ (
        .a(new_Jinkela_wire_4645),
        .b(new_Jinkela_wire_10137),
        .c(n_0853_)
    );

    and_bi n_2299_ (
        .a(new_Jinkela_wire_5877),
        .b(new_Jinkela_wire_4232),
        .c(n_0175_)
    );

    spl2 new_Jinkela_splitter_541 (
        .a(new_Jinkela_wire_7648),
        .b(new_Jinkela_wire_7649),
        .c(new_Jinkela_wire_7650)
    );

    and_bi n_1586_ (
        .a(n_0852_),
        .b(n_0853_),
        .c(n_0854_)
    );

    and_bi n_2300_ (
        .a(new_Jinkela_wire_6603),
        .b(n_0175_),
        .c(n_0176_)
    );

    bfr new_Jinkela_buffer_6321 (
        .din(new_Jinkela_wire_7702),
        .dout(new_Jinkela_wire_7703)
    );

    or_ii n_1587_ (
        .a(new_Jinkela_wire_2072),
        .b(new_Jinkela_wire_1359),
        .c(n_0855_)
    );

    or_bb n_2301_ (
        .a(new_Jinkela_wire_7020),
        .b(new_Jinkela_wire_4393),
        .c(n_0177_)
    );

    bfr new_Jinkela_buffer_6357 (
        .din(new_Jinkela_wire_7753),
        .dout(new_Jinkela_wire_7754)
    );

    and_bi n_1588_ (
        .a(new_Jinkela_wire_598),
        .b(new_Jinkela_wire_1226),
        .c(n_0856_)
    );

    and_bi n_2302_ (
        .a(new_Jinkela_wire_9137),
        .b(new_Jinkela_wire_4626),
        .c(n_0178_)
    );

    bfr new_Jinkela_buffer_6356 (
        .din(n_0676_),
        .dout(new_Jinkela_wire_7753)
    );

    and_bi n_1589_ (
        .a(new_Jinkela_wire_5555),
        .b(new_Jinkela_wire_4985),
        .c(n_0857_)
    );

    and_bi n_2303_ (
        .a(new_Jinkela_wire_10627),
        .b(new_Jinkela_wire_4923),
        .c(new_net_2489)
    );

    bfr new_Jinkela_buffer_6322 (
        .din(new_Jinkela_wire_7703),
        .dout(new_Jinkela_wire_7704)
    );

    and_bb n_1590_ (
        .a(new_Jinkela_wire_3362),
        .b(new_Jinkela_wire_1290),
        .c(n_0858_)
    );

    or_bi n_2304_ (
        .a(new_Jinkela_wire_349),
        .b(new_Jinkela_wire_3520),
        .c(n_0179_)
    );

    spl2 new_Jinkela_splitter_552 (
        .a(n_0029_),
        .b(new_Jinkela_wire_7766),
        .c(new_Jinkela_wire_7767)
    );

    spl2 new_Jinkela_splitter_553 (
        .a(n_0055_),
        .b(new_Jinkela_wire_7772),
        .c(new_Jinkela_wire_7773)
    );

    and_bi n_1591_ (
        .a(new_Jinkela_wire_799),
        .b(new_Jinkela_wire_1309),
        .c(n_0859_)
    );

    or_bb n_2305_ (
        .a(new_Jinkela_wire_7682),
        .b(new_Jinkela_wire_7824),
        .c(n_0180_)
    );

    bfr new_Jinkela_buffer_6323 (
        .din(new_Jinkela_wire_7704),
        .dout(new_Jinkela_wire_7705)
    );

    and_ii n_1592_ (
        .a(new_Jinkela_wire_8328),
        .b(new_Jinkela_wire_9767),
        .c(n_0860_)
    );

    and_bb n_2306_ (
        .a(new_Jinkela_wire_10100),
        .b(new_Jinkela_wire_9540),
        .c(n_0181_)
    );

    bfr new_Jinkela_buffer_6355 (
        .din(new_Jinkela_wire_7751),
        .dout(new_Jinkela_wire_7752)
    );

    and_ii n_1593_ (
        .a(new_Jinkela_wire_9923),
        .b(new_Jinkela_wire_10364),
        .c(n_0861_)
    );

    or_bb n_2307_ (
        .a(new_Jinkela_wire_3866),
        .b(new_Jinkela_wire_8289),
        .c(n_0182_)
    );

    bfr new_Jinkela_buffer_6324 (
        .din(new_Jinkela_wire_7705),
        .dout(new_Jinkela_wire_7706)
    );

    and_bb n_1594_ (
        .a(new_Jinkela_wire_9924),
        .b(new_Jinkela_wire_10362),
        .c(n_0862_)
    );

    and_ii n_2308_ (
        .a(new_Jinkela_wire_5640),
        .b(new_Jinkela_wire_4010),
        .c(n_0183_)
    );

    and_ii n_1595_ (
        .a(n_0862_),
        .b(n_0861_),
        .c(n_0863_)
    );

    or_bb n_2309_ (
        .a(new_Jinkela_wire_763),
        .b(new_Jinkela_wire_2586),
        .c(n_0184_)
    );

    bfr new_Jinkela_buffer_6325 (
        .din(new_Jinkela_wire_7706),
        .dout(new_Jinkela_wire_7707)
    );

    or_bb n_1596_ (
        .a(new_Jinkela_wire_9017),
        .b(new_Jinkela_wire_9771),
        .c(n_0864_)
    );

    and_bi n_2310_ (
        .a(new_Jinkela_wire_9380),
        .b(new_Jinkela_wire_8365),
        .c(n_0185_)
    );

    bfr new_Jinkela_buffer_6358 (
        .din(new_Jinkela_wire_7754),
        .dout(new_Jinkela_wire_7755)
    );

    and_bb n_1597_ (
        .a(new_Jinkela_wire_9016),
        .b(new_Jinkela_wire_9770),
        .c(n_0865_)
    );

    and_bi n_2311_ (
        .a(new_Jinkela_wire_769),
        .b(new_Jinkela_wire_9296),
        .c(n_0186_)
    );

    bfr new_Jinkela_buffer_6326 (
        .din(new_Jinkela_wire_7707),
        .dout(new_Jinkela_wire_7708)
    );

    and_bi n_1598_ (
        .a(n_0864_),
        .b(n_0865_),
        .c(n_0866_)
    );

    or_bb n_2312_ (
        .a(n_0186_),
        .b(n_0185_),
        .c(n_0187_)
    );

    spl2 new_Jinkela_splitter_554 (
        .a(n_0451_),
        .b(new_Jinkela_wire_7804),
        .c(new_Jinkela_wire_7805)
    );

    and_bb n_1599_ (
        .a(new_Jinkela_wire_2160),
        .b(new_Jinkela_wire_1293),
        .c(n_0867_)
    );

    or_bb n_2313_ (
        .a(new_Jinkela_wire_10386),
        .b(n_0183_),
        .c(n_0188_)
    );

    bfr new_Jinkela_buffer_6327 (
        .din(new_Jinkela_wire_7708),
        .dout(new_Jinkela_wire_7709)
    );

    and_bi n_1600_ (
        .a(new_Jinkela_wire_359),
        .b(new_Jinkela_wire_1268),
        .c(n_0868_)
    );

    and_bb n_2314_ (
        .a(new_Jinkela_wire_7273),
        .b(new_Jinkela_wire_6786),
        .c(n_0189_)
    );

    bfr new_Jinkela_buffer_6398 (
        .din(n_1340_),
        .dout(new_Jinkela_wire_7806)
    );

    and_ii n_1601_ (
        .a(new_Jinkela_wire_4535),
        .b(new_Jinkela_wire_5502),
        .c(n_0869_)
    );

    and_bb n_2315_ (
        .a(new_Jinkela_wire_5639),
        .b(new_Jinkela_wire_4011),
        .c(n_0190_)
    );

    bfr new_Jinkela_buffer_6328 (
        .din(new_Jinkela_wire_7709),
        .dout(new_Jinkela_wire_7710)
    );

    or_ii n_1602_ (
        .a(new_Jinkela_wire_1705),
        .b(new_Jinkela_wire_1183),
        .c(n_0870_)
    );

    or_bb n_2316_ (
        .a(n_0190_),
        .b(n_0189_),
        .c(n_0191_)
    );

    bfr new_Jinkela_buffer_6359 (
        .din(new_Jinkela_wire_7755),
        .dout(new_Jinkela_wire_7756)
    );

    and_bi n_1603_ (
        .a(new_Jinkela_wire_762),
        .b(new_Jinkela_wire_1361),
        .c(n_0871_)
    );

    and_bi n_2317_ (
        .a(n_0188_),
        .b(n_0191_),
        .c(n_0192_)
    );

    bfr new_Jinkela_buffer_6329 (
        .din(new_Jinkela_wire_7710),
        .dout(new_Jinkela_wire_7711)
    );

    and_bi n_1604_ (
        .a(new_Jinkela_wire_8392),
        .b(new_Jinkela_wire_8276),
        .c(n_0872_)
    );

    and_ii n_2318_ (
        .a(new_Jinkela_wire_7271),
        .b(new_Jinkela_wire_6787),
        .c(n_0193_)
    );

    bfr new_Jinkela_buffer_6365 (
        .din(new_Jinkela_wire_7768),
        .dout(new_Jinkela_wire_7769)
    );

    and_bb n_1605_ (
        .a(new_Jinkela_wire_9765),
        .b(new_Jinkela_wire_5574),
        .c(n_0873_)
    );

    and_ii n_2319_ (
        .a(new_Jinkela_wire_10422),
        .b(new_Jinkela_wire_8193),
        .c(n_0194_)
    );

    bfr new_Jinkela_buffer_6330 (
        .din(new_Jinkela_wire_7711),
        .dout(new_Jinkela_wire_7712)
    );

    and_ii n_1606_ (
        .a(new_Jinkela_wire_9766),
        .b(new_Jinkela_wire_5573),
        .c(n_0874_)
    );

    or_bb n_2320_ (
        .a(n_0194_),
        .b(n_0193_),
        .c(n_0195_)
    );

    bfr new_Jinkela_buffer_6364 (
        .din(new_Jinkela_wire_7767),
        .dout(new_Jinkela_wire_7768)
    );

    spl3L new_Jinkela_splitter_550 (
        .a(new_Jinkela_wire_7756),
        .d(new_Jinkela_wire_7757),
        .b(new_Jinkela_wire_7758),
        .c(new_Jinkela_wire_7759)
    );

    and_ii n_1607_ (
        .a(n_0874_),
        .b(n_0873_),
        .c(n_0875_)
    );

    or_bb n_2321_ (
        .a(new_Jinkela_wire_9148),
        .b(n_0192_),
        .c(n_0196_)
    );

    bfr new_Jinkela_buffer_6331 (
        .din(new_Jinkela_wire_7712),
        .dout(new_Jinkela_wire_7713)
    );

    and_bb n_1608_ (
        .a(new_Jinkela_wire_2901),
        .b(new_Jinkela_wire_1327),
        .c(n_0876_)
    );

    and_bb n_2322_ (
        .a(new_Jinkela_wire_3867),
        .b(new_Jinkela_wire_8288),
        .c(n_0197_)
    );

    and_bi n_1609_ (
        .a(new_Jinkela_wire_3546),
        .b(new_Jinkela_wire_1192),
        .c(n_0877_)
    );

    and_bb n_2323_ (
        .a(new_Jinkela_wire_10419),
        .b(new_Jinkela_wire_8194),
        .c(n_0198_)
    );

    bfr new_Jinkela_buffer_6332 (
        .din(new_Jinkela_wire_7713),
        .dout(new_Jinkela_wire_7714)
    );

    and_ii n_1610_ (
        .a(new_Jinkela_wire_3837),
        .b(new_Jinkela_wire_8383),
        .c(n_0878_)
    );

    or_bb n_2324_ (
        .a(n_0198_),
        .b(n_0197_),
        .c(n_0199_)
    );

    bfr new_Jinkela_buffer_6368 (
        .din(new_Jinkela_wire_7773),
        .dout(new_Jinkela_wire_7774)
    );

    bfr new_Jinkela_buffer_7120 (
        .din(new_Jinkela_wire_8803),
        .dout(new_Jinkela_wire_8804)
    );

    bfr new_Jinkela_buffer_7144 (
        .din(new_Jinkela_wire_8838),
        .dout(new_Jinkela_wire_8839)
    );

    bfr new_Jinkela_buffer_7121 (
        .din(new_Jinkela_wire_8804),
        .dout(new_Jinkela_wire_8805)
    );

    bfr new_Jinkela_buffer_7169 (
        .din(n_0564_),
        .dout(new_Jinkela_wire_8875)
    );

    spl2 new_Jinkela_splitter_684 (
        .a(n_1146_),
        .b(new_Jinkela_wire_8881),
        .c(new_Jinkela_wire_8882)
    );

    bfr new_Jinkela_buffer_7122 (
        .din(new_Jinkela_wire_8805),
        .dout(new_Jinkela_wire_8806)
    );

    bfr new_Jinkela_buffer_7145 (
        .din(new_Jinkela_wire_8839),
        .dout(new_Jinkela_wire_8840)
    );

    bfr new_Jinkela_buffer_7123 (
        .din(new_Jinkela_wire_8806),
        .dout(new_Jinkela_wire_8807)
    );

    bfr new_Jinkela_buffer_7156 (
        .din(new_Jinkela_wire_8857),
        .dout(new_Jinkela_wire_8858)
    );

    bfr new_Jinkela_buffer_7124 (
        .din(new_Jinkela_wire_8807),
        .dout(new_Jinkela_wire_8808)
    );

    bfr new_Jinkela_buffer_7146 (
        .din(new_Jinkela_wire_8840),
        .dout(new_Jinkela_wire_8841)
    );

    bfr new_Jinkela_buffer_7125 (
        .din(new_Jinkela_wire_8808),
        .dout(new_Jinkela_wire_8809)
    );

    bfr new_Jinkela_buffer_7167 (
        .din(new_Jinkela_wire_8872),
        .dout(new_Jinkela_wire_8873)
    );

    spl2 new_Jinkela_splitter_673 (
        .a(new_Jinkela_wire_8809),
        .b(new_Jinkela_wire_8810),
        .c(new_Jinkela_wire_8811)
    );

    bfr new_Jinkela_buffer_7157 (
        .din(new_Jinkela_wire_8858),
        .dout(new_Jinkela_wire_8859)
    );

    bfr new_Jinkela_buffer_7147 (
        .din(new_Jinkela_wire_8841),
        .dout(new_Jinkela_wire_8842)
    );

    bfr new_Jinkela_buffer_7158 (
        .din(new_Jinkela_wire_8859),
        .dout(new_Jinkela_wire_8860)
    );

    spl2 new_Jinkela_splitter_685 (
        .a(n_0585_),
        .b(new_Jinkela_wire_8883),
        .c(new_Jinkela_wire_8884)
    );

    bfr new_Jinkela_buffer_7170 (
        .din(new_Jinkela_wire_8875),
        .dout(new_Jinkela_wire_8876)
    );

    bfr new_Jinkela_buffer_7159 (
        .din(new_Jinkela_wire_8860),
        .dout(new_Jinkela_wire_8861)
    );

    spl2 new_Jinkela_splitter_686 (
        .a(n_1268_),
        .b(new_Jinkela_wire_8885),
        .c(new_Jinkela_wire_8886)
    );

    bfr new_Jinkela_buffer_7160 (
        .din(new_Jinkela_wire_8861),
        .dout(new_Jinkela_wire_8862)
    );

    bfr new_Jinkela_buffer_7171 (
        .din(new_Jinkela_wire_8876),
        .dout(new_Jinkela_wire_8877)
    );

    bfr new_Jinkela_buffer_7161 (
        .din(new_Jinkela_wire_8862),
        .dout(new_Jinkela_wire_8863)
    );

    bfr new_Jinkela_buffer_7162 (
        .din(new_Jinkela_wire_8863),
        .dout(new_Jinkela_wire_8864)
    );

    bfr new_Jinkela_buffer_7174 (
        .din(new_Jinkela_wire_8887),
        .dout(new_Jinkela_wire_8888)
    );

    bfr new_Jinkela_buffer_7172 (
        .din(new_Jinkela_wire_8877),
        .dout(new_Jinkela_wire_8878)
    );

    bfr new_Jinkela_buffer_7163 (
        .din(new_Jinkela_wire_8864),
        .dout(new_Jinkela_wire_8865)
    );

    bfr new_Jinkela_buffer_7164 (
        .din(new_Jinkela_wire_8865),
        .dout(new_Jinkela_wire_8866)
    );

    bfr new_Jinkela_buffer_7173 (
        .din(n_0557_),
        .dout(new_Jinkela_wire_8887)
    );

    spl2 new_Jinkela_splitter_683 (
        .a(new_Jinkela_wire_8878),
        .b(new_Jinkela_wire_8879),
        .c(new_Jinkela_wire_8880)
    );

    bfr new_Jinkela_buffer_7165 (
        .din(new_Jinkela_wire_8866),
        .dout(new_Jinkela_wire_8867)
    );

    bfr new_Jinkela_buffer_7210 (
        .din(n_0640_),
        .dout(new_Jinkela_wire_8924)
    );

    bfr new_Jinkela_buffer_7178 (
        .din(new_net_2543),
        .dout(new_Jinkela_wire_8892)
    );

    bfr new_Jinkela_buffer_7175 (
        .din(new_Jinkela_wire_8888),
        .dout(new_Jinkela_wire_8889)
    );

    bfr new_Jinkela_buffer_7179 (
        .din(new_Jinkela_wire_8892),
        .dout(new_Jinkela_wire_8893)
    );

    bfr new_Jinkela_buffer_7176 (
        .din(new_Jinkela_wire_8889),
        .dout(new_Jinkela_wire_8890)
    );

    spl2 new_Jinkela_splitter_687 (
        .a(n_0572_),
        .b(new_Jinkela_wire_8925),
        .c(new_Jinkela_wire_8926)
    );

    bfr new_Jinkela_buffer_7211 (
        .din(n_0981_),
        .dout(new_Jinkela_wire_8927)
    );

    bfr new_Jinkela_buffer_7177 (
        .din(new_Jinkela_wire_8890),
        .dout(new_Jinkela_wire_8891)
    );

    bfr new_Jinkela_buffer_7180 (
        .din(new_Jinkela_wire_8893),
        .dout(new_Jinkela_wire_8894)
    );

    bfr new_Jinkela_buffer_7181 (
        .din(new_Jinkela_wire_8894),
        .dout(new_Jinkela_wire_8895)
    );

    bfr new_Jinkela_buffer_764 (
        .din(new_Jinkela_wire_824),
        .dout(new_Jinkela_wire_825)
    );

    bfr new_Jinkela_buffer_8311 (
        .din(new_Jinkela_wire_10450),
        .dout(new_Jinkela_wire_10451)
    );

    bfr new_Jinkela_buffer_1015 (
        .din(N121),
        .dout(new_Jinkela_wire_1090)
    );

    bfr new_Jinkela_buffer_1012 (
        .din(new_Jinkela_wire_1086),
        .dout(new_Jinkela_wire_1087)
    );

    bfr new_Jinkela_buffer_8347 (
        .din(new_Jinkela_wire_10486),
        .dout(new_Jinkela_wire_10487)
    );

    bfr new_Jinkela_buffer_765 (
        .din(new_Jinkela_wire_825),
        .dout(new_Jinkela_wire_826)
    );

    bfr new_Jinkela_buffer_8312 (
        .din(new_Jinkela_wire_10451),
        .dout(new_Jinkela_wire_10452)
    );

    bfr new_Jinkela_buffer_824 (
        .din(new_Jinkela_wire_886),
        .dout(new_Jinkela_wire_887)
    );

    spl4L new_Jinkela_splitter_864 (
        .a(n_1310_),
        .d(new_Jinkela_wire_10527),
        .b(new_Jinkela_wire_10528),
        .e(new_Jinkela_wire_10529),
        .c(new_Jinkela_wire_10530)
    );

    bfr new_Jinkela_buffer_766 (
        .din(new_Jinkela_wire_826),
        .dout(new_Jinkela_wire_827)
    );

    bfr new_Jinkela_buffer_8313 (
        .din(new_Jinkela_wire_10452),
        .dout(new_Jinkela_wire_10453)
    );

    bfr new_Jinkela_buffer_886 (
        .din(new_Jinkela_wire_953),
        .dout(new_Jinkela_wire_954)
    );

    bfr new_Jinkela_buffer_8348 (
        .din(new_Jinkela_wire_10487),
        .dout(new_Jinkela_wire_10488)
    );

    bfr new_Jinkela_buffer_767 (
        .din(new_Jinkela_wire_827),
        .dout(new_Jinkela_wire_828)
    );

    bfr new_Jinkela_buffer_8314 (
        .din(new_Jinkela_wire_10453),
        .dout(new_Jinkela_wire_10454)
    );

    spl3L new_Jinkela_splitter_28 (
        .a(new_Jinkela_wire_887),
        .d(new_Jinkela_wire_888),
        .b(new_Jinkela_wire_889),
        .c(new_Jinkela_wire_890)
    );

    bfr new_Jinkela_buffer_768 (
        .din(new_Jinkela_wire_828),
        .dout(new_Jinkela_wire_829)
    );

    bfr new_Jinkela_buffer_8315 (
        .din(new_Jinkela_wire_10454),
        .dout(new_Jinkela_wire_10455)
    );

    bfr new_Jinkela_buffer_8349 (
        .din(new_Jinkela_wire_10488),
        .dout(new_Jinkela_wire_10489)
    );

    bfr new_Jinkela_buffer_769 (
        .din(new_Jinkela_wire_829),
        .dout(new_Jinkela_wire_830)
    );

    bfr new_Jinkela_buffer_8316 (
        .din(new_Jinkela_wire_10455),
        .dout(new_Jinkela_wire_10456)
    );

    bfr new_Jinkela_buffer_825 (
        .din(new_Jinkela_wire_890),
        .dout(new_Jinkela_wire_891)
    );

    spl3L new_Jinkela_splitter_866 (
        .a(n_0915_),
        .d(new_Jinkela_wire_10556),
        .b(new_Jinkela_wire_10557),
        .c(new_Jinkela_wire_10558)
    );

    spl2 new_Jinkela_splitter_861 (
        .a(new_Jinkela_wire_10503),
        .b(new_Jinkela_wire_10504),
        .c(new_Jinkela_wire_10505)
    );

    bfr new_Jinkela_buffer_770 (
        .din(new_Jinkela_wire_830),
        .dout(new_Jinkela_wire_831)
    );

    bfr new_Jinkela_buffer_8317 (
        .din(new_Jinkela_wire_10456),
        .dout(new_Jinkela_wire_10457)
    );

    spl2 new_Jinkela_splitter_29 (
        .a(new_Jinkela_wire_951),
        .b(new_Jinkela_wire_952),
        .c(new_Jinkela_wire_953)
    );

    bfr new_Jinkela_buffer_8350 (
        .din(new_Jinkela_wire_10489),
        .dout(new_Jinkela_wire_10490)
    );

    bfr new_Jinkela_buffer_771 (
        .din(new_Jinkela_wire_831),
        .dout(new_Jinkela_wire_832)
    );

    bfr new_Jinkela_buffer_8318 (
        .din(new_Jinkela_wire_10457),
        .dout(new_Jinkela_wire_10458)
    );

    bfr new_Jinkela_buffer_826 (
        .din(new_Jinkela_wire_891),
        .dout(new_Jinkela_wire_892)
    );

    bfr new_Jinkela_buffer_8362 (
        .din(new_Jinkela_wire_10505),
        .dout(new_Jinkela_wire_10506)
    );

    spl4L new_Jinkela_splitter_863 (
        .a(n_1165_),
        .d(new_Jinkela_wire_10523),
        .b(new_Jinkela_wire_10524),
        .e(new_Jinkela_wire_10525),
        .c(new_Jinkela_wire_10526)
    );

    bfr new_Jinkela_buffer_772 (
        .din(new_Jinkela_wire_832),
        .dout(new_Jinkela_wire_833)
    );

    bfr new_Jinkela_buffer_8319 (
        .din(new_Jinkela_wire_10458),
        .dout(new_Jinkela_wire_10459)
    );

    bfr new_Jinkela_buffer_948 (
        .din(new_Jinkela_wire_1020),
        .dout(new_Jinkela_wire_1021)
    );

    bfr new_Jinkela_buffer_8351 (
        .din(new_Jinkela_wire_10490),
        .dout(new_Jinkela_wire_10491)
    );

    bfr new_Jinkela_buffer_773 (
        .din(new_Jinkela_wire_833),
        .dout(new_Jinkela_wire_834)
    );

    bfr new_Jinkela_buffer_8320 (
        .din(new_Jinkela_wire_10459),
        .dout(new_Jinkela_wire_10460)
    );

    bfr new_Jinkela_buffer_827 (
        .din(new_Jinkela_wire_892),
        .dout(new_Jinkela_wire_893)
    );

    bfr new_Jinkela_buffer_774 (
        .din(new_Jinkela_wire_834),
        .dout(new_Jinkela_wire_835)
    );

    bfr new_Jinkela_buffer_8321 (
        .din(new_Jinkela_wire_10460),
        .dout(new_Jinkela_wire_10461)
    );

    bfr new_Jinkela_buffer_887 (
        .din(new_Jinkela_wire_954),
        .dout(new_Jinkela_wire_955)
    );

    bfr new_Jinkela_buffer_8352 (
        .din(new_Jinkela_wire_10491),
        .dout(new_Jinkela_wire_10492)
    );

    bfr new_Jinkela_buffer_775 (
        .din(new_Jinkela_wire_835),
        .dout(new_Jinkela_wire_836)
    );

    bfr new_Jinkela_buffer_8322 (
        .din(new_Jinkela_wire_10461),
        .dout(new_Jinkela_wire_10462)
    );

    bfr new_Jinkela_buffer_828 (
        .din(new_Jinkela_wire_893),
        .dout(new_Jinkela_wire_894)
    );

    spl2 new_Jinkela_splitter_865 (
        .a(n_0369_),
        .b(new_Jinkela_wire_10554),
        .c(new_Jinkela_wire_10555)
    );

    bfr new_Jinkela_buffer_776 (
        .din(new_Jinkela_wire_836),
        .dout(new_Jinkela_wire_837)
    );

    bfr new_Jinkela_buffer_8323 (
        .din(new_Jinkela_wire_10462),
        .dout(new_Jinkela_wire_10463)
    );

    bfr new_Jinkela_buffer_1019 (
        .din(N78),
        .dout(new_Jinkela_wire_1094)
    );

    bfr new_Jinkela_buffer_8353 (
        .din(new_Jinkela_wire_10492),
        .dout(new_Jinkela_wire_10493)
    );

    bfr new_Jinkela_buffer_777 (
        .din(new_Jinkela_wire_837),
        .dout(new_Jinkela_wire_838)
    );

    bfr new_Jinkela_buffer_8324 (
        .din(new_Jinkela_wire_10463),
        .dout(new_Jinkela_wire_10464)
    );

    bfr new_Jinkela_buffer_829 (
        .din(new_Jinkela_wire_894),
        .dout(new_Jinkela_wire_895)
    );

    bfr new_Jinkela_buffer_8377 (
        .din(new_Jinkela_wire_10530),
        .dout(new_Jinkela_wire_10531)
    );

    bfr new_Jinkela_buffer_8363 (
        .din(new_Jinkela_wire_10506),
        .dout(new_Jinkela_wire_10507)
    );

    bfr new_Jinkela_buffer_778 (
        .din(new_Jinkela_wire_838),
        .dout(new_Jinkela_wire_839)
    );

    bfr new_Jinkela_buffer_8325 (
        .din(new_Jinkela_wire_10464),
        .dout(new_Jinkela_wire_10465)
    );

    bfr new_Jinkela_buffer_888 (
        .din(new_Jinkela_wire_955),
        .dout(new_Jinkela_wire_956)
    );

    bfr new_Jinkela_buffer_8354 (
        .din(new_Jinkela_wire_10493),
        .dout(new_Jinkela_wire_10494)
    );

    bfr new_Jinkela_buffer_779 (
        .din(new_Jinkela_wire_839),
        .dout(new_Jinkela_wire_840)
    );

    bfr new_Jinkela_buffer_8326 (
        .din(new_Jinkela_wire_10465),
        .dout(new_Jinkela_wire_10466)
    );

    bfr new_Jinkela_buffer_830 (
        .din(new_Jinkela_wire_895),
        .dout(new_Jinkela_wire_896)
    );

    spl3L new_Jinkela_splitter_868 (
        .a(n_1213_),
        .d(new_Jinkela_wire_10561),
        .b(new_Jinkela_wire_10562),
        .c(new_Jinkela_wire_10563)
    );

    bfr new_Jinkela_buffer_780 (
        .din(new_Jinkela_wire_840),
        .dout(new_Jinkela_wire_841)
    );

    bfr new_Jinkela_buffer_8327 (
        .din(new_Jinkela_wire_10466),
        .dout(new_Jinkela_wire_10467)
    );

    spl2 new_Jinkela_splitter_32 (
        .a(new_Jinkela_wire_1021),
        .b(new_Jinkela_wire_1022),
        .c(new_Jinkela_wire_1023)
    );

    bfr new_Jinkela_buffer_8355 (
        .din(new_Jinkela_wire_10494),
        .dout(new_Jinkela_wire_10495)
    );

    bfr new_Jinkela_buffer_781 (
        .din(new_Jinkela_wire_841),
        .dout(new_Jinkela_wire_842)
    );

    bfr new_Jinkela_buffer_8328 (
        .din(new_Jinkela_wire_10467),
        .dout(new_Jinkela_wire_10468)
    );

    bfr new_Jinkela_buffer_831 (
        .din(new_Jinkela_wire_896),
        .dout(new_Jinkela_wire_897)
    );

    spl2 new_Jinkela_splitter_862 (
        .a(new_Jinkela_wire_10507),
        .b(new_Jinkela_wire_10508),
        .c(new_Jinkela_wire_10509)
    );

    bfr new_Jinkela_buffer_782 (
        .din(new_Jinkela_wire_842),
        .dout(new_Jinkela_wire_843)
    );

    bfr new_Jinkela_buffer_8329 (
        .din(new_Jinkela_wire_10468),
        .dout(new_Jinkela_wire_10469)
    );

    spl3L new_Jinkela_splitter_30 (
        .a(new_Jinkela_wire_956),
        .d(new_Jinkela_wire_957),
        .b(new_Jinkela_wire_958),
        .c(new_Jinkela_wire_959)
    );

    bfr new_Jinkela_buffer_8356 (
        .din(new_Jinkela_wire_10495),
        .dout(new_Jinkela_wire_10496)
    );

    bfr new_Jinkela_buffer_783 (
        .din(new_Jinkela_wire_843),
        .dout(new_Jinkela_wire_844)
    );

    bfr new_Jinkela_buffer_8330 (
        .din(new_Jinkela_wire_10469),
        .dout(new_Jinkela_wire_10470)
    );

    bfr new_Jinkela_buffer_832 (
        .din(new_Jinkela_wire_897),
        .dout(new_Jinkela_wire_898)
    );

    bfr new_Jinkela_buffer_8364 (
        .din(new_Jinkela_wire_10509),
        .dout(new_Jinkela_wire_10510)
    );

    bfr new_Jinkela_buffer_784 (
        .din(new_Jinkela_wire_844),
        .dout(new_Jinkela_wire_845)
    );

    bfr new_Jinkela_buffer_8331 (
        .din(new_Jinkela_wire_10470),
        .dout(new_Jinkela_wire_10471)
    );

    bfr new_Jinkela_buffer_949 (
        .din(new_Jinkela_wire_1023),
        .dout(new_Jinkela_wire_1024)
    );

    bfr new_Jinkela_buffer_8357 (
        .din(new_Jinkela_wire_10496),
        .dout(new_Jinkela_wire_10497)
    );

    bfr new_Jinkela_buffer_5566 (
        .din(new_Jinkela_wire_6676),
        .dout(new_Jinkela_wire_6677)
    );

    bfr new_Jinkela_buffer_5489 (
        .din(new_Jinkela_wire_6590),
        .dout(new_Jinkela_wire_6591)
    );

    bfr new_Jinkela_buffer_5513 (
        .din(new_Jinkela_wire_6617),
        .dout(new_Jinkela_wire_6618)
    );

    bfr new_Jinkela_buffer_5490 (
        .din(new_Jinkela_wire_6591),
        .dout(new_Jinkela_wire_6592)
    );

    bfr new_Jinkela_buffer_5541 (
        .din(new_Jinkela_wire_6645),
        .dout(new_Jinkela_wire_6646)
    );

    bfr new_Jinkela_buffer_5491 (
        .din(new_Jinkela_wire_6592),
        .dout(new_Jinkela_wire_6593)
    );

    bfr new_Jinkela_buffer_5514 (
        .din(new_Jinkela_wire_6618),
        .dout(new_Jinkela_wire_6619)
    );

    bfr new_Jinkela_buffer_5492 (
        .din(new_Jinkela_wire_6593),
        .dout(new_Jinkela_wire_6594)
    );

    spl3L new_Jinkela_splitter_434 (
        .a(n_0001_),
        .d(new_Jinkela_wire_6745),
        .b(new_Jinkela_wire_6746),
        .c(new_Jinkela_wire_6747)
    );

    bfr new_Jinkela_buffer_5493 (
        .din(new_Jinkela_wire_6594),
        .dout(new_Jinkela_wire_6595)
    );

    bfr new_Jinkela_buffer_5596 (
        .din(new_Jinkela_wire_6710),
        .dout(new_Jinkela_wire_6711)
    );

    bfr new_Jinkela_buffer_5515 (
        .din(new_Jinkela_wire_6619),
        .dout(new_Jinkela_wire_6620)
    );

    bfr new_Jinkela_buffer_5494 (
        .din(new_Jinkela_wire_6595),
        .dout(new_Jinkela_wire_6596)
    );

    bfr new_Jinkela_buffer_5542 (
        .din(new_Jinkela_wire_6646),
        .dout(new_Jinkela_wire_6647)
    );

    bfr new_Jinkela_buffer_5495 (
        .din(new_Jinkela_wire_6596),
        .dout(new_Jinkela_wire_6597)
    );

    bfr new_Jinkela_buffer_5516 (
        .din(new_Jinkela_wire_6620),
        .dout(new_Jinkela_wire_6621)
    );

    bfr new_Jinkela_buffer_5496 (
        .din(new_Jinkela_wire_6597),
        .dout(new_Jinkela_wire_6598)
    );

    bfr new_Jinkela_buffer_5567 (
        .din(new_Jinkela_wire_6677),
        .dout(new_Jinkela_wire_6678)
    );

    bfr new_Jinkela_buffer_5497 (
        .din(new_Jinkela_wire_6598),
        .dout(new_Jinkela_wire_6599)
    );

    bfr new_Jinkela_buffer_5517 (
        .din(new_Jinkela_wire_6621),
        .dout(new_Jinkela_wire_6622)
    );

    bfr new_Jinkela_buffer_5498 (
        .din(new_Jinkela_wire_6599),
        .dout(new_Jinkela_wire_6600)
    );

    bfr new_Jinkela_buffer_5543 (
        .din(new_Jinkela_wire_6647),
        .dout(new_Jinkela_wire_6648)
    );

    bfr new_Jinkela_buffer_5499 (
        .din(new_Jinkela_wire_6600),
        .dout(new_Jinkela_wire_6601)
    );

    bfr new_Jinkela_buffer_5518 (
        .din(new_Jinkela_wire_6622),
        .dout(new_Jinkela_wire_6623)
    );

    bfr new_Jinkela_buffer_5500 (
        .din(new_Jinkela_wire_6601),
        .dout(new_Jinkela_wire_6602)
    );

    bfr new_Jinkela_buffer_5501 (
        .din(new_Jinkela_wire_6602),
        .dout(new_Jinkela_wire_6603)
    );

    spl3L new_Jinkela_splitter_433 (
        .a(n_0727_),
        .d(new_Jinkela_wire_6742),
        .b(new_Jinkela_wire_6743),
        .c(new_Jinkela_wire_6744)
    );

    bfr new_Jinkela_buffer_5519 (
        .din(new_Jinkela_wire_6623),
        .dout(new_Jinkela_wire_6624)
    );

    bfr new_Jinkela_buffer_5544 (
        .din(new_Jinkela_wire_6648),
        .dout(new_Jinkela_wire_6649)
    );

    bfr new_Jinkela_buffer_5520 (
        .din(new_Jinkela_wire_6624),
        .dout(new_Jinkela_wire_6625)
    );

    bfr new_Jinkela_buffer_5568 (
        .din(new_Jinkela_wire_6678),
        .dout(new_Jinkela_wire_6679)
    );

    bfr new_Jinkela_buffer_5521 (
        .din(new_Jinkela_wire_6625),
        .dout(new_Jinkela_wire_6626)
    );

    bfr new_Jinkela_buffer_5545 (
        .din(new_Jinkela_wire_6649),
        .dout(new_Jinkela_wire_6650)
    );

    bfr new_Jinkela_buffer_5522 (
        .din(new_Jinkela_wire_6626),
        .dout(new_Jinkela_wire_6627)
    );

    bfr new_Jinkela_buffer_5523 (
        .din(new_Jinkela_wire_6627),
        .dout(new_Jinkela_wire_6628)
    );

    bfr new_Jinkela_buffer_5546 (
        .din(new_Jinkela_wire_6650),
        .dout(new_Jinkela_wire_6651)
    );

    bfr new_Jinkela_buffer_5524 (
        .din(new_Jinkela_wire_6628),
        .dout(new_Jinkela_wire_6629)
    );

    bfr new_Jinkela_buffer_1450 (
        .din(N80),
        .dout(new_Jinkela_wire_1783)
    );

    bfr new_Jinkela_buffer_5569 (
        .din(new_Jinkela_wire_6679),
        .dout(new_Jinkela_wire_6680)
    );

    bfr new_Jinkela_buffer_5525 (
        .din(new_Jinkela_wire_6629),
        .dout(new_Jinkela_wire_6630)
    );

    bfr new_Jinkela_buffer_5547 (
        .din(new_Jinkela_wire_6651),
        .dout(new_Jinkela_wire_6652)
    );

    bfr new_Jinkela_buffer_5526 (
        .din(new_Jinkela_wire_6630),
        .dout(new_Jinkela_wire_6631)
    );

    bfr new_Jinkela_buffer_5644 (
        .din(n_0757_),
        .dout(new_Jinkela_wire_6767)
    );

    bfr new_Jinkela_buffer_2045 (
        .din(new_Jinkela_wire_2414),
        .dout(new_Jinkela_wire_2415)
    );

    spl2 new_Jinkela_splitter_123 (
        .a(N367),
        .b(new_Jinkela_wire_2556),
        .c(new_Jinkela_wire_2557)
    );

    bfr new_Jinkela_buffer_2046 (
        .din(new_Jinkela_wire_2415),
        .dout(new_Jinkela_wire_2416)
    );

    bfr new_Jinkela_buffer_2111 (
        .din(new_Jinkela_wire_2480),
        .dout(new_Jinkela_wire_2481)
    );

    bfr new_Jinkela_buffer_2174 (
        .din(new_Jinkela_wire_2548),
        .dout(new_Jinkela_wire_2549)
    );

    bfr new_Jinkela_buffer_2047 (
        .din(new_Jinkela_wire_2416),
        .dout(new_Jinkela_wire_2417)
    );

    bfr new_Jinkela_buffer_2110 (
        .din(new_Jinkela_wire_2479),
        .dout(new_Jinkela_wire_2480)
    );

    bfr new_Jinkela_buffer_2048 (
        .din(new_Jinkela_wire_2417),
        .dout(new_Jinkela_wire_2418)
    );

    spl2 new_Jinkela_splitter_121 (
        .a(new_Jinkela_wire_2481),
        .b(new_Jinkela_wire_2482),
        .c(new_Jinkela_wire_2483)
    );

    bfr new_Jinkela_buffer_2049 (
        .din(new_Jinkela_wire_2418),
        .dout(new_Jinkela_wire_2419)
    );

    bfr new_Jinkela_buffer_2112 (
        .din(new_Jinkela_wire_2483),
        .dout(new_Jinkela_wire_2484)
    );

    bfr new_Jinkela_buffer_2050 (
        .din(new_Jinkela_wire_2419),
        .dout(new_Jinkela_wire_2420)
    );

    spl2 new_Jinkela_splitter_126 (
        .a(N70),
        .b(new_Jinkela_wire_2586),
        .c(new_Jinkela_wire_2587)
    );

    bfr new_Jinkela_buffer_2051 (
        .din(new_Jinkela_wire_2420),
        .dout(new_Jinkela_wire_2421)
    );

    bfr new_Jinkela_buffer_2175 (
        .din(new_Jinkela_wire_2549),
        .dout(new_Jinkela_wire_2550)
    );

    bfr new_Jinkela_buffer_2052 (
        .din(new_Jinkela_wire_2421),
        .dout(new_Jinkela_wire_2422)
    );

    bfr new_Jinkela_buffer_2178 (
        .din(new_Jinkela_wire_2552),
        .dout(new_Jinkela_wire_2553)
    );

    bfr new_Jinkela_buffer_2053 (
        .din(new_Jinkela_wire_2422),
        .dout(new_Jinkela_wire_2423)
    );

    bfr new_Jinkela_buffer_2113 (
        .din(new_Jinkela_wire_2484),
        .dout(new_Jinkela_wire_2485)
    );

    bfr new_Jinkela_buffer_2054 (
        .din(new_Jinkela_wire_2423),
        .dout(new_Jinkela_wire_2424)
    );

    bfr new_Jinkela_buffer_2176 (
        .din(new_Jinkela_wire_2550),
        .dout(new_Jinkela_wire_2551)
    );

    bfr new_Jinkela_buffer_2055 (
        .din(new_Jinkela_wire_2424),
        .dout(new_Jinkela_wire_2425)
    );

    bfr new_Jinkela_buffer_2114 (
        .din(new_Jinkela_wire_2485),
        .dout(new_Jinkela_wire_2486)
    );

    bfr new_Jinkela_buffer_2056 (
        .din(new_Jinkela_wire_2425),
        .dout(new_Jinkela_wire_2426)
    );

    bfr new_Jinkela_buffer_2181 (
        .din(new_Jinkela_wire_2557),
        .dout(new_Jinkela_wire_2558)
    );

    bfr new_Jinkela_buffer_2057 (
        .din(new_Jinkela_wire_2426),
        .dout(new_Jinkela_wire_2427)
    );

    spl3L new_Jinkela_splitter_122 (
        .a(new_Jinkela_wire_2486),
        .d(new_Jinkela_wire_2487),
        .b(new_Jinkela_wire_2488),
        .c(new_Jinkela_wire_2489)
    );

    bfr new_Jinkela_buffer_2058 (
        .din(new_Jinkela_wire_2427),
        .dout(new_Jinkela_wire_2428)
    );

    bfr new_Jinkela_buffer_2179 (
        .din(new_Jinkela_wire_2553),
        .dout(new_Jinkela_wire_2554)
    );

    bfr new_Jinkela_buffer_2059 (
        .din(new_Jinkela_wire_2428),
        .dout(new_Jinkela_wire_2429)
    );

    bfr new_Jinkela_buffer_2115 (
        .din(new_Jinkela_wire_2489),
        .dout(new_Jinkela_wire_2490)
    );

    bfr new_Jinkela_buffer_2060 (
        .din(new_Jinkela_wire_2429),
        .dout(new_Jinkela_wire_2430)
    );

    spl2 new_Jinkela_splitter_127 (
        .a(N277),
        .b(new_Jinkela_wire_2591),
        .c(new_Jinkela_wire_2592)
    );

    bfr new_Jinkela_buffer_2061 (
        .din(new_Jinkela_wire_2430),
        .dout(new_Jinkela_wire_2431)
    );

    bfr new_Jinkela_buffer_2116 (
        .din(new_Jinkela_wire_2490),
        .dout(new_Jinkela_wire_2491)
    );

    bfr new_Jinkela_buffer_2062 (
        .din(new_Jinkela_wire_2431),
        .dout(new_Jinkela_wire_2432)
    );

    bfr new_Jinkela_buffer_2180 (
        .din(new_Jinkela_wire_2554),
        .dout(new_Jinkela_wire_2555)
    );

    bfr new_Jinkela_buffer_2063 (
        .din(new_Jinkela_wire_2432),
        .dout(new_Jinkela_wire_2433)
    );

    bfr new_Jinkela_buffer_2117 (
        .din(new_Jinkela_wire_2491),
        .dout(new_Jinkela_wire_2492)
    );

    bfr new_Jinkela_buffer_2064 (
        .din(new_Jinkela_wire_2433),
        .dout(new_Jinkela_wire_2434)
    );

    bfr new_Jinkela_buffer_2201 (
        .din(N66),
        .dout(new_Jinkela_wire_2582)
    );

    bfr new_Jinkela_buffer_2065 (
        .din(new_Jinkela_wire_2434),
        .dout(new_Jinkela_wire_2435)
    );

    bfr new_Jinkela_buffer_2118 (
        .din(new_Jinkela_wire_2492),
        .dout(new_Jinkela_wire_2493)
    );

    bfr new_Jinkela_buffer_4653 (
        .din(new_Jinkela_wire_5533),
        .dout(new_Jinkela_wire_5534)
    );

    bfr new_Jinkela_buffer_3082 (
        .din(new_Jinkela_wire_3511),
        .dout(new_Jinkela_wire_3512)
    );

    bfr new_Jinkela_buffer_8332 (
        .din(new_Jinkela_wire_10471),
        .dout(new_Jinkela_wire_10472)
    );

    bfr new_Jinkela_buffer_2958 (
        .din(new_Jinkela_wire_3385),
        .dout(new_Jinkela_wire_3386)
    );

    bfr new_Jinkela_buffer_8378 (
        .din(new_Jinkela_wire_10531),
        .dout(new_Jinkela_wire_10532)
    );

    bfr new_Jinkela_buffer_4654 (
        .din(new_Jinkela_wire_5534),
        .dout(new_Jinkela_wire_5535)
    );

    bfr new_Jinkela_buffer_3085 (
        .din(new_Jinkela_wire_3514),
        .dout(new_Jinkela_wire_3515)
    );

    bfr new_Jinkela_buffer_3019 (
        .din(new_Jinkela_wire_3448),
        .dout(new_Jinkela_wire_3449)
    );

    bfr new_Jinkela_buffer_8333 (
        .din(new_Jinkela_wire_10472),
        .dout(new_Jinkela_wire_10473)
    );

    bfr new_Jinkela_buffer_4691 (
        .din(new_Jinkela_wire_5596),
        .dout(new_Jinkela_wire_5597)
    );

    bfr new_Jinkela_buffer_2959 (
        .din(new_Jinkela_wire_3386),
        .dout(new_Jinkela_wire_3387)
    );

    bfr new_Jinkela_buffer_4687 (
        .din(new_Jinkela_wire_5585),
        .dout(new_Jinkela_wire_5586)
    );

    bfr new_Jinkela_buffer_8358 (
        .din(new_Jinkela_wire_10497),
        .dout(new_Jinkela_wire_10498)
    );

    bfr new_Jinkela_buffer_4655 (
        .din(new_Jinkela_wire_5535),
        .dout(new_Jinkela_wire_5536)
    );

    bfr new_Jinkela_buffer_8334 (
        .din(new_Jinkela_wire_10473),
        .dout(new_Jinkela_wire_10474)
    );

    bfr new_Jinkela_buffer_2960 (
        .din(new_Jinkela_wire_3387),
        .dout(new_Jinkela_wire_3388)
    );

    spl2 new_Jinkela_splitter_869 (
        .a(n_1359_),
        .b(new_Jinkela_wire_10564),
        .c(new_Jinkela_wire_10565)
    );

    bfr new_Jinkela_buffer_4656 (
        .din(new_Jinkela_wire_5536),
        .dout(new_Jinkela_wire_5537)
    );

    bfr new_Jinkela_buffer_3083 (
        .din(new_Jinkela_wire_3512),
        .dout(new_Jinkela_wire_3513)
    );

    bfr new_Jinkela_buffer_3020 (
        .din(new_Jinkela_wire_3449),
        .dout(new_Jinkela_wire_3450)
    );

    bfr new_Jinkela_buffer_8335 (
        .din(new_Jinkela_wire_10474),
        .dout(new_Jinkela_wire_10475)
    );

    spl2 new_Jinkela_splitter_354 (
        .a(n_1317_),
        .b(new_Jinkela_wire_5731),
        .c(new_Jinkela_wire_5732)
    );

    bfr new_Jinkela_buffer_2961 (
        .din(new_Jinkela_wire_3388),
        .dout(new_Jinkela_wire_3389)
    );

    bfr new_Jinkela_buffer_4688 (
        .din(new_Jinkela_wire_5586),
        .dout(new_Jinkela_wire_5587)
    );

    bfr new_Jinkela_buffer_8359 (
        .din(new_Jinkela_wire_10498),
        .dout(new_Jinkela_wire_10499)
    );

    bfr new_Jinkela_buffer_4657 (
        .din(new_Jinkela_wire_5537),
        .dout(new_Jinkela_wire_5538)
    );

    bfr new_Jinkela_buffer_8336 (
        .din(new_Jinkela_wire_10475),
        .dout(new_Jinkela_wire_10476)
    );

    bfr new_Jinkela_buffer_2962 (
        .din(new_Jinkela_wire_3389),
        .dout(new_Jinkela_wire_3390)
    );

    spl2 new_Jinkela_splitter_348 (
        .a(n_0049_),
        .b(new_Jinkela_wire_5643),
        .c(new_Jinkela_wire_5644)
    );

    bfr new_Jinkela_buffer_8365 (
        .din(new_Jinkela_wire_10510),
        .dout(new_Jinkela_wire_10511)
    );

    bfr new_Jinkela_buffer_4658 (
        .din(new_Jinkela_wire_5538),
        .dout(new_Jinkela_wire_5539)
    );

    bfr new_Jinkela_buffer_3021 (
        .din(new_Jinkela_wire_3450),
        .dout(new_Jinkela_wire_3451)
    );

    bfr new_Jinkela_buffer_8337 (
        .din(new_Jinkela_wire_10476),
        .dout(new_Jinkela_wire_10477)
    );

    bfr new_Jinkela_buffer_4692 (
        .din(new_Jinkela_wire_5597),
        .dout(new_Jinkela_wire_5598)
    );

    bfr new_Jinkela_buffer_2963 (
        .din(new_Jinkela_wire_3390),
        .dout(new_Jinkela_wire_3391)
    );

    bfr new_Jinkela_buffer_8360 (
        .din(new_Jinkela_wire_10499),
        .dout(new_Jinkela_wire_10500)
    );

    bfr new_Jinkela_buffer_4659 (
        .din(new_Jinkela_wire_5539),
        .dout(new_Jinkela_wire_5540)
    );

    bfr new_Jinkela_buffer_3088 (
        .din(new_Jinkela_wire_3521),
        .dout(new_Jinkela_wire_3522)
    );

    bfr new_Jinkela_buffer_8338 (
        .din(new_Jinkela_wire_10477),
        .dout(new_Jinkela_wire_10478)
    );

    bfr new_Jinkela_buffer_2964 (
        .din(new_Jinkela_wire_3391),
        .dout(new_Jinkela_wire_3392)
    );

    bfr new_Jinkela_buffer_4727 (
        .din(new_net_2547),
        .dout(new_Jinkela_wire_5647)
    );

    bfr new_Jinkela_buffer_8379 (
        .din(new_Jinkela_wire_10532),
        .dout(new_Jinkela_wire_10533)
    );

    bfr new_Jinkela_buffer_4660 (
        .din(new_Jinkela_wire_5540),
        .dout(new_Jinkela_wire_5541)
    );

    bfr new_Jinkela_buffer_3086 (
        .din(new_Jinkela_wire_3515),
        .dout(new_Jinkela_wire_3516)
    );

    bfr new_Jinkela_buffer_3022 (
        .din(new_Jinkela_wire_3451),
        .dout(new_Jinkela_wire_3452)
    );

    bfr new_Jinkela_buffer_8339 (
        .din(new_Jinkela_wire_10478),
        .dout(new_Jinkela_wire_10479)
    );

    bfr new_Jinkela_buffer_4693 (
        .din(new_Jinkela_wire_5598),
        .dout(new_Jinkela_wire_5599)
    );

    bfr new_Jinkela_buffer_2965 (
        .din(new_Jinkela_wire_3392),
        .dout(new_Jinkela_wire_3393)
    );

    bfr new_Jinkela_buffer_8361 (
        .din(new_Jinkela_wire_10500),
        .dout(new_Jinkela_wire_10501)
    );

    bfr new_Jinkela_buffer_4661 (
        .din(new_Jinkela_wire_5541),
        .dout(new_Jinkela_wire_5542)
    );

    bfr new_Jinkela_buffer_8340 (
        .din(new_Jinkela_wire_10479),
        .dout(new_Jinkela_wire_10480)
    );

    bfr new_Jinkela_buffer_2966 (
        .din(new_Jinkela_wire_3393),
        .dout(new_Jinkela_wire_3394)
    );

    spl2 new_Jinkela_splitter_349 (
        .a(n_0009_),
        .b(new_Jinkela_wire_5645),
        .c(new_Jinkela_wire_5646)
    );

    bfr new_Jinkela_buffer_8366 (
        .din(new_Jinkela_wire_10511),
        .dout(new_Jinkela_wire_10512)
    );

    bfr new_Jinkela_buffer_4662 (
        .din(new_Jinkela_wire_5542),
        .dout(new_Jinkela_wire_5543)
    );

    bfr new_Jinkela_buffer_3023 (
        .din(new_Jinkela_wire_3452),
        .dout(new_Jinkela_wire_3453)
    );

    bfr new_Jinkela_buffer_8341 (
        .din(new_Jinkela_wire_10480),
        .dout(new_Jinkela_wire_10481)
    );

    bfr new_Jinkela_buffer_4694 (
        .din(new_Jinkela_wire_5599),
        .dout(new_Jinkela_wire_5600)
    );

    bfr new_Jinkela_buffer_2967 (
        .din(new_Jinkela_wire_3394),
        .dout(new_Jinkela_wire_3395)
    );

    bfr new_Jinkela_buffer_8401 (
        .din(new_Jinkela_wire_10566),
        .dout(new_Jinkela_wire_10567)
    );

    bfr new_Jinkela_buffer_4663 (
        .din(new_Jinkela_wire_5543),
        .dout(new_Jinkela_wire_5544)
    );

    bfr new_Jinkela_buffer_8342 (
        .din(new_Jinkela_wire_10481),
        .dout(new_Jinkela_wire_10482)
    );

    bfr new_Jinkela_buffer_4728 (
        .din(new_Jinkela_wire_5647),
        .dout(new_Jinkela_wire_5648)
    );

    bfr new_Jinkela_buffer_2968 (
        .din(new_Jinkela_wire_3395),
        .dout(new_Jinkela_wire_3396)
    );

    bfr new_Jinkela_buffer_8367 (
        .din(new_Jinkela_wire_10512),
        .dout(new_Jinkela_wire_10513)
    );

    bfr new_Jinkela_buffer_4664 (
        .din(new_Jinkela_wire_5544),
        .dout(new_Jinkela_wire_5545)
    );

    bfr new_Jinkela_buffer_3087 (
        .din(new_Jinkela_wire_3516),
        .dout(new_Jinkela_wire_3517)
    );

    bfr new_Jinkela_buffer_3024 (
        .din(new_Jinkela_wire_3453),
        .dout(new_Jinkela_wire_3454)
    );

    bfr new_Jinkela_buffer_8343 (
        .din(new_Jinkela_wire_10482),
        .dout(new_Jinkela_wire_10483)
    );

    bfr new_Jinkela_buffer_4695 (
        .din(new_Jinkela_wire_5600),
        .dout(new_Jinkela_wire_5601)
    );

    bfr new_Jinkela_buffer_2969 (
        .din(new_Jinkela_wire_3396),
        .dout(new_Jinkela_wire_3397)
    );

    bfr new_Jinkela_buffer_8380 (
        .din(new_Jinkela_wire_10533),
        .dout(new_Jinkela_wire_10534)
    );

    bfr new_Jinkela_buffer_4665 (
        .din(new_Jinkela_wire_5545),
        .dout(new_Jinkela_wire_5546)
    );

    bfr new_Jinkela_buffer_8344 (
        .din(new_Jinkela_wire_10483),
        .dout(new_Jinkela_wire_10484)
    );

    spl2 new_Jinkela_splitter_350 (
        .a(n_0121_),
        .b(new_Jinkela_wire_5676),
        .c(new_Jinkela_wire_5677)
    );

    bfr new_Jinkela_buffer_2970 (
        .din(new_Jinkela_wire_3397),
        .dout(new_Jinkela_wire_3398)
    );

    bfr new_Jinkela_buffer_8368 (
        .din(new_Jinkela_wire_10513),
        .dout(new_Jinkela_wire_10514)
    );

    bfr new_Jinkela_buffer_4666 (
        .din(new_Jinkela_wire_5546),
        .dout(new_Jinkela_wire_5547)
    );

    bfr new_Jinkela_buffer_3091 (
        .din(new_Jinkela_wire_3524),
        .dout(new_Jinkela_wire_3525)
    );

    bfr new_Jinkela_buffer_3025 (
        .din(new_Jinkela_wire_3454),
        .dout(new_Jinkela_wire_3455)
    );

    bfr new_Jinkela_buffer_4696 (
        .din(new_Jinkela_wire_5601),
        .dout(new_Jinkela_wire_5602)
    );

    bfr new_Jinkela_buffer_2971 (
        .din(new_Jinkela_wire_3398),
        .dout(new_Jinkela_wire_3399)
    );

    spl2 new_Jinkela_splitter_867 (
        .a(new_Jinkela_wire_10558),
        .b(new_Jinkela_wire_10559),
        .c(new_Jinkela_wire_10560)
    );

    bfr new_Jinkela_buffer_8369 (
        .din(new_Jinkela_wire_10514),
        .dout(new_Jinkela_wire_10515)
    );

    bfr new_Jinkela_buffer_4667 (
        .din(new_Jinkela_wire_5547),
        .dout(new_Jinkela_wire_5548)
    );

    bfr new_Jinkela_buffer_3094 (
        .din(N169),
        .dout(new_Jinkela_wire_3528)
    );

    bfr new_Jinkela_buffer_8381 (
        .din(new_Jinkela_wire_10534),
        .dout(new_Jinkela_wire_10535)
    );

    bfr new_Jinkela_buffer_2972 (
        .din(new_Jinkela_wire_3399),
        .dout(new_Jinkela_wire_3400)
    );

    bfr new_Jinkela_buffer_8370 (
        .din(new_Jinkela_wire_10515),
        .dout(new_Jinkela_wire_10516)
    );

    bfr new_Jinkela_buffer_4668 (
        .din(new_Jinkela_wire_5548),
        .dout(new_Jinkela_wire_5549)
    );

    bfr new_Jinkela_buffer_3026 (
        .din(new_Jinkela_wire_3455),
        .dout(new_Jinkela_wire_3456)
    );

    bfr new_Jinkela_buffer_4697 (
        .din(new_Jinkela_wire_5602),
        .dout(new_Jinkela_wire_5603)
    );

    bfr new_Jinkela_buffer_2973 (
        .din(new_Jinkela_wire_3400),
        .dout(new_Jinkela_wire_3401)
    );

    bfr new_Jinkela_buffer_8371 (
        .din(new_Jinkela_wire_10516),
        .dout(new_Jinkela_wire_10517)
    );

    bfr new_Jinkela_buffer_4669 (
        .din(new_Jinkela_wire_5549),
        .dout(new_Jinkela_wire_5550)
    );

    bfr new_Jinkela_buffer_3089 (
        .din(new_Jinkela_wire_3522),
        .dout(new_Jinkela_wire_3523)
    );

    bfr new_Jinkela_buffer_8382 (
        .din(new_Jinkela_wire_10535),
        .dout(new_Jinkela_wire_10536)
    );

    bfr new_Jinkela_buffer_4729 (
        .din(new_Jinkela_wire_5648),
        .dout(new_Jinkela_wire_5649)
    );

    bfr new_Jinkela_buffer_2974 (
        .din(new_Jinkela_wire_3401),
        .dout(new_Jinkela_wire_3402)
    );

    bfr new_Jinkela_buffer_8372 (
        .din(new_Jinkela_wire_10517),
        .dout(new_Jinkela_wire_10518)
    );

    bfr new_Jinkela_buffer_4670 (
        .din(new_Jinkela_wire_5550),
        .dout(new_Jinkela_wire_5551)
    );

    bfr new_Jinkela_buffer_3027 (
        .din(new_Jinkela_wire_3456),
        .dout(new_Jinkela_wire_3457)
    );

    spl2 new_Jinkela_splitter_871 (
        .a(n_0728_),
        .b(new_Jinkela_wire_10629),
        .c(new_Jinkela_wire_10630)
    );

    bfr new_Jinkela_buffer_4698 (
        .din(new_Jinkela_wire_5603),
        .dout(new_Jinkela_wire_5604)
    );

    bfr new_Jinkela_buffer_2975 (
        .din(new_Jinkela_wire_3402),
        .dout(new_Jinkela_wire_3403)
    );

    bfr new_Jinkela_buffer_8373 (
        .din(new_Jinkela_wire_10518),
        .dout(new_Jinkela_wire_10519)
    );

    bfr new_Jinkela_buffer_4671 (
        .din(new_Jinkela_wire_5551),
        .dout(new_Jinkela_wire_5552)
    );

    bfr new_Jinkela_buffer_8383 (
        .din(new_Jinkela_wire_10536),
        .dout(new_Jinkela_wire_10537)
    );

    spl3L new_Jinkela_splitter_355 (
        .a(n_0112_),
        .d(new_Jinkela_wire_5755),
        .b(new_Jinkela_wire_5756),
        .c(new_Jinkela_wire_5757)
    );

    bfr new_Jinkela_buffer_2976 (
        .din(new_Jinkela_wire_3403),
        .dout(new_Jinkela_wire_3404)
    );

    bfr new_Jinkela_buffer_4800 (
        .din(n_0318_),
        .dout(new_Jinkela_wire_5730)
    );

    bfr new_Jinkela_buffer_8374 (
        .din(new_Jinkela_wire_10519),
        .dout(new_Jinkela_wire_10520)
    );

    bfr new_Jinkela_buffer_4672 (
        .din(new_Jinkela_wire_5552),
        .dout(new_Jinkela_wire_5553)
    );

    bfr new_Jinkela_buffer_3098 (
        .din(N35),
        .dout(new_Jinkela_wire_3532)
    );

    bfr new_Jinkela_buffer_3028 (
        .din(new_Jinkela_wire_3457),
        .dout(new_Jinkela_wire_3458)
    );

    bfr new_Jinkela_buffer_8400 (
        .din(n_0163_),
        .dout(new_Jinkela_wire_10566)
    );

    bfr new_Jinkela_buffer_4699 (
        .din(new_Jinkela_wire_5604),
        .dout(new_Jinkela_wire_5605)
    );

    bfr new_Jinkela_buffer_2977 (
        .din(new_Jinkela_wire_3404),
        .dout(new_Jinkela_wire_3405)
    );

    bfr new_Jinkela_buffer_8375 (
        .din(new_Jinkela_wire_10520),
        .dout(new_Jinkela_wire_10521)
    );

    bfr new_Jinkela_buffer_4730 (
        .din(new_Jinkela_wire_5649),
        .dout(new_Jinkela_wire_5650)
    );

    bfr new_Jinkela_buffer_8384 (
        .din(new_Jinkela_wire_10537),
        .dout(new_Jinkela_wire_10538)
    );

    bfr new_Jinkela_buffer_4700 (
        .din(new_Jinkela_wire_5605),
        .dout(new_Jinkela_wire_5606)
    );

    bfr new_Jinkela_buffer_2978 (
        .din(new_Jinkela_wire_3405),
        .dout(new_Jinkela_wire_3406)
    );

    bfr new_Jinkela_buffer_785 (
        .din(new_Jinkela_wire_845),
        .dout(new_Jinkela_wire_846)
    );

    bfr new_Jinkela_buffer_833 (
        .din(new_Jinkela_wire_898),
        .dout(new_Jinkela_wire_899)
    );

    bfr new_Jinkela_buffer_7213 (
        .din(n_0669_),
        .dout(new_Jinkela_wire_8934)
    );

    bfr new_Jinkela_buffer_7182 (
        .din(new_Jinkela_wire_8895),
        .dout(new_Jinkela_wire_8896)
    );

    bfr new_Jinkela_buffer_786 (
        .din(new_Jinkela_wire_846),
        .dout(new_Jinkela_wire_847)
    );

    bfr new_Jinkela_buffer_889 (
        .din(new_Jinkela_wire_959),
        .dout(new_Jinkela_wire_960)
    );

    bfr new_Jinkela_buffer_7183 (
        .din(new_Jinkela_wire_8896),
        .dout(new_Jinkela_wire_8897)
    );

    bfr new_Jinkela_buffer_787 (
        .din(new_Jinkela_wire_847),
        .dout(new_Jinkela_wire_848)
    );

    spl3L new_Jinkela_splitter_692 (
        .a(n_0152_),
        .d(new_Jinkela_wire_8942),
        .b(new_Jinkela_wire_8943),
        .c(new_Jinkela_wire_8944)
    );

    bfr new_Jinkela_buffer_834 (
        .din(new_Jinkela_wire_899),
        .dout(new_Jinkela_wire_900)
    );

    spl3L new_Jinkela_splitter_688 (
        .a(new_Jinkela_wire_8927),
        .d(new_Jinkela_wire_8928),
        .b(new_Jinkela_wire_8929),
        .c(new_Jinkela_wire_8930)
    );

    bfr new_Jinkela_buffer_7184 (
        .din(new_Jinkela_wire_8897),
        .dout(new_Jinkela_wire_8898)
    );

    bfr new_Jinkela_buffer_788 (
        .din(new_Jinkela_wire_848),
        .dout(new_Jinkela_wire_849)
    );

    spl3L new_Jinkela_splitter_690 (
        .a(n_0692_),
        .d(new_Jinkela_wire_8936),
        .b(new_Jinkela_wire_8937),
        .c(new_Jinkela_wire_8938)
    );

    bfr new_Jinkela_buffer_1013 (
        .din(new_Jinkela_wire_1087),
        .dout(new_Jinkela_wire_1088)
    );

    bfr new_Jinkela_buffer_7212 (
        .din(new_Jinkela_wire_8930),
        .dout(new_Jinkela_wire_8931)
    );

    bfr new_Jinkela_buffer_7185 (
        .din(new_Jinkela_wire_8898),
        .dout(new_Jinkela_wire_8899)
    );

    bfr new_Jinkela_buffer_789 (
        .din(new_Jinkela_wire_849),
        .dout(new_Jinkela_wire_850)
    );

    bfr new_Jinkela_buffer_835 (
        .din(new_Jinkela_wire_900),
        .dout(new_Jinkela_wire_901)
    );

    bfr new_Jinkela_buffer_7214 (
        .din(n_0698_),
        .dout(new_Jinkela_wire_8935)
    );

    bfr new_Jinkela_buffer_7186 (
        .din(new_Jinkela_wire_8899),
        .dout(new_Jinkela_wire_8900)
    );

    bfr new_Jinkela_buffer_790 (
        .din(new_Jinkela_wire_850),
        .dout(new_Jinkela_wire_851)
    );

    spl2 new_Jinkela_splitter_693 (
        .a(n_1224_),
        .b(new_Jinkela_wire_8946),
        .c(new_Jinkela_wire_8947)
    );

    bfr new_Jinkela_buffer_890 (
        .din(new_Jinkela_wire_960),
        .dout(new_Jinkela_wire_961)
    );

    bfr new_Jinkela_buffer_7216 (
        .din(n_0499_),
        .dout(new_Jinkela_wire_8945)
    );

    bfr new_Jinkela_buffer_7187 (
        .din(new_Jinkela_wire_8900),
        .dout(new_Jinkela_wire_8901)
    );

    bfr new_Jinkela_buffer_791 (
        .din(new_Jinkela_wire_851),
        .dout(new_Jinkela_wire_852)
    );

    spl2 new_Jinkela_splitter_689 (
        .a(new_Jinkela_wire_8931),
        .b(new_Jinkela_wire_8932),
        .c(new_Jinkela_wire_8933)
    );

    bfr new_Jinkela_buffer_836 (
        .din(new_Jinkela_wire_901),
        .dout(new_Jinkela_wire_902)
    );

    bfr new_Jinkela_buffer_7188 (
        .din(new_Jinkela_wire_8901),
        .dout(new_Jinkela_wire_8902)
    );

    bfr new_Jinkela_buffer_792 (
        .din(new_Jinkela_wire_852),
        .dout(new_Jinkela_wire_853)
    );

    bfr new_Jinkela_buffer_7215 (
        .din(new_Jinkela_wire_8938),
        .dout(new_Jinkela_wire_8939)
    );

    bfr new_Jinkela_buffer_1016 (
        .din(new_Jinkela_wire_1090),
        .dout(new_Jinkela_wire_1091)
    );

    bfr new_Jinkela_buffer_7217 (
        .din(new_net_2511),
        .dout(new_Jinkela_wire_8948)
    );

    bfr new_Jinkela_buffer_7189 (
        .din(new_Jinkela_wire_8902),
        .dout(new_Jinkela_wire_8903)
    );

    bfr new_Jinkela_buffer_793 (
        .din(new_Jinkela_wire_853),
        .dout(new_Jinkela_wire_854)
    );

    bfr new_Jinkela_buffer_837 (
        .din(new_Jinkela_wire_902),
        .dout(new_Jinkela_wire_903)
    );

    bfr new_Jinkela_buffer_7190 (
        .din(new_Jinkela_wire_8903),
        .dout(new_Jinkela_wire_8904)
    );

    bfr new_Jinkela_buffer_794 (
        .din(new_Jinkela_wire_854),
        .dout(new_Jinkela_wire_855)
    );

    bfr new_Jinkela_buffer_7218 (
        .din(new_Jinkela_wire_8948),
        .dout(new_Jinkela_wire_8949)
    );

    bfr new_Jinkela_buffer_891 (
        .din(new_Jinkela_wire_961),
        .dout(new_Jinkela_wire_962)
    );

    bfr new_Jinkela_buffer_7191 (
        .din(new_Jinkela_wire_8904),
        .dout(new_Jinkela_wire_8905)
    );

    bfr new_Jinkela_buffer_795 (
        .din(new_Jinkela_wire_855),
        .dout(new_Jinkela_wire_856)
    );

    spl2 new_Jinkela_splitter_691 (
        .a(new_Jinkela_wire_8939),
        .b(new_Jinkela_wire_8940),
        .c(new_Jinkela_wire_8941)
    );

    bfr new_Jinkela_buffer_838 (
        .din(new_Jinkela_wire_903),
        .dout(new_Jinkela_wire_904)
    );

    bfr new_Jinkela_buffer_7192 (
        .din(new_Jinkela_wire_8905),
        .dout(new_Jinkela_wire_8906)
    );

    bfr new_Jinkela_buffer_796 (
        .din(new_Jinkela_wire_856),
        .dout(new_Jinkela_wire_857)
    );

    bfr new_Jinkela_buffer_950 (
        .din(new_Jinkela_wire_1024),
        .dout(new_Jinkela_wire_1025)
    );

    bfr new_Jinkela_buffer_7193 (
        .din(new_Jinkela_wire_8906),
        .dout(new_Jinkela_wire_8907)
    );

    bfr new_Jinkela_buffer_797 (
        .din(new_Jinkela_wire_857),
        .dout(new_Jinkela_wire_858)
    );

    bfr new_Jinkela_buffer_839 (
        .din(new_Jinkela_wire_904),
        .dout(new_Jinkela_wire_905)
    );

    bfr new_Jinkela_buffer_7194 (
        .din(new_Jinkela_wire_8907),
        .dout(new_Jinkela_wire_8908)
    );

    bfr new_Jinkela_buffer_798 (
        .din(new_Jinkela_wire_858),
        .dout(new_Jinkela_wire_859)
    );

    bfr new_Jinkela_buffer_7247 (
        .din(n_0427_),
        .dout(new_Jinkela_wire_8978)
    );

    bfr new_Jinkela_buffer_892 (
        .din(new_Jinkela_wire_962),
        .dout(new_Jinkela_wire_963)
    );

    bfr new_Jinkela_buffer_7195 (
        .din(new_Jinkela_wire_8908),
        .dout(new_Jinkela_wire_8909)
    );

    bfr new_Jinkela_buffer_799 (
        .din(new_Jinkela_wire_859),
        .dout(new_Jinkela_wire_860)
    );

    bfr new_Jinkela_buffer_7264 (
        .din(n_0254_),
        .dout(new_Jinkela_wire_8995)
    );

    bfr new_Jinkela_buffer_840 (
        .din(new_Jinkela_wire_905),
        .dout(new_Jinkela_wire_906)
    );

    bfr new_Jinkela_buffer_7196 (
        .din(new_Jinkela_wire_8909),
        .dout(new_Jinkela_wire_8910)
    );

    bfr new_Jinkela_buffer_800 (
        .din(new_Jinkela_wire_860),
        .dout(new_Jinkela_wire_861)
    );

    bfr new_Jinkela_buffer_7219 (
        .din(new_Jinkela_wire_8949),
        .dout(new_Jinkela_wire_8950)
    );

    bfr new_Jinkela_buffer_1014 (
        .din(new_Jinkela_wire_1088),
        .dout(new_Jinkela_wire_1089)
    );

    bfr new_Jinkela_buffer_7197 (
        .din(new_Jinkela_wire_8910),
        .dout(new_Jinkela_wire_8911)
    );

    bfr new_Jinkela_buffer_801 (
        .din(new_Jinkela_wire_861),
        .dout(new_Jinkela_wire_862)
    );

    bfr new_Jinkela_buffer_7248 (
        .din(new_Jinkela_wire_8978),
        .dout(new_Jinkela_wire_8979)
    );

    bfr new_Jinkela_buffer_841 (
        .din(new_Jinkela_wire_906),
        .dout(new_Jinkela_wire_907)
    );

    bfr new_Jinkela_buffer_7198 (
        .din(new_Jinkela_wire_8911),
        .dout(new_Jinkela_wire_8912)
    );

    bfr new_Jinkela_buffer_802 (
        .din(new_Jinkela_wire_862),
        .dout(new_Jinkela_wire_863)
    );

    bfr new_Jinkela_buffer_7220 (
        .din(new_Jinkela_wire_8950),
        .dout(new_Jinkela_wire_8951)
    );

    bfr new_Jinkela_buffer_893 (
        .din(new_Jinkela_wire_963),
        .dout(new_Jinkela_wire_964)
    );

    bfr new_Jinkela_buffer_7199 (
        .din(new_Jinkela_wire_8912),
        .dout(new_Jinkela_wire_8913)
    );

    bfr new_Jinkela_buffer_803 (
        .din(new_Jinkela_wire_863),
        .dout(new_Jinkela_wire_864)
    );

    spl2 new_Jinkela_splitter_694 (
        .a(n_0842_),
        .b(new_Jinkela_wire_8996),
        .c(new_Jinkela_wire_8997)
    );

    bfr new_Jinkela_buffer_842 (
        .din(new_Jinkela_wire_907),
        .dout(new_Jinkela_wire_908)
    );

    spl2 new_Jinkela_splitter_695 (
        .a(n_0847_),
        .b(new_Jinkela_wire_8998),
        .c(new_Jinkela_wire_8999)
    );

    bfr new_Jinkela_buffer_7200 (
        .din(new_Jinkela_wire_8913),
        .dout(new_Jinkela_wire_8914)
    );

    bfr new_Jinkela_buffer_804 (
        .din(new_Jinkela_wire_864),
        .dout(new_Jinkela_wire_865)
    );

    bfr new_Jinkela_buffer_7221 (
        .din(new_Jinkela_wire_8951),
        .dout(new_Jinkela_wire_8952)
    );

    bfr new_Jinkela_buffer_951 (
        .din(new_Jinkela_wire_1025),
        .dout(new_Jinkela_wire_1026)
    );

    bfr new_Jinkela_buffer_7201 (
        .din(new_Jinkela_wire_8914),
        .dout(new_Jinkela_wire_8915)
    );

    bfr new_Jinkela_buffer_805 (
        .din(new_Jinkela_wire_865),
        .dout(new_Jinkela_wire_866)
    );

    bfr new_Jinkela_buffer_7249 (
        .din(new_Jinkela_wire_8979),
        .dout(new_Jinkela_wire_8980)
    );

    bfr new_Jinkela_buffer_843 (
        .din(new_Jinkela_wire_908),
        .dout(new_Jinkela_wire_909)
    );

    bfr new_Jinkela_buffer_7202 (
        .din(new_Jinkela_wire_8915),
        .dout(new_Jinkela_wire_8916)
    );

    bfr new_Jinkela_buffer_3836 (
        .din(new_Jinkela_wire_4469),
        .dout(new_Jinkela_wire_4470)
    );

    bfr new_Jinkela_buffer_2066 (
        .din(new_Jinkela_wire_2435),
        .dout(new_Jinkela_wire_2436)
    );

    bfr new_Jinkela_buffer_6360 (
        .din(new_Jinkela_wire_7759),
        .dout(new_Jinkela_wire_7760)
    );

    bfr new_Jinkela_buffer_6333 (
        .din(new_Jinkela_wire_7714),
        .dout(new_Jinkela_wire_7715)
    );

    bfr new_Jinkela_buffer_2202 (
        .din(new_Jinkela_wire_2582),
        .dout(new_Jinkela_wire_2583)
    );

    bfr new_Jinkela_buffer_3864 (
        .din(new_Jinkela_wire_4499),
        .dout(new_Jinkela_wire_4500)
    );

    bfr new_Jinkela_buffer_3837 (
        .din(new_Jinkela_wire_4470),
        .dout(new_Jinkela_wire_4471)
    );

    bfr new_Jinkela_buffer_2067 (
        .din(new_Jinkela_wire_2436),
        .dout(new_Jinkela_wire_2437)
    );

    bfr new_Jinkela_buffer_6334 (
        .din(new_Jinkela_wire_7715),
        .dout(new_Jinkela_wire_7716)
    );

    bfr new_Jinkela_buffer_2119 (
        .din(new_Jinkela_wire_2493),
        .dout(new_Jinkela_wire_2494)
    );

    bfr new_Jinkela_buffer_6366 (
        .din(new_Jinkela_wire_7769),
        .dout(new_Jinkela_wire_7770)
    );

    bfr new_Jinkela_buffer_3838 (
        .din(new_Jinkela_wire_4471),
        .dout(new_Jinkela_wire_4472)
    );

    bfr new_Jinkela_buffer_2068 (
        .din(new_Jinkela_wire_2437),
        .dout(new_Jinkela_wire_2438)
    );

    bfr new_Jinkela_buffer_6361 (
        .din(new_Jinkela_wire_7760),
        .dout(new_Jinkela_wire_7761)
    );

    bfr new_Jinkela_buffer_6335 (
        .din(new_Jinkela_wire_7716),
        .dout(new_Jinkela_wire_7717)
    );

    bfr new_Jinkela_buffer_3872 (
        .din(new_Jinkela_wire_4524),
        .dout(new_Jinkela_wire_4525)
    );

    bfr new_Jinkela_buffer_2182 (
        .din(new_Jinkela_wire_2558),
        .dout(new_Jinkela_wire_2559)
    );

    bfr new_Jinkela_buffer_3865 (
        .din(new_Jinkela_wire_4500),
        .dout(new_Jinkela_wire_4501)
    );

    bfr new_Jinkela_buffer_3839 (
        .din(new_Jinkela_wire_4472),
        .dout(new_Jinkela_wire_4473)
    );

    bfr new_Jinkela_buffer_2069 (
        .din(new_Jinkela_wire_2438),
        .dout(new_Jinkela_wire_2439)
    );

    bfr new_Jinkela_buffer_6336 (
        .din(new_Jinkela_wire_7717),
        .dout(new_Jinkela_wire_7718)
    );

    bfr new_Jinkela_buffer_2120 (
        .din(new_Jinkela_wire_2494),
        .dout(new_Jinkela_wire_2495)
    );

    bfr new_Jinkela_buffer_3840 (
        .din(new_Jinkela_wire_4473),
        .dout(new_Jinkela_wire_4474)
    );

    bfr new_Jinkela_buffer_2070 (
        .din(new_Jinkela_wire_2439),
        .dout(new_Jinkela_wire_2440)
    );

    bfr new_Jinkela_buffer_6362 (
        .din(new_Jinkela_wire_7761),
        .dout(new_Jinkela_wire_7762)
    );

    bfr new_Jinkela_buffer_6337 (
        .din(new_Jinkela_wire_7718),
        .dout(new_Jinkela_wire_7719)
    );

    spl2 new_Jinkela_splitter_237 (
        .a(n_0769_),
        .b(new_Jinkela_wire_4527),
        .c(new_Jinkela_wire_4528)
    );

    bfr new_Jinkela_buffer_2205 (
        .din(new_Jinkela_wire_2587),
        .dout(new_Jinkela_wire_2588)
    );

    spl3L new_Jinkela_splitter_238 (
        .a(n_0074_),
        .d(new_Jinkela_wire_4529),
        .b(new_Jinkela_wire_4530),
        .c(new_Jinkela_wire_4531)
    );

    bfr new_Jinkela_buffer_3841 (
        .din(new_Jinkela_wire_4474),
        .dout(new_Jinkela_wire_4475)
    );

    bfr new_Jinkela_buffer_2071 (
        .din(new_Jinkela_wire_2440),
        .dout(new_Jinkela_wire_2441)
    );

    spl2 new_Jinkela_splitter_557 (
        .a(n_0939_),
        .b(new_Jinkela_wire_7824),
        .c(new_Jinkela_wire_7825)
    );

    bfr new_Jinkela_buffer_6338 (
        .din(new_Jinkela_wire_7719),
        .dout(new_Jinkela_wire_7720)
    );

    spl2 new_Jinkela_splitter_240 (
        .a(n_0868_),
        .b(new_Jinkela_wire_4534),
        .c(new_Jinkela_wire_4535)
    );

    bfr new_Jinkela_buffer_2121 (
        .din(new_Jinkela_wire_2495),
        .dout(new_Jinkela_wire_2496)
    );

    spl2 new_Jinkela_splitter_242 (
        .a(n_0809_),
        .b(new_Jinkela_wire_4539),
        .c(new_Jinkela_wire_4540)
    );

    bfr new_Jinkela_buffer_6367 (
        .din(new_Jinkela_wire_7770),
        .dout(new_Jinkela_wire_7771)
    );

    bfr new_Jinkela_buffer_3842 (
        .din(new_Jinkela_wire_4475),
        .dout(new_Jinkela_wire_4476)
    );

    bfr new_Jinkela_buffer_2072 (
        .din(new_Jinkela_wire_2441),
        .dout(new_Jinkela_wire_2442)
    );

    bfr new_Jinkela_buffer_6363 (
        .din(new_Jinkela_wire_7762),
        .dout(new_Jinkela_wire_7763)
    );

    bfr new_Jinkela_buffer_6339 (
        .din(new_Jinkela_wire_7720),
        .dout(new_Jinkela_wire_7721)
    );

    bfr new_Jinkela_buffer_2183 (
        .din(new_Jinkela_wire_2559),
        .dout(new_Jinkela_wire_2560)
    );

    bfr new_Jinkela_buffer_2204 (
        .din(new_Jinkela_wire_2584),
        .dout(new_Jinkela_wire_2585)
    );

    spl2 new_Jinkela_splitter_239 (
        .a(n_0442_),
        .b(new_Jinkela_wire_4532),
        .c(new_Jinkela_wire_4533)
    );

    bfr new_Jinkela_buffer_3843 (
        .din(new_Jinkela_wire_4476),
        .dout(new_Jinkela_wire_4477)
    );

    bfr new_Jinkela_buffer_2073 (
        .din(new_Jinkela_wire_2442),
        .dout(new_Jinkela_wire_2443)
    );

    bfr new_Jinkela_buffer_6340 (
        .din(new_Jinkela_wire_7721),
        .dout(new_Jinkela_wire_7722)
    );

    bfr new_Jinkela_buffer_2122 (
        .din(new_Jinkela_wire_2496),
        .dout(new_Jinkela_wire_2497)
    );

    bfr new_Jinkela_buffer_6369 (
        .din(new_Jinkela_wire_7774),
        .dout(new_Jinkela_wire_7775)
    );

    bfr new_Jinkela_buffer_3844 (
        .din(new_Jinkela_wire_4477),
        .dout(new_Jinkela_wire_4478)
    );

    bfr new_Jinkela_buffer_2074 (
        .din(new_Jinkela_wire_2443),
        .dout(new_Jinkela_wire_2444)
    );

    spl2 new_Jinkela_splitter_551 (
        .a(new_Jinkela_wire_7763),
        .b(new_Jinkela_wire_7764),
        .c(new_Jinkela_wire_7765)
    );

    bfr new_Jinkela_buffer_6341 (
        .din(new_Jinkela_wire_7722),
        .dout(new_Jinkela_wire_7723)
    );

    bfr new_Jinkela_buffer_2203 (
        .din(new_Jinkela_wire_2583),
        .dout(new_Jinkela_wire_2584)
    );

    bfr new_Jinkela_buffer_3845 (
        .din(new_Jinkela_wire_4478),
        .dout(new_Jinkela_wire_4479)
    );

    bfr new_Jinkela_buffer_2075 (
        .din(new_Jinkela_wire_2444),
        .dout(new_Jinkela_wire_2445)
    );

    bfr new_Jinkela_buffer_6400 (
        .din(new_Jinkela_wire_7807),
        .dout(new_Jinkela_wire_7808)
    );

    bfr new_Jinkela_buffer_6342 (
        .din(new_Jinkela_wire_7723),
        .dout(new_Jinkela_wire_7724)
    );

    spl3L new_Jinkela_splitter_241 (
        .a(n_0053_),
        .d(new_Jinkela_wire_4536),
        .b(new_Jinkela_wire_4537),
        .c(new_Jinkela_wire_4538)
    );

    bfr new_Jinkela_buffer_2123 (
        .din(new_Jinkela_wire_2497),
        .dout(new_Jinkela_wire_2498)
    );

    spl2 new_Jinkela_splitter_243 (
        .a(n_0488_),
        .b(new_Jinkela_wire_4541),
        .c(new_Jinkela_wire_4542)
    );

    bfr new_Jinkela_buffer_6370 (
        .din(new_Jinkela_wire_7775),
        .dout(new_Jinkela_wire_7776)
    );

    bfr new_Jinkela_buffer_3846 (
        .din(new_Jinkela_wire_4479),
        .dout(new_Jinkela_wire_4480)
    );

    bfr new_Jinkela_buffer_2076 (
        .din(new_Jinkela_wire_2445),
        .dout(new_Jinkela_wire_2446)
    );

    bfr new_Jinkela_buffer_6343 (
        .din(new_Jinkela_wire_7724),
        .dout(new_Jinkela_wire_7725)
    );

    bfr new_Jinkela_buffer_2184 (
        .din(new_Jinkela_wire_2560),
        .dout(new_Jinkela_wire_2561)
    );

    bfr new_Jinkela_buffer_6410 (
        .din(n_1143_),
        .dout(new_Jinkela_wire_7820)
    );

    bfr new_Jinkela_buffer_3847 (
        .din(new_Jinkela_wire_4480),
        .dout(new_Jinkela_wire_4481)
    );

    bfr new_Jinkela_buffer_2124 (
        .din(new_Jinkela_wire_2498),
        .dout(new_Jinkela_wire_2499)
    );

    spl2 new_Jinkela_splitter_544 (
        .a(new_Jinkela_wire_7725),
        .b(new_Jinkela_wire_7726),
        .c(new_Jinkela_wire_7727)
    );

    bfr new_Jinkela_buffer_2272 (
        .din(N233),
        .dout(new_Jinkela_wire_2659)
    );

    bfr new_Jinkela_buffer_6371 (
        .din(new_Jinkela_wire_7776),
        .dout(new_Jinkela_wire_7777)
    );

    bfr new_Jinkela_buffer_3848 (
        .din(new_Jinkela_wire_4481),
        .dout(new_Jinkela_wire_4482)
    );

    bfr new_Jinkela_buffer_2125 (
        .din(new_Jinkela_wire_2499),
        .dout(new_Jinkela_wire_2500)
    );

    bfr new_Jinkela_buffer_6399 (
        .din(new_Jinkela_wire_7806),
        .dout(new_Jinkela_wire_7807)
    );

    spl2 new_Jinkela_splitter_244 (
        .a(n_0244_),
        .b(new_Jinkela_wire_4543),
        .c(new_Jinkela_wire_4544)
    );

    bfr new_Jinkela_buffer_2185 (
        .din(new_Jinkela_wire_2561),
        .dout(new_Jinkela_wire_2562)
    );

    bfr new_Jinkela_buffer_3875 (
        .din(new_Jinkela_wire_4545),
        .dout(new_Jinkela_wire_4546)
    );

    bfr new_Jinkela_buffer_3849 (
        .din(new_Jinkela_wire_4482),
        .dout(new_Jinkela_wire_4483)
    );

    bfr new_Jinkela_buffer_2126 (
        .din(new_Jinkela_wire_2500),
        .dout(new_Jinkela_wire_2501)
    );

    bfr new_Jinkela_buffer_6415 (
        .din(n_1156_),
        .dout(new_Jinkela_wire_7829)
    );

    bfr new_Jinkela_buffer_6372 (
        .din(new_Jinkela_wire_7777),
        .dout(new_Jinkela_wire_7778)
    );

    bfr new_Jinkela_buffer_3874 (
        .din(new_net_2539),
        .dout(new_Jinkela_wire_4545)
    );

    bfr new_Jinkela_buffer_3850 (
        .din(new_Jinkela_wire_4483),
        .dout(new_Jinkela_wire_4484)
    );

    bfr new_Jinkela_buffer_2127 (
        .din(new_Jinkela_wire_2501),
        .dout(new_Jinkela_wire_2502)
    );

    bfr new_Jinkela_buffer_6373 (
        .din(new_Jinkela_wire_7778),
        .dout(new_Jinkela_wire_7779)
    );

    bfr new_Jinkela_buffer_3899 (
        .din(n_0165_),
        .dout(new_Jinkela_wire_4570)
    );

    bfr new_Jinkela_buffer_2186 (
        .din(new_Jinkela_wire_2562),
        .dout(new_Jinkela_wire_2563)
    );

    bfr new_Jinkela_buffer_6411 (
        .din(new_Jinkela_wire_7820),
        .dout(new_Jinkela_wire_7821)
    );

    bfr new_Jinkela_buffer_3851 (
        .din(new_Jinkela_wire_4484),
        .dout(new_Jinkela_wire_4485)
    );

    bfr new_Jinkela_buffer_2128 (
        .din(new_Jinkela_wire_2502),
        .dout(new_Jinkela_wire_2503)
    );

    bfr new_Jinkela_buffer_6374 (
        .din(new_Jinkela_wire_7779),
        .dout(new_Jinkela_wire_7780)
    );

    spl2 new_Jinkela_splitter_245 (
        .a(n_1099_),
        .b(new_Jinkela_wire_4627),
        .c(new_Jinkela_wire_4628)
    );

    bfr new_Jinkela_buffer_3956 (
        .din(n_0256_),
        .dout(new_Jinkela_wire_4629)
    );

    bfr new_Jinkela_buffer_6401 (
        .din(new_Jinkela_wire_7808),
        .dout(new_Jinkela_wire_7809)
    );

    bfr new_Jinkela_buffer_3876 (
        .din(new_Jinkela_wire_4546),
        .dout(new_Jinkela_wire_4547)
    );

    bfr new_Jinkela_buffer_2129 (
        .din(new_Jinkela_wire_2503),
        .dout(new_Jinkela_wire_2504)
    );

    bfr new_Jinkela_buffer_6375 (
        .din(new_Jinkela_wire_7780),
        .dout(new_Jinkela_wire_7781)
    );

    bfr new_Jinkela_buffer_3900 (
        .din(new_Jinkela_wire_4570),
        .dout(new_Jinkela_wire_4571)
    );

    bfr new_Jinkela_buffer_2187 (
        .din(new_Jinkela_wire_2563),
        .dout(new_Jinkela_wire_2564)
    );

    bfr new_Jinkela_buffer_3877 (
        .din(new_Jinkela_wire_4547),
        .dout(new_Jinkela_wire_4548)
    );

    bfr new_Jinkela_buffer_2130 (
        .din(new_Jinkela_wire_2504),
        .dout(new_Jinkela_wire_2505)
    );

    spl2 new_Jinkela_splitter_559 (
        .a(n_0324_),
        .b(new_Jinkela_wire_7834),
        .c(new_Jinkela_wire_7835)
    );

    bfr new_Jinkela_buffer_6376 (
        .din(new_Jinkela_wire_7781),
        .dout(new_Jinkela_wire_7782)
    );

    bfr new_Jinkela_buffer_3957 (
        .din(n_0805_),
        .dout(new_Jinkela_wire_4630)
    );

    bfr new_Jinkela_buffer_2206 (
        .din(new_Jinkela_wire_2588),
        .dout(new_Jinkela_wire_2589)
    );

    bfr new_Jinkela_buffer_6402 (
        .din(new_Jinkela_wire_7809),
        .dout(new_Jinkela_wire_7810)
    );

    bfr new_Jinkela_buffer_3878 (
        .din(new_Jinkela_wire_4548),
        .dout(new_Jinkela_wire_4549)
    );

    bfr new_Jinkela_buffer_2131 (
        .din(new_Jinkela_wire_2505),
        .dout(new_Jinkela_wire_2506)
    );

    bfr new_Jinkela_buffer_6377 (
        .din(new_Jinkela_wire_7782),
        .dout(new_Jinkela_wire_7783)
    );

    bfr new_Jinkela_buffer_3901 (
        .din(new_Jinkela_wire_4571),
        .dout(new_Jinkela_wire_4572)
    );

    bfr new_Jinkela_buffer_673 (
        .din(new_Jinkela_wire_725),
        .dout(new_Jinkela_wire_726)
    );

    bfr new_Jinkela_buffer_2188 (
        .din(new_Jinkela_wire_2564),
        .dout(new_Jinkela_wire_2565)
    );

    spl2 new_Jinkela_splitter_556 (
        .a(new_Jinkela_wire_7821),
        .b(new_Jinkela_wire_7822),
        .c(new_Jinkela_wire_7823)
    );

    bfr new_Jinkela_buffer_3879 (
        .din(new_Jinkela_wire_4549),
        .dout(new_Jinkela_wire_4550)
    );

    bfr new_Jinkela_buffer_2132 (
        .din(new_Jinkela_wire_2506),
        .dout(new_Jinkela_wire_2507)
    );

    bfr new_Jinkela_buffer_6378 (
        .din(new_Jinkela_wire_7783),
        .dout(new_Jinkela_wire_7784)
    );

    bfr new_Jinkela_buffer_2276 (
        .din(N299),
        .dout(new_Jinkela_wire_2663)
    );

    bfr new_Jinkela_buffer_6403 (
        .din(new_Jinkela_wire_7810),
        .dout(new_Jinkela_wire_7811)
    );

    bfr new_Jinkela_buffer_3880 (
        .din(new_Jinkela_wire_4550),
        .dout(new_Jinkela_wire_4551)
    );

    bfr new_Jinkela_buffer_2133 (
        .din(new_Jinkela_wire_2507),
        .dout(new_Jinkela_wire_2508)
    );

    bfr new_Jinkela_buffer_6379 (
        .din(new_Jinkela_wire_7784),
        .dout(new_Jinkela_wire_7785)
    );

    bfr new_Jinkela_buffer_3902 (
        .din(new_Jinkela_wire_4572),
        .dout(new_Jinkela_wire_4573)
    );

    bfr new_Jinkela_buffer_2208 (
        .din(new_Jinkela_wire_2592),
        .dout(new_Jinkela_wire_2593)
    );

    spl2 new_Jinkela_splitter_124 (
        .a(new_Jinkela_wire_2565),
        .b(new_Jinkela_wire_2566),
        .c(new_Jinkela_wire_2567)
    );

    bfr new_Jinkela_buffer_6412 (
        .din(new_Jinkela_wire_7825),
        .dout(new_Jinkela_wire_7826)
    );

    bfr new_Jinkela_buffer_3092 (
        .din(new_Jinkela_wire_3525),
        .dout(new_Jinkela_wire_3526)
    );

    and_bb n_1611_ (
        .a(new_Jinkela_wire_434),
        .b(new_Jinkela_wire_1253),
        .c(n_0879_)
    );

    and_bi n_2325_ (
        .a(n_0196_),
        .b(new_Jinkela_wire_3941),
        .c(n_0200_)
    );

    bfr new_Jinkela_buffer_3029 (
        .din(new_Jinkela_wire_3458),
        .dout(new_Jinkela_wire_3459)
    );

    bfr new_Jinkela_buffer_7222 (
        .din(new_Jinkela_wire_8952),
        .dout(new_Jinkela_wire_8953)
    );

    bfr new_Jinkela_buffer_2979 (
        .din(new_Jinkela_wire_3406),
        .dout(new_Jinkela_wire_3407)
    );

    and_bi n_1612_ (
        .a(new_Jinkela_wire_2585),
        .b(new_Jinkela_wire_1319),
        .c(n_0880_)
    );

    and_bi n_2326_ (
        .a(new_Jinkela_wire_6527),
        .b(n_0200_),
        .c(n_0201_)
    );

    bfr new_Jinkela_buffer_7203 (
        .din(new_Jinkela_wire_8916),
        .dout(new_Jinkela_wire_8917)
    );

    and_ii n_1613_ (
        .a(new_Jinkela_wire_8718),
        .b(new_Jinkela_wire_8753),
        .c(n_0881_)
    );

    and_ii n_2327_ (
        .a(n_0201_),
        .b(new_Jinkela_wire_9374),
        .c(n_0202_)
    );

    bfr new_Jinkela_buffer_2980 (
        .din(new_Jinkela_wire_3407),
        .dout(new_Jinkela_wire_3408)
    );

    and_bi n_1614_ (
        .a(new_Jinkela_wire_5230),
        .b(new_Jinkela_wire_5294),
        .c(n_0882_)
    );

    and_ii n_2328_ (
        .a(new_Jinkela_wire_8577),
        .b(new_Jinkela_wire_8929),
        .c(n_0203_)
    );

    bfr new_Jinkela_buffer_7204 (
        .din(new_Jinkela_wire_8917),
        .dout(new_Jinkela_wire_8918)
    );

    bfr new_Jinkela_buffer_3095 (
        .din(new_Jinkela_wire_3528),
        .dout(new_Jinkela_wire_3529)
    );

    and_bi n_1615_ (
        .a(new_Jinkela_wire_5292),
        .b(new_Jinkela_wire_5231),
        .c(n_0883_)
    );

    and_ii n_2329_ (
        .a(new_Jinkela_wire_10098),
        .b(new_Jinkela_wire_9539),
        .c(n_0204_)
    );

    bfr new_Jinkela_buffer_3030 (
        .din(new_Jinkela_wire_3459),
        .dout(new_Jinkela_wire_3460)
    );

    bfr new_Jinkela_buffer_7223 (
        .din(new_Jinkela_wire_8953),
        .dout(new_Jinkela_wire_8954)
    );

    bfr new_Jinkela_buffer_2981 (
        .din(new_Jinkela_wire_3408),
        .dout(new_Jinkela_wire_3409)
    );

    and_ii n_1616_ (
        .a(n_0883_),
        .b(n_0882_),
        .c(n_0884_)
    );

    or_bb n_2330_ (
        .a(n_0204_),
        .b(n_0203_),
        .c(n_0205_)
    );

    bfr new_Jinkela_buffer_7205 (
        .din(new_Jinkela_wire_8918),
        .dout(new_Jinkela_wire_8919)
    );

    or_ii n_1617_ (
        .a(new_Jinkela_wire_3517),
        .b(new_Jinkela_wire_1224),
        .c(n_0885_)
    );

    and_ii n_2331_ (
        .a(new_Jinkela_wire_5932),
        .b(n_0202_),
        .c(n_0206_)
    );

    bfr new_Jinkela_buffer_7250 (
        .din(new_Jinkela_wire_8980),
        .dout(new_Jinkela_wire_8981)
    );

    bfr new_Jinkela_buffer_2982 (
        .din(new_Jinkela_wire_3409),
        .dout(new_Jinkela_wire_3410)
    );

    and_bi n_1618_ (
        .a(new_Jinkela_wire_3535),
        .b(new_Jinkela_wire_1373),
        .c(n_0886_)
    );

    and_bb n_2332_ (
        .a(new_Jinkela_wire_3695),
        .b(new_Jinkela_wire_6011),
        .c(n_0207_)
    );

    bfr new_Jinkela_buffer_7206 (
        .din(new_Jinkela_wire_8919),
        .dout(new_Jinkela_wire_8920)
    );

    bfr new_Jinkela_buffer_3093 (
        .din(new_Jinkela_wire_3526),
        .dout(new_Jinkela_wire_3527)
    );

    and_bi n_1619_ (
        .a(new_Jinkela_wire_3578),
        .b(new_Jinkela_wire_4522),
        .c(n_0887_)
    );

    and_ii n_2333_ (
        .a(new_Jinkela_wire_8293),
        .b(new_Jinkela_wire_6402),
        .c(n_0208_)
    );

    bfr new_Jinkela_buffer_3031 (
        .din(new_Jinkela_wire_3460),
        .dout(new_Jinkela_wire_3461)
    );

    bfr new_Jinkela_buffer_7224 (
        .din(new_Jinkela_wire_8954),
        .dout(new_Jinkela_wire_8955)
    );

    bfr new_Jinkela_buffer_2983 (
        .din(new_Jinkela_wire_3410),
        .dout(new_Jinkela_wire_3411)
    );

    or_ii n_1620_ (
        .a(new_Jinkela_wire_2462),
        .b(new_Jinkela_wire_1310),
        .c(n_0888_)
    );

    or_bb n_2334_ (
        .a(new_Jinkela_wire_4632),
        .b(new_Jinkela_wire_4861),
        .c(n_0209_)
    );

    bfr new_Jinkela_buffer_7207 (
        .din(new_Jinkela_wire_8920),
        .dout(new_Jinkela_wire_8921)
    );

    and_bi n_1621_ (
        .a(new_Jinkela_wire_2068),
        .b(new_Jinkela_wire_1382),
        .c(n_0889_)
    );

    and_bb n_2335_ (
        .a(new_Jinkela_wire_8574),
        .b(new_Jinkela_wire_8928),
        .c(n_0210_)
    );

    bfr new_Jinkela_buffer_2984 (
        .din(new_Jinkela_wire_3411),
        .dout(new_Jinkela_wire_3412)
    );

    and_bi n_1622_ (
        .a(new_Jinkela_wire_3577),
        .b(new_Jinkela_wire_7928),
        .c(n_0890_)
    );

    and_bb n_2336_ (
        .a(new_Jinkela_wire_8291),
        .b(new_Jinkela_wire_6401),
        .c(n_0211_)
    );

    bfr new_Jinkela_buffer_7208 (
        .din(new_Jinkela_wire_8921),
        .dout(new_Jinkela_wire_8922)
    );

    spl3L new_Jinkela_splitter_148 (
        .a(N5),
        .d(new_Jinkela_wire_3536),
        .b(new_Jinkela_wire_3537),
        .c(new_Jinkela_wire_3538)
    );

    and_ii n_1623_ (
        .a(new_Jinkela_wire_7685),
        .b(new_Jinkela_wire_9471),
        .c(n_0891_)
    );

    or_bb n_2337_ (
        .a(n_0211_),
        .b(n_0210_),
        .c(n_0212_)
    );

    bfr new_Jinkela_buffer_3032 (
        .din(new_Jinkela_wire_3461),
        .dout(new_Jinkela_wire_3462)
    );

    bfr new_Jinkela_buffer_7225 (
        .din(new_Jinkela_wire_8955),
        .dout(new_Jinkela_wire_8956)
    );

    bfr new_Jinkela_buffer_2985 (
        .din(new_Jinkela_wire_3412),
        .dout(new_Jinkela_wire_3413)
    );

    and_bb n_1624_ (
        .a(new_Jinkela_wire_7686),
        .b(new_Jinkela_wire_9470),
        .c(n_0892_)
    );

    or_bb n_2338_ (
        .a(new_Jinkela_wire_9925),
        .b(n_0209_),
        .c(n_0213_)
    );

    bfr new_Jinkela_buffer_7209 (
        .din(new_Jinkela_wire_8922),
        .dout(new_Jinkela_wire_8923)
    );

    and_ii n_1625_ (
        .a(n_0892_),
        .b(n_0891_),
        .c(n_0893_)
    );

    and_ii n_2339_ (
        .a(new_Jinkela_wire_6434),
        .b(n_0206_),
        .c(n_0214_)
    );

    bfr new_Jinkela_buffer_3102 (
        .din(N114),
        .dout(new_Jinkela_wire_3539)
    );

    bfr new_Jinkela_buffer_7251 (
        .din(new_Jinkela_wire_8981),
        .dout(new_Jinkela_wire_8982)
    );

    bfr new_Jinkela_buffer_2986 (
        .din(new_Jinkela_wire_3413),
        .dout(new_Jinkela_wire_3414)
    );

    and_bi n_1626_ (
        .a(new_Jinkela_wire_9301),
        .b(new_Jinkela_wire_4976),
        .c(n_0894_)
    );

    and_bi n_2340_ (
        .a(new_Jinkela_wire_4631),
        .b(new_Jinkela_wire_4860),
        .c(n_0215_)
    );

    bfr new_Jinkela_buffer_7226 (
        .din(new_Jinkela_wire_8956),
        .dout(new_Jinkela_wire_8957)
    );

    bfr new_Jinkela_buffer_3096 (
        .din(new_Jinkela_wire_3529),
        .dout(new_Jinkela_wire_3530)
    );

    and_bi n_1627_ (
        .a(new_Jinkela_wire_4975),
        .b(new_Jinkela_wire_9300),
        .c(n_0895_)
    );

    and_ii n_2341_ (
        .a(new_Jinkela_wire_3694),
        .b(new_Jinkela_wire_6012),
        .c(n_0216_)
    );

    bfr new_Jinkela_buffer_3033 (
        .din(new_Jinkela_wire_3462),
        .dout(new_Jinkela_wire_3463)
    );

    spl2 new_Jinkela_splitter_696 (
        .a(n_0644_),
        .b(new_Jinkela_wire_9000),
        .c(new_Jinkela_wire_9001)
    );

    bfr new_Jinkela_buffer_2987 (
        .din(new_Jinkela_wire_3414),
        .dout(new_Jinkela_wire_3415)
    );

    spl2 new_Jinkela_splitter_700 (
        .a(n_0863_),
        .b(new_Jinkela_wire_9016),
        .c(new_Jinkela_wire_9017)
    );

    and_ii n_1628_ (
        .a(n_0895_),
        .b(n_0894_),
        .c(n_0896_)
    );

    and_ii n_2342_ (
        .a(new_Jinkela_wire_6391),
        .b(new_Jinkela_wire_4236),
        .c(n_0217_)
    );

    bfr new_Jinkela_buffer_7227 (
        .din(new_Jinkela_wire_8957),
        .dout(new_Jinkela_wire_8958)
    );

    and_bi n_1629_ (
        .a(new_Jinkela_wire_7245),
        .b(new_Jinkela_wire_3704),
        .c(n_0897_)
    );

    or_bb n_2343_ (
        .a(n_0217_),
        .b(n_0216_),
        .c(n_0218_)
    );

    bfr new_Jinkela_buffer_7252 (
        .din(new_Jinkela_wire_8982),
        .dout(new_Jinkela_wire_8983)
    );

    bfr new_Jinkela_buffer_2988 (
        .din(new_Jinkela_wire_3415),
        .dout(new_Jinkela_wire_3416)
    );

    and_bi n_1630_ (
        .a(new_Jinkela_wire_3703),
        .b(new_Jinkela_wire_7244),
        .c(n_0898_)
    );

    or_bb n_2344_ (
        .a(new_Jinkela_wire_5012),
        .b(n_0215_),
        .c(n_0219_)
    );

    bfr new_Jinkela_buffer_7228 (
        .din(new_Jinkela_wire_8958),
        .dout(new_Jinkela_wire_8959)
    );

    bfr new_Jinkela_buffer_3099 (
        .din(new_Jinkela_wire_3532),
        .dout(new_Jinkela_wire_3533)
    );

    and_ii n_1631_ (
        .a(n_0898_),
        .b(n_0897_),
        .c(n_0899_)
    );

    and_ii n_2345_ (
        .a(new_Jinkela_wire_8101),
        .b(n_0214_),
        .c(n_0220_)
    );

    bfr new_Jinkela_buffer_3034 (
        .din(new_Jinkela_wire_3463),
        .dout(new_Jinkela_wire_3464)
    );

    bfr new_Jinkela_buffer_7265 (
        .din(new_net_2519),
        .dout(new_Jinkela_wire_9002)
    );

    bfr new_Jinkela_buffer_2989 (
        .din(new_Jinkela_wire_3416),
        .dout(new_Jinkela_wire_3417)
    );

    spl2 new_Jinkela_splitter_698 (
        .a(n_1231_),
        .b(new_Jinkela_wire_9007),
        .c(new_Jinkela_wire_9008)
    );

    or_bi n_1632_ (
        .a(new_Jinkela_wire_3777),
        .b(new_Jinkela_wire_3852),
        .c(n_0900_)
    );

    and_ii n_2346_ (
        .a(new_Jinkela_wire_7277),
        .b(new_Jinkela_wire_8274),
        .c(n_0221_)
    );

    bfr new_Jinkela_buffer_7229 (
        .din(new_Jinkela_wire_8959),
        .dout(new_Jinkela_wire_8960)
    );

    and_bi n_1633_ (
        .a(new_Jinkela_wire_3776),
        .b(new_Jinkela_wire_3851),
        .c(n_0901_)
    );

    and_ii n_2347_ (
        .a(new_Jinkela_wire_8187),
        .b(new_Jinkela_wire_8002),
        .c(n_0222_)
    );

    bfr new_Jinkela_buffer_7253 (
        .din(new_Jinkela_wire_8983),
        .dout(new_Jinkela_wire_8984)
    );

    bfr new_Jinkela_buffer_2990 (
        .din(new_Jinkela_wire_3417),
        .dout(new_Jinkela_wire_3418)
    );

    and_bi n_1634_ (
        .a(n_0900_),
        .b(n_0901_),
        .c(n_0902_)
    );

    or_bb n_2348_ (
        .a(n_0222_),
        .b(n_0221_),
        .c(n_0223_)
    );

    bfr new_Jinkela_buffer_7230 (
        .din(new_Jinkela_wire_8960),
        .dout(new_Jinkela_wire_8961)
    );

    bfr new_Jinkela_buffer_3097 (
        .din(new_Jinkela_wire_3530),
        .dout(new_Jinkela_wire_3531)
    );

    or_bb n_1635_ (
        .a(n_0902_),
        .b(n_0845_),
        .c(n_0903_)
    );

    and_bb n_2349_ (
        .a(new_Jinkela_wire_3582),
        .b(new_Jinkela_wire_6338),
        .c(n_0224_)
    );

    bfr new_Jinkela_buffer_3035 (
        .din(new_Jinkela_wire_3464),
        .dout(new_Jinkela_wire_3465)
    );

    spl4L new_Jinkela_splitter_697 (
        .a(n_1151_),
        .d(new_Jinkela_wire_9003),
        .b(new_Jinkela_wire_9004),
        .e(new_Jinkela_wire_9005),
        .c(new_Jinkela_wire_9006)
    );

    bfr new_Jinkela_buffer_2991 (
        .din(new_Jinkela_wire_3418),
        .dout(new_Jinkela_wire_3419)
    );

    or_bb n_1636_ (
        .a(n_0903_),
        .b(n_0801_),
        .c(new_net_4)
    );

    and_bb n_2350_ (
        .a(new_Jinkela_wire_7276),
        .b(new_Jinkela_wire_8273),
        .c(n_0225_)
    );

    bfr new_Jinkela_buffer_7231 (
        .din(new_Jinkela_wire_8961),
        .dout(new_Jinkela_wire_8962)
    );

    or_bi n_1637_ (
        .a(new_Jinkela_wire_1204),
        .b(new_Jinkela_wire_3542),
        .c(n_0904_)
    );

    and_bb n_2351_ (
        .a(new_Jinkela_wire_8184),
        .b(new_Jinkela_wire_8001),
        .c(n_0226_)
    );

    bfr new_Jinkela_buffer_7254 (
        .din(new_Jinkela_wire_8984),
        .dout(new_Jinkela_wire_8985)
    );

    bfr new_Jinkela_buffer_2992 (
        .din(new_Jinkela_wire_3419),
        .dout(new_Jinkela_wire_3420)
    );

    and_bi n_1638_ (
        .a(new_Jinkela_wire_1257),
        .b(new_Jinkela_wire_2001),
        .c(n_0905_)
    );

    or_bb n_2352_ (
        .a(new_Jinkela_wire_8298),
        .b(new_Jinkela_wire_9648),
        .c(n_0227_)
    );

    bfr new_Jinkela_buffer_7232 (
        .din(new_Jinkela_wire_8962),
        .dout(new_Jinkela_wire_8963)
    );

    and_bi n_1639_ (
        .a(n_0904_),
        .b(n_0905_),
        .c(n_0906_)
    );

    or_bb n_2353_ (
        .a(n_0227_),
        .b(new_Jinkela_wire_10381),
        .c(n_0228_)
    );

    bfr new_Jinkela_buffer_3036 (
        .din(new_Jinkela_wire_3465),
        .dout(new_Jinkela_wire_3466)
    );

    bfr new_Jinkela_buffer_7269 (
        .din(n_0570_),
        .dout(new_Jinkela_wire_9014)
    );

    bfr new_Jinkela_buffer_2993 (
        .din(new_Jinkela_wire_3420),
        .dout(new_Jinkela_wire_3421)
    );

    and_bi n_1640_ (
        .a(new_Jinkela_wire_1826),
        .b(new_Jinkela_wire_1336),
        .c(n_0907_)
    );

    and_ii n_2354_ (
        .a(n_0228_),
        .b(new_Jinkela_wire_7502),
        .c(n_0229_)
    );

    bfr new_Jinkela_buffer_7233 (
        .din(new_Jinkela_wire_8963),
        .dout(new_Jinkela_wire_8964)
    );

    and_bi n_1641_ (
        .a(new_Jinkela_wire_1213),
        .b(new_Jinkela_wire_2820),
        .c(n_0908_)
    );

    and_ii n_2355_ (
        .a(new_Jinkela_wire_9004),
        .b(new_Jinkela_wire_4518),
        .c(n_0230_)
    );

    bfr new_Jinkela_buffer_7255 (
        .din(new_Jinkela_wire_8985),
        .dout(new_Jinkela_wire_8986)
    );

    bfr new_Jinkela_buffer_2994 (
        .din(new_Jinkela_wire_3421),
        .dout(new_Jinkela_wire_3422)
    );

    and_ii n_1642_ (
        .a(n_0908_),
        .b(n_0907_),
        .c(n_0909_)
    );

    and_ii n_2356_ (
        .a(new_Jinkela_wire_3579),
        .b(new_Jinkela_wire_6339),
        .c(n_0231_)
    );

    bfr new_Jinkela_buffer_7234 (
        .din(new_Jinkela_wire_8964),
        .dout(new_Jinkela_wire_8965)
    );

    bfr new_Jinkela_buffer_3100 (
        .din(new_Jinkela_wire_3533),
        .dout(new_Jinkela_wire_3534)
    );

    and_ii n_1643_ (
        .a(new_Jinkela_wire_8765),
        .b(new_Jinkela_wire_5576),
        .c(n_0910_)
    );

    and_ii n_2357_ (
        .a(n_0231_),
        .b(n_0230_),
        .c(n_0232_)
    );

    bfr new_Jinkela_buffer_3037 (
        .din(new_Jinkela_wire_3466),
        .dout(new_Jinkela_wire_3467)
    );

    bfr new_Jinkela_buffer_7266 (
        .din(n_1241_),
        .dout(new_Jinkela_wire_9009)
    );

    bfr new_Jinkela_buffer_2995 (
        .din(new_Jinkela_wire_3422),
        .dout(new_Jinkela_wire_3423)
    );

    and_bb n_1644_ (
        .a(new_Jinkela_wire_8764),
        .b(new_Jinkela_wire_5575),
        .c(n_0911_)
    );

    and_bb n_2358_ (
        .a(new_Jinkela_wire_6393),
        .b(new_Jinkela_wire_4237),
        .c(n_0233_)
    );

    bfr new_Jinkela_buffer_7235 (
        .din(new_Jinkela_wire_8965),
        .dout(new_Jinkela_wire_8966)
    );

    and_ii n_1645_ (
        .a(n_0911_),
        .b(n_0910_),
        .c(n_0912_)
    );

    and_bb n_2359_ (
        .a(new_Jinkela_wire_9003),
        .b(new_Jinkela_wire_4519),
        .c(n_0234_)
    );

    bfr new_Jinkela_buffer_7256 (
        .din(new_Jinkela_wire_8986),
        .dout(new_Jinkela_wire_8987)
    );

    bfr new_Jinkela_buffer_2996 (
        .din(new_Jinkela_wire_3423),
        .dout(new_Jinkela_wire_3424)
    );

    and_bi n_1646_ (
        .a(new_Jinkela_wire_1822),
        .b(new_Jinkela_wire_1345),
        .c(n_0913_)
    );

    and_ii n_2360_ (
        .a(n_0234_),
        .b(n_0233_),
        .c(n_0235_)
    );

    bfr new_Jinkela_buffer_7236 (
        .din(new_Jinkela_wire_8966),
        .dout(new_Jinkela_wire_8967)
    );

    and_bi n_1647_ (
        .a(new_Jinkela_wire_1368),
        .b(new_Jinkela_wire_2482),
        .c(n_0914_)
    );

    and_bb n_2361_ (
        .a(new_Jinkela_wire_9468),
        .b(new_Jinkela_wire_9291),
        .c(n_0236_)
    );

    bfr new_Jinkela_buffer_3038 (
        .din(new_Jinkela_wire_3467),
        .dout(new_Jinkela_wire_3468)
    );

    bfr new_Jinkela_buffer_7267 (
        .din(new_Jinkela_wire_9009),
        .dout(new_Jinkela_wire_9010)
    );

    bfr new_Jinkela_buffer_2997 (
        .din(new_Jinkela_wire_3424),
        .dout(new_Jinkela_wire_3425)
    );

    and_ii n_1648_ (
        .a(n_0914_),
        .b(n_0913_),
        .c(n_0915_)
    );

    or_ii n_2362_ (
        .a(new_Jinkela_wire_8570),
        .b(new_Jinkela_wire_8440),
        .c(n_0237_)
    );

    bfr new_Jinkela_buffer_7237 (
        .din(new_Jinkela_wire_8967),
        .dout(new_Jinkela_wire_8968)
    );

    or_bi n_1649_ (
        .a(new_Jinkela_wire_1314),
        .b(new_Jinkela_wire_604),
        .c(n_0916_)
    );

    and_ii n_2363_ (
        .a(new_Jinkela_wire_5009),
        .b(n_0220_),
        .c(n_0238_)
    );

    bfr new_Jinkela_buffer_3106 (
        .din(N50),
        .dout(new_Jinkela_wire_3543)
    );

    bfr new_Jinkela_buffer_7257 (
        .din(new_Jinkela_wire_8987),
        .dout(new_Jinkela_wire_8988)
    );

    bfr new_Jinkela_buffer_2998 (
        .din(new_Jinkela_wire_3425),
        .dout(new_Jinkela_wire_3426)
    );

    and_bi n_1650_ (
        .a(new_Jinkela_wire_1324),
        .b(new_Jinkela_wire_613),
        .c(n_0917_)
    );

    and_bi n_2364_ (
        .a(new_Jinkela_wire_8439),
        .b(new_Jinkela_wire_9295),
        .c(n_0239_)
    );

    bfr new_Jinkela_buffer_7238 (
        .din(new_Jinkela_wire_8968),
        .dout(new_Jinkela_wire_8969)
    );

    bfr new_Jinkela_buffer_3101 (
        .din(new_Jinkela_wire_3534),
        .dout(new_Jinkela_wire_3535)
    );

    and_bi n_1651_ (
        .a(n_0916_),
        .b(n_0917_),
        .c(n_0918_)
    );

    and_bi n_2365_ (
        .a(new_Jinkela_wire_7500),
        .b(new_Jinkela_wire_8300),
        .c(n_0240_)
    );

    bfr new_Jinkela_buffer_3039 (
        .din(new_Jinkela_wire_3468),
        .dout(new_Jinkela_wire_3469)
    );

    spl4L new_Jinkela_splitter_701 (
        .a(n_0804_),
        .d(new_Jinkela_wire_9018),
        .b(new_Jinkela_wire_9019),
        .e(new_Jinkela_wire_9020),
        .c(new_Jinkela_wire_9021)
    );

    bfr new_Jinkela_buffer_2999 (
        .din(new_Jinkela_wire_3426),
        .dout(new_Jinkela_wire_3427)
    );

    and_bi n_1652_ (
        .a(new_Jinkela_wire_10557),
        .b(new_Jinkela_wire_9151),
        .c(n_0919_)
    );

    or_bb n_2366_ (
        .a(new_Jinkela_wire_8360),
        .b(n_0239_),
        .c(n_0241_)
    );

    bfr new_Jinkela_buffer_7239 (
        .din(new_Jinkela_wire_8969),
        .dout(new_Jinkela_wire_8970)
    );

    bfr new_Jinkela_buffer_8376 (
        .din(new_Jinkela_wire_10521),
        .dout(new_Jinkela_wire_10522)
    );

    bfr new_Jinkela_buffer_8459 (
        .din(new_Jinkela_wire_10630),
        .dout(new_Jinkela_wire_10631)
    );

    bfr new_Jinkela_buffer_8385 (
        .din(new_Jinkela_wire_10538),
        .dout(new_Jinkela_wire_10539)
    );

    bfr new_Jinkela_buffer_8402 (
        .din(new_Jinkela_wire_10567),
        .dout(new_Jinkela_wire_10568)
    );

    bfr new_Jinkela_buffer_8386 (
        .din(new_Jinkela_wire_10539),
        .dout(new_Jinkela_wire_10540)
    );

    bfr new_Jinkela_buffer_8387 (
        .din(new_Jinkela_wire_10540),
        .dout(new_Jinkela_wire_10541)
    );

    bfr new_Jinkela_buffer_8403 (
        .din(new_Jinkela_wire_10568),
        .dout(new_Jinkela_wire_10569)
    );

    bfr new_Jinkela_buffer_8388 (
        .din(new_Jinkela_wire_10541),
        .dout(new_Jinkela_wire_10542)
    );

    bfr new_Jinkela_buffer_8389 (
        .din(new_Jinkela_wire_10542),
        .dout(new_Jinkela_wire_10543)
    );

    bfr new_Jinkela_buffer_8404 (
        .din(new_Jinkela_wire_10569),
        .dout(new_Jinkela_wire_10570)
    );

    bfr new_Jinkela_buffer_8390 (
        .din(new_Jinkela_wire_10543),
        .dout(new_Jinkela_wire_10544)
    );

    bfr new_Jinkela_buffer_8460 (
        .din(new_Jinkela_wire_10631),
        .dout(new_Jinkela_wire_10632)
    );

    bfr new_Jinkela_buffer_8391 (
        .din(new_Jinkela_wire_10544),
        .dout(new_Jinkela_wire_10545)
    );

    bfr new_Jinkela_buffer_8405 (
        .din(new_Jinkela_wire_10570),
        .dout(new_Jinkela_wire_10571)
    );

    bfr new_Jinkela_buffer_8392 (
        .din(new_Jinkela_wire_10545),
        .dout(new_Jinkela_wire_10546)
    );

    bfr new_Jinkela_buffer_8393 (
        .din(new_Jinkela_wire_10546),
        .dout(new_Jinkela_wire_10547)
    );

    bfr new_Jinkela_buffer_8406 (
        .din(new_Jinkela_wire_10571),
        .dout(new_Jinkela_wire_10572)
    );

    bfr new_Jinkela_buffer_8394 (
        .din(new_Jinkela_wire_10547),
        .dout(new_Jinkela_wire_10548)
    );

    bfr new_Jinkela_buffer_8395 (
        .din(new_Jinkela_wire_10548),
        .dout(new_Jinkela_wire_10549)
    );

    bfr new_Jinkela_buffer_8407 (
        .din(new_Jinkela_wire_10572),
        .dout(new_Jinkela_wire_10573)
    );

    bfr new_Jinkela_buffer_8396 (
        .din(new_Jinkela_wire_10549),
        .dout(new_Jinkela_wire_10550)
    );

    bfr new_Jinkela_buffer_8397 (
        .din(new_Jinkela_wire_10550),
        .dout(new_Jinkela_wire_10551)
    );

    bfr new_Jinkela_buffer_8408 (
        .din(new_Jinkela_wire_10573),
        .dout(new_Jinkela_wire_10574)
    );

    bfr new_Jinkela_buffer_8398 (
        .din(new_Jinkela_wire_10551),
        .dout(new_Jinkela_wire_10552)
    );

    bfr new_Jinkela_buffer_8399 (
        .din(new_Jinkela_wire_10552),
        .dout(new_Jinkela_wire_10553)
    );

    bfr new_Jinkela_buffer_8409 (
        .din(new_Jinkela_wire_10574),
        .dout(new_Jinkela_wire_10575)
    );

    bfr new_Jinkela_buffer_8410 (
        .din(new_Jinkela_wire_10575),
        .dout(new_Jinkela_wire_10576)
    );

    bfr new_Jinkela_buffer_8411 (
        .din(new_Jinkela_wire_10576),
        .dout(new_Jinkela_wire_10577)
    );

    bfr new_Jinkela_buffer_8412 (
        .din(new_Jinkela_wire_10577),
        .dout(new_Jinkela_wire_10578)
    );

    bfr new_Jinkela_buffer_8413 (
        .din(new_Jinkela_wire_10578),
        .dout(new_Jinkela_wire_10579)
    );

    bfr new_Jinkela_buffer_8414 (
        .din(new_Jinkela_wire_10579),
        .dout(new_Jinkela_wire_10580)
    );

    bfr new_Jinkela_buffer_5597 (
        .din(new_Jinkela_wire_6711),
        .dout(new_Jinkela_wire_6712)
    );

    bfr new_Jinkela_buffer_5527 (
        .din(new_Jinkela_wire_6631),
        .dout(new_Jinkela_wire_6632)
    );

    bfr new_Jinkela_buffer_5548 (
        .din(new_Jinkela_wire_6652),
        .dout(new_Jinkela_wire_6653)
    );

    bfr new_Jinkela_buffer_5528 (
        .din(new_Jinkela_wire_6632),
        .dout(new_Jinkela_wire_6633)
    );

    bfr new_Jinkela_buffer_5570 (
        .din(new_Jinkela_wire_6680),
        .dout(new_Jinkela_wire_6681)
    );

    bfr new_Jinkela_buffer_5529 (
        .din(new_Jinkela_wire_6633),
        .dout(new_Jinkela_wire_6634)
    );

    bfr new_Jinkela_buffer_5549 (
        .din(new_Jinkela_wire_6653),
        .dout(new_Jinkela_wire_6654)
    );

    bfr new_Jinkela_buffer_5530 (
        .din(new_Jinkela_wire_6634),
        .dout(new_Jinkela_wire_6635)
    );

    bfr new_Jinkela_buffer_5531 (
        .din(new_Jinkela_wire_6635),
        .dout(new_Jinkela_wire_6636)
    );

    bfr new_Jinkela_buffer_5550 (
        .din(new_Jinkela_wire_6654),
        .dout(new_Jinkela_wire_6655)
    );

    bfr new_Jinkela_buffer_5532 (
        .din(new_Jinkela_wire_6636),
        .dout(new_Jinkela_wire_6637)
    );

    bfr new_Jinkela_buffer_5571 (
        .din(new_Jinkela_wire_6681),
        .dout(new_Jinkela_wire_6682)
    );

    bfr new_Jinkela_buffer_5533 (
        .din(new_Jinkela_wire_6637),
        .dout(new_Jinkela_wire_6638)
    );

    bfr new_Jinkela_buffer_5551 (
        .din(new_Jinkela_wire_6655),
        .dout(new_Jinkela_wire_6656)
    );

    bfr new_Jinkela_buffer_5534 (
        .din(new_Jinkela_wire_6638),
        .dout(new_Jinkela_wire_6639)
    );

    bfr new_Jinkela_buffer_5598 (
        .din(new_Jinkela_wire_6712),
        .dout(new_Jinkela_wire_6713)
    );

    bfr new_Jinkela_buffer_5552 (
        .din(new_Jinkela_wire_6656),
        .dout(new_Jinkela_wire_6657)
    );

    bfr new_Jinkela_buffer_5572 (
        .din(new_Jinkela_wire_6682),
        .dout(new_Jinkela_wire_6683)
    );

    bfr new_Jinkela_buffer_5553 (
        .din(new_Jinkela_wire_6657),
        .dout(new_Jinkela_wire_6658)
    );

    bfr new_Jinkela_buffer_5554 (
        .din(new_Jinkela_wire_6658),
        .dout(new_Jinkela_wire_6659)
    );

    bfr new_Jinkela_buffer_5573 (
        .din(new_Jinkela_wire_6683),
        .dout(new_Jinkela_wire_6684)
    );

    bfr new_Jinkela_buffer_5555 (
        .din(new_Jinkela_wire_6659),
        .dout(new_Jinkela_wire_6660)
    );

    bfr new_Jinkela_buffer_5599 (
        .din(new_Jinkela_wire_6713),
        .dout(new_Jinkela_wire_6714)
    );

    bfr new_Jinkela_buffer_5556 (
        .din(new_Jinkela_wire_6660),
        .dout(new_Jinkela_wire_6661)
    );

    bfr new_Jinkela_buffer_5574 (
        .din(new_Jinkela_wire_6684),
        .dout(new_Jinkela_wire_6685)
    );

    bfr new_Jinkela_buffer_5557 (
        .din(new_Jinkela_wire_6661),
        .dout(new_Jinkela_wire_6662)
    );

    spl2 new_Jinkela_splitter_439 (
        .a(new_Jinkela_wire_6785),
        .b(new_Jinkela_wire_6786),
        .c(new_Jinkela_wire_6787)
    );

    bfr new_Jinkela_buffer_5558 (
        .din(new_Jinkela_wire_6662),
        .dout(new_Jinkela_wire_6663)
    );

    bfr new_Jinkela_buffer_5575 (
        .din(new_Jinkela_wire_6685),
        .dout(new_Jinkela_wire_6686)
    );

    bfr new_Jinkela_buffer_5559 (
        .din(new_Jinkela_wire_6663),
        .dout(new_Jinkela_wire_6664)
    );

    bfr new_Jinkela_buffer_5627 (
        .din(new_Jinkela_wire_6747),
        .dout(new_Jinkela_wire_6748)
    );

    bfr new_Jinkela_buffer_5600 (
        .din(new_Jinkela_wire_6714),
        .dout(new_Jinkela_wire_6715)
    );

    bfr new_Jinkela_buffer_5560 (
        .din(new_Jinkela_wire_6664),
        .dout(new_Jinkela_wire_6665)
    );

    bfr new_Jinkela_buffer_5576 (
        .din(new_Jinkela_wire_6686),
        .dout(new_Jinkela_wire_6687)
    );

    bfr new_Jinkela_buffer_5561 (
        .din(new_Jinkela_wire_6665),
        .dout(new_Jinkela_wire_6666)
    );

    bfr new_Jinkela_buffer_5562 (
        .din(new_Jinkela_wire_6666),
        .dout(new_Jinkela_wire_6667)
    );

    bfr new_Jinkela_buffer_5577 (
        .din(new_Jinkela_wire_6687),
        .dout(new_Jinkela_wire_6688)
    );

    bfr new_Jinkela_buffer_5563 (
        .din(new_Jinkela_wire_6667),
        .dout(new_Jinkela_wire_6668)
    );

    bfr new_Jinkela_buffer_5647 (
        .din(new_Jinkela_wire_6771),
        .dout(new_Jinkela_wire_6772)
    );

    bfr new_Jinkela_buffer_5601 (
        .din(new_Jinkela_wire_6715),
        .dout(new_Jinkela_wire_6716)
    );

    bfr new_Jinkela_buffer_5564 (
        .din(new_Jinkela_wire_6668),
        .dout(new_Jinkela_wire_6669)
    );

    bfr new_Jinkela_buffer_5578 (
        .din(new_Jinkela_wire_6688),
        .dout(new_Jinkela_wire_6689)
    );

    bfr new_Jinkela_buffer_806 (
        .din(new_Jinkela_wire_866),
        .dout(new_Jinkela_wire_867)
    );

    bfr new_Jinkela_buffer_894 (
        .din(new_Jinkela_wire_964),
        .dout(new_Jinkela_wire_965)
    );

    bfr new_Jinkela_buffer_844 (
        .din(new_Jinkela_wire_909),
        .dout(new_Jinkela_wire_910)
    );

    bfr new_Jinkela_buffer_1023 (
        .din(N307),
        .dout(new_Jinkela_wire_1098)
    );

    spl2 new_Jinkela_splitter_34 (
        .a(N245),
        .b(new_Jinkela_wire_1165),
        .c(new_Jinkela_wire_1166)
    );

    bfr new_Jinkela_buffer_845 (
        .din(new_Jinkela_wire_910),
        .dout(new_Jinkela_wire_911)
    );

    bfr new_Jinkela_buffer_895 (
        .din(new_Jinkela_wire_965),
        .dout(new_Jinkela_wire_966)
    );

    bfr new_Jinkela_buffer_846 (
        .din(new_Jinkela_wire_911),
        .dout(new_Jinkela_wire_912)
    );

    bfr new_Jinkela_buffer_952 (
        .din(new_Jinkela_wire_1026),
        .dout(new_Jinkela_wire_1027)
    );

    bfr new_Jinkela_buffer_847 (
        .din(new_Jinkela_wire_912),
        .dout(new_Jinkela_wire_913)
    );

    bfr new_Jinkela_buffer_896 (
        .din(new_Jinkela_wire_966),
        .dout(new_Jinkela_wire_967)
    );

    bfr new_Jinkela_buffer_848 (
        .din(new_Jinkela_wire_913),
        .dout(new_Jinkela_wire_914)
    );

    bfr new_Jinkela_buffer_1017 (
        .din(new_Jinkela_wire_1091),
        .dout(new_Jinkela_wire_1092)
    );

    bfr new_Jinkela_buffer_849 (
        .din(new_Jinkela_wire_914),
        .dout(new_Jinkela_wire_915)
    );

    bfr new_Jinkela_buffer_897 (
        .din(new_Jinkela_wire_967),
        .dout(new_Jinkela_wire_968)
    );

    bfr new_Jinkela_buffer_850 (
        .din(new_Jinkela_wire_915),
        .dout(new_Jinkela_wire_916)
    );

    bfr new_Jinkela_buffer_953 (
        .din(new_Jinkela_wire_1027),
        .dout(new_Jinkela_wire_1028)
    );

    bfr new_Jinkela_buffer_851 (
        .din(new_Jinkela_wire_916),
        .dout(new_Jinkela_wire_917)
    );

    bfr new_Jinkela_buffer_898 (
        .din(new_Jinkela_wire_968),
        .dout(new_Jinkela_wire_969)
    );

    bfr new_Jinkela_buffer_852 (
        .din(new_Jinkela_wire_917),
        .dout(new_Jinkela_wire_918)
    );

    bfr new_Jinkela_buffer_1020 (
        .din(new_Jinkela_wire_1094),
        .dout(new_Jinkela_wire_1095)
    );

    bfr new_Jinkela_buffer_853 (
        .din(new_Jinkela_wire_918),
        .dout(new_Jinkela_wire_919)
    );

    bfr new_Jinkela_buffer_899 (
        .din(new_Jinkela_wire_969),
        .dout(new_Jinkela_wire_970)
    );

    bfr new_Jinkela_buffer_854 (
        .din(new_Jinkela_wire_919),
        .dout(new_Jinkela_wire_920)
    );

    bfr new_Jinkela_buffer_954 (
        .din(new_Jinkela_wire_1028),
        .dout(new_Jinkela_wire_1029)
    );

    bfr new_Jinkela_buffer_855 (
        .din(new_Jinkela_wire_920),
        .dout(new_Jinkela_wire_921)
    );

    bfr new_Jinkela_buffer_900 (
        .din(new_Jinkela_wire_970),
        .dout(new_Jinkela_wire_971)
    );

    bfr new_Jinkela_buffer_856 (
        .din(new_Jinkela_wire_921),
        .dout(new_Jinkela_wire_922)
    );

    bfr new_Jinkela_buffer_1018 (
        .din(new_Jinkela_wire_1092),
        .dout(new_Jinkela_wire_1093)
    );

    bfr new_Jinkela_buffer_857 (
        .din(new_Jinkela_wire_922),
        .dout(new_Jinkela_wire_923)
    );

    bfr new_Jinkela_buffer_901 (
        .din(new_Jinkela_wire_971),
        .dout(new_Jinkela_wire_972)
    );

    bfr new_Jinkela_buffer_858 (
        .din(new_Jinkela_wire_923),
        .dout(new_Jinkela_wire_924)
    );

    bfr new_Jinkela_buffer_955 (
        .din(new_Jinkela_wire_1029),
        .dout(new_Jinkela_wire_1030)
    );

    bfr new_Jinkela_buffer_859 (
        .din(new_Jinkela_wire_924),
        .dout(new_Jinkela_wire_925)
    );

    bfr new_Jinkela_buffer_902 (
        .din(new_Jinkela_wire_972),
        .dout(new_Jinkela_wire_973)
    );

    bfr new_Jinkela_buffer_860 (
        .din(new_Jinkela_wire_925),
        .dout(new_Jinkela_wire_926)
    );

    bfr new_Jinkela_buffer_861 (
        .din(new_Jinkela_wire_926),
        .dout(new_Jinkela_wire_927)
    );

    bfr new_Jinkela_buffer_903 (
        .din(new_Jinkela_wire_973),
        .dout(new_Jinkela_wire_974)
    );

    bfr new_Jinkela_buffer_862 (
        .din(new_Jinkela_wire_927),
        .dout(new_Jinkela_wire_928)
    );

    bfr new_Jinkela_buffer_956 (
        .din(new_Jinkela_wire_1030),
        .dout(new_Jinkela_wire_1031)
    );

    bfr new_Jinkela_buffer_863 (
        .din(new_Jinkela_wire_928),
        .dout(new_Jinkela_wire_929)
    );

    bfr new_Jinkela_buffer_904 (
        .din(new_Jinkela_wire_974),
        .dout(new_Jinkela_wire_975)
    );

    bfr new_Jinkela_buffer_7258 (
        .din(new_Jinkela_wire_8988),
        .dout(new_Jinkela_wire_8989)
    );

    bfr new_Jinkela_buffer_3000 (
        .din(new_Jinkela_wire_3427),
        .dout(new_Jinkela_wire_3428)
    );

    bfr new_Jinkela_buffer_4701 (
        .din(new_Jinkela_wire_5606),
        .dout(new_Jinkela_wire_5607)
    );

    bfr new_Jinkela_buffer_7240 (
        .din(new_Jinkela_wire_8970),
        .dout(new_Jinkela_wire_8971)
    );

    bfr new_Jinkela_buffer_4731 (
        .din(new_Jinkela_wire_5650),
        .dout(new_Jinkela_wire_5651)
    );

    bfr new_Jinkela_buffer_3040 (
        .din(new_Jinkela_wire_3469),
        .dout(new_Jinkela_wire_3470)
    );

    bfr new_Jinkela_buffer_7270 (
        .din(new_Jinkela_wire_9014),
        .dout(new_Jinkela_wire_9015)
    );

    bfr new_Jinkela_buffer_3001 (
        .din(new_Jinkela_wire_3428),
        .dout(new_Jinkela_wire_3429)
    );

    bfr new_Jinkela_buffer_4702 (
        .din(new_Jinkela_wire_5607),
        .dout(new_Jinkela_wire_5608)
    );

    bfr new_Jinkela_buffer_7268 (
        .din(new_Jinkela_wire_9010),
        .dout(new_Jinkela_wire_9011)
    );

    bfr new_Jinkela_buffer_7241 (
        .din(new_Jinkela_wire_8971),
        .dout(new_Jinkela_wire_8972)
    );

    bfr new_Jinkela_buffer_4801 (
        .din(new_Jinkela_wire_5732),
        .dout(new_Jinkela_wire_5733)
    );

    bfr new_Jinkela_buffer_3103 (
        .din(new_Jinkela_wire_3539),
        .dout(new_Jinkela_wire_3540)
    );

    bfr new_Jinkela_buffer_7259 (
        .din(new_Jinkela_wire_8989),
        .dout(new_Jinkela_wire_8990)
    );

    bfr new_Jinkela_buffer_3002 (
        .din(new_Jinkela_wire_3429),
        .dout(new_Jinkela_wire_3430)
    );

    bfr new_Jinkela_buffer_4703 (
        .din(new_Jinkela_wire_5608),
        .dout(new_Jinkela_wire_5609)
    );

    bfr new_Jinkela_buffer_7242 (
        .din(new_Jinkela_wire_8972),
        .dout(new_Jinkela_wire_8973)
    );

    bfr new_Jinkela_buffer_3110 (
        .din(N209),
        .dout(new_Jinkela_wire_3547)
    );

    bfr new_Jinkela_buffer_4732 (
        .din(new_Jinkela_wire_5651),
        .dout(new_Jinkela_wire_5652)
    );

    bfr new_Jinkela_buffer_3041 (
        .din(new_Jinkela_wire_3470),
        .dout(new_Jinkela_wire_3471)
    );

    bfr new_Jinkela_buffer_4704 (
        .din(new_Jinkela_wire_5609),
        .dout(new_Jinkela_wire_5610)
    );

    bfr new_Jinkela_buffer_7243 (
        .din(new_Jinkela_wire_8973),
        .dout(new_Jinkela_wire_8974)
    );

    bfr new_Jinkela_buffer_3104 (
        .din(new_Jinkela_wire_3540),
        .dout(new_Jinkela_wire_3541)
    );

    bfr new_Jinkela_buffer_3042 (
        .din(new_Jinkela_wire_3471),
        .dout(new_Jinkela_wire_3472)
    );

    bfr new_Jinkela_buffer_4868 (
        .din(new_net_11),
        .dout(new_Jinkela_wire_5805)
    );

    bfr new_Jinkela_buffer_7260 (
        .din(new_Jinkela_wire_8990),
        .dout(new_Jinkela_wire_8991)
    );

    bfr new_Jinkela_buffer_4705 (
        .din(new_Jinkela_wire_5610),
        .dout(new_Jinkela_wire_5611)
    );

    bfr new_Jinkela_buffer_7244 (
        .din(new_Jinkela_wire_8974),
        .dout(new_Jinkela_wire_8975)
    );

    bfr new_Jinkela_buffer_3107 (
        .din(new_Jinkela_wire_3543),
        .dout(new_Jinkela_wire_3544)
    );

    bfr new_Jinkela_buffer_4733 (
        .din(new_Jinkela_wire_5652),
        .dout(new_Jinkela_wire_5653)
    );

    bfr new_Jinkela_buffer_3043 (
        .din(new_Jinkela_wire_3472),
        .dout(new_Jinkela_wire_3473)
    );

    bfr new_Jinkela_buffer_4706 (
        .din(new_Jinkela_wire_5611),
        .dout(new_Jinkela_wire_5612)
    );

    spl2 new_Jinkela_splitter_699 (
        .a(new_Jinkela_wire_9011),
        .b(new_Jinkela_wire_9012),
        .c(new_Jinkela_wire_9013)
    );

    bfr new_Jinkela_buffer_7245 (
        .din(new_Jinkela_wire_8975),
        .dout(new_Jinkela_wire_8976)
    );

    bfr new_Jinkela_buffer_3105 (
        .din(new_Jinkela_wire_3541),
        .dout(new_Jinkela_wire_3542)
    );

    spl3L new_Jinkela_splitter_352 (
        .a(new_Jinkela_wire_5680),
        .d(new_Jinkela_wire_5681),
        .b(new_Jinkela_wire_5682),
        .c(new_Jinkela_wire_5683)
    );

    bfr new_Jinkela_buffer_3044 (
        .din(new_Jinkela_wire_3473),
        .dout(new_Jinkela_wire_3474)
    );

    bfr new_Jinkela_buffer_7261 (
        .din(new_Jinkela_wire_8991),
        .dout(new_Jinkela_wire_8992)
    );

    bfr new_Jinkela_buffer_4707 (
        .din(new_Jinkela_wire_5612),
        .dout(new_Jinkela_wire_5613)
    );

    bfr new_Jinkela_buffer_7246 (
        .din(new_Jinkela_wire_8976),
        .dout(new_Jinkela_wire_8977)
    );

    bfr new_Jinkela_buffer_3114 (
        .din(N215),
        .dout(new_Jinkela_wire_3551)
    );

    bfr new_Jinkela_buffer_4734 (
        .din(new_Jinkela_wire_5653),
        .dout(new_Jinkela_wire_5654)
    );

    bfr new_Jinkela_buffer_3045 (
        .din(new_Jinkela_wire_3474),
        .dout(new_Jinkela_wire_3475)
    );

    bfr new_Jinkela_buffer_4708 (
        .din(new_Jinkela_wire_5613),
        .dout(new_Jinkela_wire_5614)
    );

    spl4L new_Jinkela_splitter_702 (
        .a(n_0683_),
        .d(new_Jinkela_wire_9022),
        .b(new_Jinkela_wire_9023),
        .e(new_Jinkela_wire_9024),
        .c(new_Jinkela_wire_9025)
    );

    bfr new_Jinkela_buffer_7262 (
        .din(new_Jinkela_wire_8992),
        .dout(new_Jinkela_wire_8993)
    );

    bfr new_Jinkela_buffer_3108 (
        .din(new_Jinkela_wire_3544),
        .dout(new_Jinkela_wire_3545)
    );

    spl3L new_Jinkela_splitter_351 (
        .a(new_Jinkela_wire_5677),
        .d(new_Jinkela_wire_5678),
        .b(new_Jinkela_wire_5679),
        .c(new_Jinkela_wire_5680)
    );

    bfr new_Jinkela_buffer_3046 (
        .din(new_Jinkela_wire_3475),
        .dout(new_Jinkela_wire_3476)
    );

    bfr new_Jinkela_buffer_4823 (
        .din(new_Jinkela_wire_5757),
        .dout(new_Jinkela_wire_5758)
    );

    spl3L new_Jinkela_splitter_705 (
        .a(n_0111_),
        .d(new_Jinkela_wire_9039),
        .b(new_Jinkela_wire_9040),
        .c(new_Jinkela_wire_9041)
    );

    bfr new_Jinkela_buffer_4709 (
        .din(new_Jinkela_wire_5614),
        .dout(new_Jinkela_wire_5615)
    );

    bfr new_Jinkela_buffer_7263 (
        .din(new_Jinkela_wire_8993),
        .dout(new_Jinkela_wire_8994)
    );

    bfr new_Jinkela_buffer_3111 (
        .din(new_Jinkela_wire_3547),
        .dout(new_Jinkela_wire_3548)
    );

    bfr new_Jinkela_buffer_4735 (
        .din(new_Jinkela_wire_5654),
        .dout(new_Jinkela_wire_5655)
    );

    bfr new_Jinkela_buffer_3047 (
        .din(new_Jinkela_wire_3476),
        .dout(new_Jinkela_wire_3477)
    );

    bfr new_Jinkela_buffer_4710 (
        .din(new_Jinkela_wire_5615),
        .dout(new_Jinkela_wire_5616)
    );

    spl2 new_Jinkela_splitter_704 (
        .a(n_0355_),
        .b(new_Jinkela_wire_9037),
        .c(new_Jinkela_wire_9038)
    );

    bfr new_Jinkela_buffer_3109 (
        .din(new_Jinkela_wire_3545),
        .dout(new_Jinkela_wire_3546)
    );

    bfr new_Jinkela_buffer_4756 (
        .din(new_Jinkela_wire_5683),
        .dout(new_Jinkela_wire_5684)
    );

    bfr new_Jinkela_buffer_7271 (
        .din(n_1358_),
        .dout(new_Jinkela_wire_9026)
    );

    bfr new_Jinkela_buffer_3048 (
        .din(new_Jinkela_wire_3477),
        .dout(new_Jinkela_wire_3478)
    );

    bfr new_Jinkela_buffer_7323 (
        .din(new_net_2495),
        .dout(new_Jinkela_wire_9093)
    );

    bfr new_Jinkela_buffer_4711 (
        .din(new_Jinkela_wire_5616),
        .dout(new_Jinkela_wire_5617)
    );

    spl2 new_Jinkela_splitter_709 (
        .a(n_0249_),
        .b(new_Jinkela_wire_9091),
        .c(new_Jinkela_wire_9092)
    );

    bfr new_Jinkela_buffer_7272 (
        .din(new_Jinkela_wire_9026),
        .dout(new_Jinkela_wire_9027)
    );

    bfr new_Jinkela_buffer_3118 (
        .din(N192),
        .dout(new_Jinkela_wire_3555)
    );

    bfr new_Jinkela_buffer_4736 (
        .din(new_Jinkela_wire_5655),
        .dout(new_Jinkela_wire_5656)
    );

    bfr new_Jinkela_buffer_3049 (
        .din(new_Jinkela_wire_3478),
        .dout(new_Jinkela_wire_3479)
    );

    spl2 new_Jinkela_splitter_708 (
        .a(n_1114_),
        .b(new_Jinkela_wire_9089),
        .c(new_Jinkela_wire_9090)
    );

    bfr new_Jinkela_buffer_4712 (
        .din(new_Jinkela_wire_5617),
        .dout(new_Jinkela_wire_5618)
    );

    bfr new_Jinkela_buffer_7273 (
        .din(new_Jinkela_wire_9027),
        .dout(new_Jinkela_wire_9028)
    );

    bfr new_Jinkela_buffer_3112 (
        .din(new_Jinkela_wire_3548),
        .dout(new_Jinkela_wire_3549)
    );

    bfr new_Jinkela_buffer_4932 (
        .din(n_0610_),
        .dout(new_Jinkela_wire_5872)
    );

    bfr new_Jinkela_buffer_3050 (
        .din(new_Jinkela_wire_3479),
        .dout(new_Jinkela_wire_3480)
    );

    bfr new_Jinkela_buffer_4802 (
        .din(new_Jinkela_wire_5733),
        .dout(new_Jinkela_wire_5734)
    );

    bfr new_Jinkela_buffer_4713 (
        .din(new_Jinkela_wire_5618),
        .dout(new_Jinkela_wire_5619)
    );

    bfr new_Jinkela_buffer_7274 (
        .din(new_Jinkela_wire_9028),
        .dout(new_Jinkela_wire_9029)
    );

    bfr new_Jinkela_buffer_3115 (
        .din(new_Jinkela_wire_3551),
        .dout(new_Jinkela_wire_3552)
    );

    bfr new_Jinkela_buffer_4737 (
        .din(new_Jinkela_wire_5656),
        .dout(new_Jinkela_wire_5657)
    );

    bfr new_Jinkela_buffer_7324 (
        .din(new_Jinkela_wire_9093),
        .dout(new_Jinkela_wire_9094)
    );

    bfr new_Jinkela_buffer_3051 (
        .din(new_Jinkela_wire_3480),
        .dout(new_Jinkela_wire_3481)
    );

    bfr new_Jinkela_buffer_7280 (
        .din(new_Jinkela_wire_9041),
        .dout(new_Jinkela_wire_9042)
    );

    bfr new_Jinkela_buffer_4714 (
        .din(new_Jinkela_wire_5619),
        .dout(new_Jinkela_wire_5620)
    );

    bfr new_Jinkela_buffer_7275 (
        .din(new_Jinkela_wire_9029),
        .dout(new_Jinkela_wire_9030)
    );

    bfr new_Jinkela_buffer_3113 (
        .din(new_Jinkela_wire_3549),
        .dout(new_Jinkela_wire_3550)
    );

    bfr new_Jinkela_buffer_4757 (
        .din(new_Jinkela_wire_5684),
        .dout(new_Jinkela_wire_5685)
    );

    bfr new_Jinkela_buffer_3052 (
        .din(new_Jinkela_wire_3481),
        .dout(new_Jinkela_wire_3482)
    );

    bfr new_Jinkela_buffer_7340 (
        .din(n_1288_),
        .dout(new_Jinkela_wire_9113)
    );

    bfr new_Jinkela_buffer_4715 (
        .din(new_Jinkela_wire_5620),
        .dout(new_Jinkela_wire_5621)
    );

    bfr new_Jinkela_buffer_7276 (
        .din(new_Jinkela_wire_9030),
        .dout(new_Jinkela_wire_9031)
    );

    bfr new_Jinkela_buffer_3122 (
        .din(N63),
        .dout(new_Jinkela_wire_3559)
    );

    bfr new_Jinkela_buffer_4738 (
        .din(new_Jinkela_wire_5657),
        .dout(new_Jinkela_wire_5658)
    );

    bfr new_Jinkela_buffer_3053 (
        .din(new_Jinkela_wire_3482),
        .dout(new_Jinkela_wire_3483)
    );

    spl2 new_Jinkela_splitter_706 (
        .a(new_Jinkela_wire_9042),
        .b(new_Jinkela_wire_9043),
        .c(new_Jinkela_wire_9044)
    );

    bfr new_Jinkela_buffer_4716 (
        .din(new_Jinkela_wire_5621),
        .dout(new_Jinkela_wire_5622)
    );

    bfr new_Jinkela_buffer_7277 (
        .din(new_Jinkela_wire_9031),
        .dout(new_Jinkela_wire_9032)
    );

    bfr new_Jinkela_buffer_3116 (
        .din(new_Jinkela_wire_3552),
        .dout(new_Jinkela_wire_3553)
    );

    bfr new_Jinkela_buffer_3054 (
        .din(new_Jinkela_wire_3483),
        .dout(new_Jinkela_wire_3484)
    );

    bfr new_Jinkela_buffer_4717 (
        .din(new_Jinkela_wire_5622),
        .dout(new_Jinkela_wire_5623)
    );

    spl2 new_Jinkela_splitter_703 (
        .a(new_Jinkela_wire_9032),
        .b(new_Jinkela_wire_9033),
        .c(new_Jinkela_wire_9034)
    );

    bfr new_Jinkela_buffer_3119 (
        .din(new_Jinkela_wire_3555),
        .dout(new_Jinkela_wire_3556)
    );

    bfr new_Jinkela_buffer_4739 (
        .din(new_Jinkela_wire_5658),
        .dout(new_Jinkela_wire_5659)
    );

    bfr new_Jinkela_buffer_7278 (
        .din(new_Jinkela_wire_9034),
        .dout(new_Jinkela_wire_9035)
    );

    bfr new_Jinkela_buffer_3055 (
        .din(new_Jinkela_wire_3484),
        .dout(new_Jinkela_wire_3485)
    );

    bfr new_Jinkela_buffer_4718 (
        .din(new_Jinkela_wire_5623),
        .dout(new_Jinkela_wire_5624)
    );

    bfr new_Jinkela_buffer_7281 (
        .din(new_Jinkela_wire_9044),
        .dout(new_Jinkela_wire_9045)
    );

    bfr new_Jinkela_buffer_3117 (
        .din(new_Jinkela_wire_3553),
        .dout(new_Jinkela_wire_3554)
    );

    bfr new_Jinkela_buffer_4758 (
        .din(new_Jinkela_wire_5685),
        .dout(new_Jinkela_wire_5686)
    );

    bfr new_Jinkela_buffer_3056 (
        .din(new_Jinkela_wire_3485),
        .dout(new_Jinkela_wire_3486)
    );

    spl3L new_Jinkela_splitter_710 (
        .a(n_0063_),
        .d(new_Jinkela_wire_9110),
        .b(new_Jinkela_wire_9111),
        .c(new_Jinkela_wire_9112)
    );

    bfr new_Jinkela_buffer_4719 (
        .din(new_Jinkela_wire_5624),
        .dout(new_Jinkela_wire_5625)
    );

    bfr new_Jinkela_buffer_7279 (
        .din(new_Jinkela_wire_9035),
        .dout(new_Jinkela_wire_9036)
    );

    spl2 new_Jinkela_splitter_149 (
        .a(n_0045_),
        .b(new_Jinkela_wire_3563),
        .c(new_Jinkela_wire_3564)
    );

    bfr new_Jinkela_buffer_4740 (
        .din(new_Jinkela_wire_5659),
        .dout(new_Jinkela_wire_5660)
    );

    bfr new_Jinkela_buffer_3057 (
        .din(new_Jinkela_wire_3486),
        .dout(new_Jinkela_wire_3487)
    );

    bfr new_Jinkela_buffer_4720 (
        .din(new_Jinkela_wire_5625),
        .dout(new_Jinkela_wire_5626)
    );

    bfr new_Jinkela_buffer_7282 (
        .din(new_Jinkela_wire_9045),
        .dout(new_Jinkela_wire_9046)
    );

    bfr new_Jinkela_buffer_3138 (
        .din(n_0888_),
        .dout(new_Jinkela_wire_3577)
    );

    bfr new_Jinkela_buffer_3120 (
        .din(new_Jinkela_wire_3556),
        .dout(new_Jinkela_wire_3557)
    );

    bfr new_Jinkela_buffer_3058 (
        .din(new_Jinkela_wire_3487),
        .dout(new_Jinkela_wire_3488)
    );

    bfr new_Jinkela_buffer_4803 (
        .din(new_Jinkela_wire_5734),
        .dout(new_Jinkela_wire_5735)
    );

    bfr new_Jinkela_buffer_7325 (
        .din(new_Jinkela_wire_9094),
        .dout(new_Jinkela_wire_9095)
    );

    bfr new_Jinkela_buffer_4721 (
        .din(new_Jinkela_wire_5626),
        .dout(new_Jinkela_wire_5627)
    );

    bfr new_Jinkela_buffer_7283 (
        .din(new_Jinkela_wire_9046),
        .dout(new_Jinkela_wire_9047)
    );

    bfr new_Jinkela_buffer_6419 (
        .din(n_0281_),
        .dout(new_Jinkela_wire_7837)
    );

    bfr new_Jinkela_buffer_6380 (
        .din(new_Jinkela_wire_7785),
        .dout(new_Jinkela_wire_7786)
    );

    spl2 new_Jinkela_splitter_555 (
        .a(new_Jinkela_wire_7811),
        .b(new_Jinkela_wire_7812),
        .c(new_Jinkela_wire_7813)
    );

    bfr new_Jinkela_buffer_6381 (
        .din(new_Jinkela_wire_7786),
        .dout(new_Jinkela_wire_7787)
    );

    bfr new_Jinkela_buffer_6404 (
        .din(new_Jinkela_wire_7813),
        .dout(new_Jinkela_wire_7814)
    );

    bfr new_Jinkela_buffer_6382 (
        .din(new_Jinkela_wire_7787),
        .dout(new_Jinkela_wire_7788)
    );

    bfr new_Jinkela_buffer_6383 (
        .din(new_Jinkela_wire_7788),
        .dout(new_Jinkela_wire_7789)
    );

    bfr new_Jinkela_buffer_6413 (
        .din(new_Jinkela_wire_7826),
        .dout(new_Jinkela_wire_7827)
    );

    bfr new_Jinkela_buffer_6384 (
        .din(new_Jinkela_wire_7789),
        .dout(new_Jinkela_wire_7790)
    );

    bfr new_Jinkela_buffer_6405 (
        .din(new_Jinkela_wire_7814),
        .dout(new_Jinkela_wire_7815)
    );

    bfr new_Jinkela_buffer_6385 (
        .din(new_Jinkela_wire_7790),
        .dout(new_Jinkela_wire_7791)
    );

    bfr new_Jinkela_buffer_6416 (
        .din(new_Jinkela_wire_7829),
        .dout(new_Jinkela_wire_7830)
    );

    bfr new_Jinkela_buffer_6386 (
        .din(new_Jinkela_wire_7791),
        .dout(new_Jinkela_wire_7792)
    );

    bfr new_Jinkela_buffer_6406 (
        .din(new_Jinkela_wire_7815),
        .dout(new_Jinkela_wire_7816)
    );

    bfr new_Jinkela_buffer_6387 (
        .din(new_Jinkela_wire_7792),
        .dout(new_Jinkela_wire_7793)
    );

    bfr new_Jinkela_buffer_6414 (
        .din(new_Jinkela_wire_7827),
        .dout(new_Jinkela_wire_7828)
    );

    bfr new_Jinkela_buffer_6388 (
        .din(new_Jinkela_wire_7793),
        .dout(new_Jinkela_wire_7794)
    );

    bfr new_Jinkela_buffer_6407 (
        .din(new_Jinkela_wire_7816),
        .dout(new_Jinkela_wire_7817)
    );

    bfr new_Jinkela_buffer_6389 (
        .din(new_Jinkela_wire_7794),
        .dout(new_Jinkela_wire_7795)
    );

    bfr new_Jinkela_buffer_6390 (
        .din(new_Jinkela_wire_7795),
        .dout(new_Jinkela_wire_7796)
    );

    bfr new_Jinkela_buffer_6408 (
        .din(new_Jinkela_wire_7817),
        .dout(new_Jinkela_wire_7818)
    );

    bfr new_Jinkela_buffer_6391 (
        .din(new_Jinkela_wire_7796),
        .dout(new_Jinkela_wire_7797)
    );

    bfr new_Jinkela_buffer_6417 (
        .din(new_Jinkela_wire_7830),
        .dout(new_Jinkela_wire_7831)
    );

    bfr new_Jinkela_buffer_6392 (
        .din(new_Jinkela_wire_7797),
        .dout(new_Jinkela_wire_7798)
    );

    bfr new_Jinkela_buffer_6409 (
        .din(new_Jinkela_wire_7818),
        .dout(new_Jinkela_wire_7819)
    );

    bfr new_Jinkela_buffer_6393 (
        .din(new_Jinkela_wire_7798),
        .dout(new_Jinkela_wire_7799)
    );

    bfr new_Jinkela_buffer_6418 (
        .din(new_Jinkela_wire_7835),
        .dout(new_Jinkela_wire_7836)
    );

    spl2 new_Jinkela_splitter_560 (
        .a(n_1327_),
        .b(new_Jinkela_wire_7838),
        .c(new_Jinkela_wire_7839)
    );

    bfr new_Jinkela_buffer_6394 (
        .din(new_Jinkela_wire_7799),
        .dout(new_Jinkela_wire_7800)
    );

    spl2 new_Jinkela_splitter_558 (
        .a(new_Jinkela_wire_7831),
        .b(new_Jinkela_wire_7832),
        .c(new_Jinkela_wire_7833)
    );

    bfr new_Jinkela_buffer_6395 (
        .din(new_Jinkela_wire_7800),
        .dout(new_Jinkela_wire_7801)
    );

    bfr new_Jinkela_buffer_6420 (
        .din(n_0282_),
        .dout(new_Jinkela_wire_7845)
    );

    bfr new_Jinkela_buffer_6396 (
        .din(new_Jinkela_wire_7801),
        .dout(new_Jinkela_wire_7802)
    );

    spl2 new_Jinkela_splitter_561 (
        .a(n_0095_),
        .b(new_Jinkela_wire_7840),
        .c(new_Jinkela_wire_7841)
    );

    bfr new_Jinkela_buffer_6424 (
        .din(n_0265_),
        .dout(new_Jinkela_wire_7851)
    );

    bfr new_Jinkela_buffer_6397 (
        .din(new_Jinkela_wire_7802),
        .dout(new_Jinkela_wire_7803)
    );

    spl3L new_Jinkela_splitter_562 (
        .a(n_1137_),
        .d(new_Jinkela_wire_7842),
        .b(new_Jinkela_wire_7843),
        .c(new_Jinkela_wire_7844)
    );

    spl2 new_Jinkela_splitter_563 (
        .a(n_0688_),
        .b(new_Jinkela_wire_7849),
        .c(new_Jinkela_wire_7850)
    );

    bfr new_Jinkela_buffer_6421 (
        .din(new_Jinkela_wire_7845),
        .dout(new_Jinkela_wire_7846)
    );

    bfr new_Jinkela_buffer_6425 (
        .din(new_net_12),
        .dout(new_Jinkela_wire_7852)
    );

    bfr new_Jinkela_buffer_6487 (
        .din(n_0615_),
        .dout(new_Jinkela_wire_7916)
    );

    bfr new_Jinkela_buffer_6422 (
        .din(new_Jinkela_wire_7846),
        .dout(new_Jinkela_wire_7847)
    );

    bfr new_Jinkela_buffer_3881 (
        .din(new_Jinkela_wire_4551),
        .dout(new_Jinkela_wire_4552)
    );

    spl2 new_Jinkela_splitter_428 (
        .a(new_Jinkela_wire_6669),
        .b(new_Jinkela_wire_6670),
        .c(new_Jinkela_wire_6671)
    );

    spl2 new_Jinkela_splitter_246 (
        .a(n_0208_),
        .b(new_Jinkela_wire_4631),
        .c(new_Jinkela_wire_4632)
    );

    spl2 new_Jinkela_splitter_247 (
        .a(n_1343_),
        .b(new_Jinkela_wire_4633),
        .c(new_Jinkela_wire_4634)
    );

    bfr new_Jinkela_buffer_5579 (
        .din(new_Jinkela_wire_6689),
        .dout(new_Jinkela_wire_6690)
    );

    bfr new_Jinkela_buffer_3882 (
        .din(new_Jinkela_wire_4552),
        .dout(new_Jinkela_wire_4553)
    );

    bfr new_Jinkela_buffer_5628 (
        .din(new_Jinkela_wire_6748),
        .dout(new_Jinkela_wire_6749)
    );

    bfr new_Jinkela_buffer_3903 (
        .din(new_Jinkela_wire_4573),
        .dout(new_Jinkela_wire_4574)
    );

    bfr new_Jinkela_buffer_5602 (
        .din(new_Jinkela_wire_6716),
        .dout(new_Jinkela_wire_6717)
    );

    bfr new_Jinkela_buffer_3883 (
        .din(new_Jinkela_wire_4553),
        .dout(new_Jinkela_wire_4554)
    );

    bfr new_Jinkela_buffer_5580 (
        .din(new_Jinkela_wire_6690),
        .dout(new_Jinkela_wire_6691)
    );

    spl4L new_Jinkela_splitter_249 (
        .a(n_0851_),
        .d(new_Jinkela_wire_4645),
        .b(new_Jinkela_wire_4646),
        .e(new_Jinkela_wire_4647),
        .c(new_Jinkela_wire_4648)
    );

    spl2 new_Jinkela_splitter_436 (
        .a(n_0674_),
        .b(new_Jinkela_wire_6768),
        .c(new_Jinkela_wire_6769)
    );

    bfr new_Jinkela_buffer_3884 (
        .din(new_Jinkela_wire_4554),
        .dout(new_Jinkela_wire_4555)
    );

    bfr new_Jinkela_buffer_5581 (
        .din(new_Jinkela_wire_6691),
        .dout(new_Jinkela_wire_6692)
    );

    bfr new_Jinkela_buffer_3904 (
        .din(new_Jinkela_wire_4574),
        .dout(new_Jinkela_wire_4575)
    );

    bfr new_Jinkela_buffer_5603 (
        .din(new_Jinkela_wire_6717),
        .dout(new_Jinkela_wire_6718)
    );

    bfr new_Jinkela_buffer_3885 (
        .din(new_Jinkela_wire_4555),
        .dout(new_Jinkela_wire_4556)
    );

    bfr new_Jinkela_buffer_5582 (
        .din(new_Jinkela_wire_6692),
        .dout(new_Jinkela_wire_6693)
    );

    bfr new_Jinkela_buffer_5629 (
        .din(new_Jinkela_wire_6749),
        .dout(new_Jinkela_wire_6750)
    );

    bfr new_Jinkela_buffer_3886 (
        .din(new_Jinkela_wire_4556),
        .dout(new_Jinkela_wire_4557)
    );

    bfr new_Jinkela_buffer_5583 (
        .din(new_Jinkela_wire_6693),
        .dout(new_Jinkela_wire_6694)
    );

    bfr new_Jinkela_buffer_3905 (
        .din(new_Jinkela_wire_4575),
        .dout(new_Jinkela_wire_4576)
    );

    bfr new_Jinkela_buffer_5604 (
        .din(new_Jinkela_wire_6718),
        .dout(new_Jinkela_wire_6719)
    );

    bfr new_Jinkela_buffer_3887 (
        .din(new_Jinkela_wire_4557),
        .dout(new_Jinkela_wire_4558)
    );

    bfr new_Jinkela_buffer_5584 (
        .din(new_Jinkela_wire_6694),
        .dout(new_Jinkela_wire_6695)
    );

    spl2 new_Jinkela_splitter_248 (
        .a(n_0532_),
        .b(new_Jinkela_wire_4643),
        .c(new_Jinkela_wire_4644)
    );

    bfr new_Jinkela_buffer_3958 (
        .din(new_Jinkela_wire_4634),
        .dout(new_Jinkela_wire_4635)
    );

    bfr new_Jinkela_buffer_3888 (
        .din(new_Jinkela_wire_4558),
        .dout(new_Jinkela_wire_4559)
    );

    bfr new_Jinkela_buffer_5585 (
        .din(new_Jinkela_wire_6695),
        .dout(new_Jinkela_wire_6696)
    );

    bfr new_Jinkela_buffer_3906 (
        .din(new_Jinkela_wire_4576),
        .dout(new_Jinkela_wire_4577)
    );

    bfr new_Jinkela_buffer_5645 (
        .din(new_Jinkela_wire_6769),
        .dout(new_Jinkela_wire_6770)
    );

    bfr new_Jinkela_buffer_5605 (
        .din(new_Jinkela_wire_6719),
        .dout(new_Jinkela_wire_6720)
    );

    bfr new_Jinkela_buffer_3889 (
        .din(new_Jinkela_wire_4559),
        .dout(new_Jinkela_wire_4560)
    );

    bfr new_Jinkela_buffer_5586 (
        .din(new_Jinkela_wire_6696),
        .dout(new_Jinkela_wire_6697)
    );

    spl2 new_Jinkela_splitter_251 (
        .a(n_1170_),
        .b(new_Jinkela_wire_4652),
        .c(new_Jinkela_wire_4653)
    );

    bfr new_Jinkela_buffer_5630 (
        .din(new_Jinkela_wire_6750),
        .dout(new_Jinkela_wire_6751)
    );

    bfr new_Jinkela_buffer_3890 (
        .din(new_Jinkela_wire_4560),
        .dout(new_Jinkela_wire_4561)
    );

    bfr new_Jinkela_buffer_5587 (
        .din(new_Jinkela_wire_6697),
        .dout(new_Jinkela_wire_6698)
    );

    bfr new_Jinkela_buffer_3907 (
        .din(new_Jinkela_wire_4577),
        .dout(new_Jinkela_wire_4578)
    );

    bfr new_Jinkela_buffer_5606 (
        .din(new_Jinkela_wire_6720),
        .dout(new_Jinkela_wire_6721)
    );

    bfr new_Jinkela_buffer_3891 (
        .din(new_Jinkela_wire_4561),
        .dout(new_Jinkela_wire_4562)
    );

    bfr new_Jinkela_buffer_5588 (
        .din(new_Jinkela_wire_6698),
        .dout(new_Jinkela_wire_6699)
    );

    bfr new_Jinkela_buffer_3959 (
        .din(new_Jinkela_wire_4635),
        .dout(new_Jinkela_wire_4636)
    );

    bfr new_Jinkela_buffer_3892 (
        .din(new_Jinkela_wire_4562),
        .dout(new_Jinkela_wire_4563)
    );

    bfr new_Jinkela_buffer_5589 (
        .din(new_Jinkela_wire_6699),
        .dout(new_Jinkela_wire_6700)
    );

    bfr new_Jinkela_buffer_3908 (
        .din(new_Jinkela_wire_4578),
        .dout(new_Jinkela_wire_4579)
    );

    bfr new_Jinkela_buffer_5607 (
        .din(new_Jinkela_wire_6721),
        .dout(new_Jinkela_wire_6722)
    );

    bfr new_Jinkela_buffer_3893 (
        .din(new_Jinkela_wire_4563),
        .dout(new_Jinkela_wire_4564)
    );

    bfr new_Jinkela_buffer_5590 (
        .din(new_Jinkela_wire_6700),
        .dout(new_Jinkela_wire_6701)
    );

    bfr new_Jinkela_buffer_5631 (
        .din(new_Jinkela_wire_6751),
        .dout(new_Jinkela_wire_6752)
    );

    bfr new_Jinkela_buffer_3894 (
        .din(new_Jinkela_wire_4564),
        .dout(new_Jinkela_wire_4565)
    );

    bfr new_Jinkela_buffer_5591 (
        .din(new_Jinkela_wire_6701),
        .dout(new_Jinkela_wire_6702)
    );

    bfr new_Jinkela_buffer_3909 (
        .din(new_Jinkela_wire_4579),
        .dout(new_Jinkela_wire_4580)
    );

    bfr new_Jinkela_buffer_5608 (
        .din(new_Jinkela_wire_6722),
        .dout(new_Jinkela_wire_6723)
    );

    bfr new_Jinkela_buffer_3895 (
        .din(new_Jinkela_wire_4565),
        .dout(new_Jinkela_wire_4566)
    );

    bfr new_Jinkela_buffer_5592 (
        .din(new_Jinkela_wire_6702),
        .dout(new_Jinkela_wire_6703)
    );

    bfr new_Jinkela_buffer_3966 (
        .din(n_0434_),
        .dout(new_Jinkela_wire_4649)
    );

    bfr new_Jinkela_buffer_3960 (
        .din(new_Jinkela_wire_4636),
        .dout(new_Jinkela_wire_4637)
    );

    spl2 new_Jinkela_splitter_440 (
        .a(n_0484_),
        .b(new_Jinkela_wire_6788),
        .c(new_Jinkela_wire_6789)
    );

    bfr new_Jinkela_buffer_3896 (
        .din(new_Jinkela_wire_4566),
        .dout(new_Jinkela_wire_4567)
    );

    bfr new_Jinkela_buffer_5593 (
        .din(new_Jinkela_wire_6703),
        .dout(new_Jinkela_wire_6704)
    );

    bfr new_Jinkela_buffer_3910 (
        .din(new_Jinkela_wire_4580),
        .dout(new_Jinkela_wire_4581)
    );

    bfr new_Jinkela_buffer_5656 (
        .din(n_0612_),
        .dout(new_Jinkela_wire_6790)
    );

    bfr new_Jinkela_buffer_5609 (
        .din(new_Jinkela_wire_6723),
        .dout(new_Jinkela_wire_6724)
    );

    bfr new_Jinkela_buffer_3897 (
        .din(new_Jinkela_wire_4567),
        .dout(new_Jinkela_wire_4568)
    );

    bfr new_Jinkela_buffer_5594 (
        .din(new_Jinkela_wire_6704),
        .dout(new_Jinkela_wire_6705)
    );

    spl2 new_Jinkela_splitter_250 (
        .a(new_Jinkela_wire_4649),
        .b(new_Jinkela_wire_4650),
        .c(new_Jinkela_wire_4651)
    );

    bfr new_Jinkela_buffer_5632 (
        .din(new_Jinkela_wire_6752),
        .dout(new_Jinkela_wire_6753)
    );

    bfr new_Jinkela_buffer_3898 (
        .din(new_Jinkela_wire_4568),
        .dout(new_Jinkela_wire_4569)
    );

    bfr new_Jinkela_buffer_5610 (
        .din(new_Jinkela_wire_6724),
        .dout(new_Jinkela_wire_6725)
    );

    bfr new_Jinkela_buffer_3911 (
        .din(new_Jinkela_wire_4581),
        .dout(new_Jinkela_wire_4582)
    );

    bfr new_Jinkela_buffer_3961 (
        .din(new_Jinkela_wire_4637),
        .dout(new_Jinkela_wire_4638)
    );

    bfr new_Jinkela_buffer_5646 (
        .din(new_Jinkela_wire_6770),
        .dout(new_Jinkela_wire_6771)
    );

    bfr new_Jinkela_buffer_5611 (
        .din(new_Jinkela_wire_6725),
        .dout(new_Jinkela_wire_6726)
    );

    bfr new_Jinkela_buffer_3912 (
        .din(new_Jinkela_wire_4582),
        .dout(new_Jinkela_wire_4583)
    );

    bfr new_Jinkela_buffer_5633 (
        .din(new_Jinkela_wire_6753),
        .dout(new_Jinkela_wire_6754)
    );

    spl2 new_Jinkela_splitter_252 (
        .a(n_1087_),
        .b(new_Jinkela_wire_4654),
        .c(new_Jinkela_wire_4655)
    );

    bfr new_Jinkela_buffer_5612 (
        .din(new_Jinkela_wire_6726),
        .dout(new_Jinkela_wire_6727)
    );

    bfr new_Jinkela_buffer_3913 (
        .din(new_Jinkela_wire_4583),
        .dout(new_Jinkela_wire_4584)
    );

    bfr new_Jinkela_buffer_3962 (
        .din(new_Jinkela_wire_4638),
        .dout(new_Jinkela_wire_4639)
    );

    spl3L new_Jinkela_splitter_438 (
        .a(n_0960_),
        .d(new_Jinkela_wire_6783),
        .b(new_Jinkela_wire_6784),
        .c(new_Jinkela_wire_6785)
    );

    bfr new_Jinkela_buffer_5613 (
        .din(new_Jinkela_wire_6727),
        .dout(new_Jinkela_wire_6728)
    );

    bfr new_Jinkela_buffer_3914 (
        .din(new_Jinkela_wire_4584),
        .dout(new_Jinkela_wire_4585)
    );

    bfr new_Jinkela_buffer_2134 (
        .din(new_Jinkela_wire_2508),
        .dout(new_Jinkela_wire_2509)
    );

    and_ii n_2367_ (
        .a(new_Jinkela_wire_8391),
        .b(n_0238_),
        .c(n_0242_)
    );

    and_bb n_2368_ (
        .a(new_Jinkela_wire_4872),
        .b(new_Jinkela_wire_5285),
        .c(n_0243_)
    );

    bfr new_Jinkela_buffer_2189 (
        .din(new_Jinkela_wire_2567),
        .dout(new_Jinkela_wire_2568)
    );

    bfr new_Jinkela_buffer_2135 (
        .din(new_Jinkela_wire_2509),
        .dout(new_Jinkela_wire_2510)
    );

    and_ii n_2369_ (
        .a(new_Jinkela_wire_3725),
        .b(new_Jinkela_wire_3953),
        .c(n_0244_)
    );

    and_ii n_2370_ (
        .a(new_Jinkela_wire_4544),
        .b(new_Jinkela_wire_8706),
        .c(n_0245_)
    );

    bfr new_Jinkela_buffer_2207 (
        .din(new_Jinkela_wire_2589),
        .dout(new_Jinkela_wire_2590)
    );

    bfr new_Jinkela_buffer_2136 (
        .din(new_Jinkela_wire_2510),
        .dout(new_Jinkela_wire_2511)
    );

    and_ii n_2371_ (
        .a(new_Jinkela_wire_4874),
        .b(new_Jinkela_wire_5286),
        .c(n_0246_)
    );

    and_bb n_2372_ (
        .a(new_Jinkela_wire_3723),
        .b(new_Jinkela_wire_3952),
        .c(n_0247_)
    );

    bfr new_Jinkela_buffer_2137 (
        .din(new_Jinkela_wire_2511),
        .dout(new_Jinkela_wire_2512)
    );

    or_bb n_2373_ (
        .a(new_Jinkela_wire_6814),
        .b(new_Jinkela_wire_9533),
        .c(n_0248_)
    );

    bfr new_Jinkela_buffer_2273 (
        .din(new_Jinkela_wire_2659),
        .dout(new_Jinkela_wire_2660)
    );

    and_bi n_2374_ (
        .a(n_0245_),
        .b(n_0248_),
        .c(n_0249_)
    );

    bfr new_Jinkela_buffer_2190 (
        .din(new_Jinkela_wire_2568),
        .dout(new_Jinkela_wire_2569)
    );

    bfr new_Jinkela_buffer_2138 (
        .din(new_Jinkela_wire_2512),
        .dout(new_Jinkela_wire_2513)
    );

    and_ii n_2375_ (
        .a(new_Jinkela_wire_5367),
        .b(new_Jinkela_wire_7080),
        .c(n_0250_)
    );

    and_ii n_2376_ (
        .a(new_Jinkela_wire_10526),
        .b(new_Jinkela_wire_8169),
        .c(n_0251_)
    );

    bfr new_Jinkela_buffer_2139 (
        .din(new_Jinkela_wire_2513),
        .dout(new_Jinkela_wire_2514)
    );

    and_ii n_2377_ (
        .a(n_0251_),
        .b(n_0250_),
        .c(n_0252_)
    );

    bfr new_Jinkela_buffer_2209 (
        .din(new_Jinkela_wire_2593),
        .dout(new_Jinkela_wire_2594)
    );

    and_bb n_2378_ (
        .a(new_Jinkela_wire_5365),
        .b(new_Jinkela_wire_7079),
        .c(n_0253_)
    );

    bfr new_Jinkela_buffer_2191 (
        .din(new_Jinkela_wire_2569),
        .dout(new_Jinkela_wire_2570)
    );

    bfr new_Jinkela_buffer_2140 (
        .din(new_Jinkela_wire_2514),
        .dout(new_Jinkela_wire_2515)
    );

    and_bb n_2379_ (
        .a(new_Jinkela_wire_10523),
        .b(new_Jinkela_wire_8168),
        .c(n_0254_)
    );

    and_ii n_2380_ (
        .a(new_Jinkela_wire_8995),
        .b(new_Jinkela_wire_7086),
        .c(n_0255_)
    );

    bfr new_Jinkela_buffer_2141 (
        .din(new_Jinkela_wire_2515),
        .dout(new_Jinkela_wire_2516)
    );

    and_bb n_2381_ (
        .a(n_0255_),
        .b(new_Jinkela_wire_3943),
        .c(n_0256_)
    );

    or_ii n_2382_ (
        .a(new_Jinkela_wire_4629),
        .b(new_Jinkela_wire_9092),
        .c(n_0257_)
    );

    bfr new_Jinkela_buffer_2192 (
        .din(new_Jinkela_wire_2570),
        .dout(new_Jinkela_wire_2571)
    );

    bfr new_Jinkela_buffer_2142 (
        .din(new_Jinkela_wire_2516),
        .dout(new_Jinkela_wire_2517)
    );

    and_ii n_2383_ (
        .a(new_Jinkela_wire_7369),
        .b(n_0242_),
        .c(n_0258_)
    );

    or_bb n_2384_ (
        .a(new_Jinkela_wire_7088),
        .b(new_Jinkela_wire_3942),
        .c(n_0259_)
    );

    bfr new_Jinkela_buffer_2412 (
        .din(N159),
        .dout(new_Jinkela_wire_2809)
    );

    bfr new_Jinkela_buffer_2143 (
        .din(new_Jinkela_wire_2517),
        .dout(new_Jinkela_wire_2518)
    );

    and_bi n_2385_ (
        .a(new_Jinkela_wire_9091),
        .b(new_Jinkela_wire_9344),
        .c(n_0260_)
    );

    spl2 new_Jinkela_splitter_128 (
        .a(new_Jinkela_wire_2594),
        .b(new_Jinkela_wire_2595),
        .c(new_Jinkela_wire_2596)
    );

    and_bi n_2386_ (
        .a(new_Jinkela_wire_4543),
        .b(new_Jinkela_wire_8705),
        .c(n_0261_)
    );

    bfr new_Jinkela_buffer_2193 (
        .din(new_Jinkela_wire_2571),
        .dout(new_Jinkela_wire_2572)
    );

    bfr new_Jinkela_buffer_2144 (
        .din(new_Jinkela_wire_2518),
        .dout(new_Jinkela_wire_2519)
    );

    or_bb n_2387_ (
        .a(n_0261_),
        .b(new_Jinkela_wire_9535),
        .c(n_0262_)
    );

    or_bb n_2388_ (
        .a(new_Jinkela_wire_5165),
        .b(n_0260_),
        .c(n_0263_)
    );

    bfr new_Jinkela_buffer_2145 (
        .din(new_Jinkela_wire_2519),
        .dout(new_Jinkela_wire_2520)
    );

    and_ii n_2389_ (
        .a(new_Jinkela_wire_8714),
        .b(n_0258_),
        .c(n_0264_)
    );

    bfr new_Jinkela_buffer_2210 (
        .din(new_Jinkela_wire_2596),
        .dout(new_Jinkela_wire_2597)
    );

    and_bi n_2390_ (
        .a(new_Jinkela_wire_6106),
        .b(new_Jinkela_wire_8750),
        .c(n_0265_)
    );

    spl2 new_Jinkela_splitter_125 (
        .a(new_Jinkela_wire_2572),
        .b(new_Jinkela_wire_2573),
        .c(new_Jinkela_wire_2574)
    );

    bfr new_Jinkela_buffer_2146 (
        .din(new_Jinkela_wire_2520),
        .dout(new_Jinkela_wire_2521)
    );

    and_ii n_2391_ (
        .a(new_Jinkela_wire_7327),
        .b(new_Jinkela_wire_3586),
        .c(n_0266_)
    );

    or_bb n_2392_ (
        .a(n_0266_),
        .b(new_Jinkela_wire_7851),
        .c(n_0267_)
    );

    bfr new_Jinkela_buffer_2194 (
        .din(new_Jinkela_wire_2574),
        .dout(new_Jinkela_wire_2575)
    );

    bfr new_Jinkela_buffer_2147 (
        .din(new_Jinkela_wire_2521),
        .dout(new_Jinkela_wire_2522)
    );

    and_bi n_2393_ (
        .a(new_Jinkela_wire_8749),
        .b(new_Jinkela_wire_6105),
        .c(n_0268_)
    );

    bfr new_Jinkela_buffer_6784 (
        .din(new_Jinkela_wire_8359),
        .dout(new_Jinkela_wire_8360)
    );

    and_bb n_2394_ (
        .a(new_Jinkela_wire_7329),
        .b(new_Jinkela_wire_3587),
        .c(n_0269_)
    );

    bfr new_Jinkela_buffer_2148 (
        .din(new_Jinkela_wire_2522),
        .dout(new_Jinkela_wire_2523)
    );

    or_bb n_2395_ (
        .a(n_0269_),
        .b(new_Jinkela_wire_7923),
        .c(n_0270_)
    );

    bfr new_Jinkela_buffer_2274 (
        .din(new_Jinkela_wire_2660),
        .dout(new_Jinkela_wire_2661)
    );

    and_ii n_2396_ (
        .a(new_Jinkela_wire_4526),
        .b(new_Jinkela_wire_10136),
        .c(n_0271_)
    );

    bfr new_Jinkela_buffer_2149 (
        .din(new_Jinkela_wire_2523),
        .dout(new_Jinkela_wire_2524)
    );

    and_ii n_2397_ (
        .a(new_Jinkela_wire_9381),
        .b(new_Jinkela_wire_8316),
        .c(n_0272_)
    );

    bfr new_Jinkela_buffer_2340 (
        .din(N234),
        .dout(new_Jinkela_wire_2732)
    );

    and_ii n_2398_ (
        .a(new_Jinkela_wire_4971),
        .b(new_Jinkela_wire_10224),
        .c(n_0273_)
    );

    bfr new_Jinkela_buffer_2195 (
        .din(new_Jinkela_wire_2575),
        .dout(new_Jinkela_wire_2576)
    );

    bfr new_Jinkela_buffer_2150 (
        .din(new_Jinkela_wire_2524),
        .dout(new_Jinkela_wire_2525)
    );

    and_ii n_2399_ (
        .a(n_0273_),
        .b(n_0272_),
        .c(n_0274_)
    );

    and_bb n_2400_ (
        .a(new_Jinkela_wire_9382),
        .b(new_Jinkela_wire_8317),
        .c(n_0275_)
    );

    bfr new_Jinkela_buffer_2151 (
        .din(new_Jinkela_wire_2525),
        .dout(new_Jinkela_wire_2526)
    );

    and_bb n_2401_ (
        .a(new_Jinkela_wire_4972),
        .b(new_Jinkela_wire_10223),
        .c(n_0276_)
    );

    bfr new_Jinkela_buffer_2211 (
        .din(new_Jinkela_wire_2597),
        .dout(new_Jinkela_wire_2598)
    );

    and_ii n_2402_ (
        .a(new_Jinkela_wire_5225),
        .b(new_Jinkela_wire_5232),
        .c(n_0277_)
    );

    bfr new_Jinkela_buffer_2196 (
        .din(new_Jinkela_wire_2576),
        .dout(new_Jinkela_wire_2577)
    );

    bfr new_Jinkela_buffer_2152 (
        .din(new_Jinkela_wire_2526),
        .dout(new_Jinkela_wire_2527)
    );

    or_ii n_2403_ (
        .a(n_0277_),
        .b(new_Jinkela_wire_5638),
        .c(n_0278_)
    );

    and_bi n_2404_ (
        .a(new_Jinkela_wire_3843),
        .b(new_Jinkela_wire_9598),
        .c(n_0279_)
    );

    bfr new_Jinkela_buffer_2153 (
        .din(new_Jinkela_wire_2527),
        .dout(new_Jinkela_wire_2528)
    );

    and_ii n_2405_ (
        .a(new_Jinkela_wire_3713),
        .b(new_Jinkela_wire_7120),
        .c(n_0280_)
    );

    bfr new_Jinkela_buffer_2275 (
        .din(new_Jinkela_wire_2661),
        .dout(new_Jinkela_wire_2662)
    );

    and_bb n_2406_ (
        .a(new_Jinkela_wire_3715),
        .b(new_Jinkela_wire_7119),
        .c(n_0281_)
    );

    bfr new_Jinkela_buffer_2197 (
        .din(new_Jinkela_wire_2577),
        .dout(new_Jinkela_wire_2578)
    );

    bfr new_Jinkela_buffer_2154 (
        .din(new_Jinkela_wire_2528),
        .dout(new_Jinkela_wire_2529)
    );

    and_ii n_2407_ (
        .a(new_Jinkela_wire_7837),
        .b(new_Jinkela_wire_6815),
        .c(n_0282_)
    );

    or_ii n_2408_ (
        .a(new_Jinkela_wire_7848),
        .b(new_Jinkela_wire_6709),
        .c(n_0283_)
    );

    bfr new_Jinkela_buffer_4741 (
        .din(new_Jinkela_wire_5660),
        .dout(new_Jinkela_wire_5661)
    );

    and_bi n_1653_ (
        .a(new_Jinkela_wire_9150),
        .b(new_Jinkela_wire_10556),
        .c(n_0920_)
    );

    bfr new_Jinkela_buffer_7356 (
        .din(n_0614_),
        .dout(new_Jinkela_wire_9135)
    );

    bfr new_Jinkela_buffer_7284 (
        .din(new_Jinkela_wire_9047),
        .dout(new_Jinkela_wire_9048)
    );

    bfr new_Jinkela_buffer_4722 (
        .din(new_Jinkela_wire_5627),
        .dout(new_Jinkela_wire_5628)
    );

    and_ii n_1654_ (
        .a(n_0920_),
        .b(n_0919_),
        .c(n_0921_)
    );

    spl2 new_Jinkela_splitter_712 (
        .a(n_1370_),
        .b(new_Jinkela_wire_9118),
        .c(new_Jinkela_wire_9119)
    );

    bfr new_Jinkela_buffer_4759 (
        .din(new_Jinkela_wire_5686),
        .dout(new_Jinkela_wire_5687)
    );

    and_ii n_1655_ (
        .a(new_Jinkela_wire_4998),
        .b(new_Jinkela_wire_3772),
        .c(n_0922_)
    );

    bfr new_Jinkela_buffer_7326 (
        .din(new_Jinkela_wire_9095),
        .dout(new_Jinkela_wire_9096)
    );

    bfr new_Jinkela_buffer_7285 (
        .din(new_Jinkela_wire_9048),
        .dout(new_Jinkela_wire_9049)
    );

    bfr new_Jinkela_buffer_4723 (
        .din(new_Jinkela_wire_5628),
        .dout(new_Jinkela_wire_5629)
    );

    and_bb n_1656_ (
        .a(new_Jinkela_wire_4997),
        .b(new_Jinkela_wire_3771),
        .c(n_0923_)
    );

    bfr new_Jinkela_buffer_4742 (
        .din(new_Jinkela_wire_5661),
        .dout(new_Jinkela_wire_5662)
    );

    or_bb n_1657_ (
        .a(n_0923_),
        .b(n_0922_),
        .c(n_0924_)
    );

    bfr new_Jinkela_buffer_7341 (
        .din(new_Jinkela_wire_9113),
        .dout(new_Jinkela_wire_9114)
    );

    bfr new_Jinkela_buffer_7286 (
        .din(new_Jinkela_wire_9049),
        .dout(new_Jinkela_wire_9050)
    );

    bfr new_Jinkela_buffer_4724 (
        .din(new_Jinkela_wire_5629),
        .dout(new_Jinkela_wire_5630)
    );

    and_bi n_1658_ (
        .a(new_Jinkela_wire_1810),
        .b(new_Jinkela_wire_1283),
        .c(n_0925_)
    );

    and_bi n_1659_ (
        .a(new_Jinkela_wire_1194),
        .b(new_Jinkela_wire_1709),
        .c(n_0926_)
    );

    spl2 new_Jinkela_splitter_358 (
        .a(n_0833_),
        .b(new_Jinkela_wire_5874),
        .c(new_Jinkela_wire_5875)
    );

    bfr new_Jinkela_buffer_7327 (
        .din(new_Jinkela_wire_9096),
        .dout(new_Jinkela_wire_9097)
    );

    bfr new_Jinkela_buffer_7287 (
        .din(new_Jinkela_wire_9050),
        .dout(new_Jinkela_wire_9051)
    );

    bfr new_Jinkela_buffer_4725 (
        .din(new_Jinkela_wire_5630),
        .dout(new_Jinkela_wire_5631)
    );

    and_ii n_1660_ (
        .a(n_0926_),
        .b(n_0925_),
        .c(n_0927_)
    );

    bfr new_Jinkela_buffer_4743 (
        .din(new_Jinkela_wire_5662),
        .dout(new_Jinkela_wire_5663)
    );

    and_bi n_1661_ (
        .a(new_Jinkela_wire_430),
        .b(new_Jinkela_wire_1231),
        .c(n_0928_)
    );

    bfr new_Jinkela_buffer_7288 (
        .din(new_Jinkela_wire_9051),
        .dout(new_Jinkela_wire_9052)
    );

    bfr new_Jinkela_buffer_4726 (
        .din(new_Jinkela_wire_5631),
        .dout(new_Jinkela_wire_5632)
    );

    and_bi n_1662_ (
        .a(new_Jinkela_wire_1311),
        .b(new_Jinkela_wire_1834),
        .c(n_0929_)
    );

    spl2 new_Jinkela_splitter_714 (
        .a(n_0177_),
        .b(new_Jinkela_wire_9136),
        .c(new_Jinkela_wire_9137)
    );

    bfr new_Jinkela_buffer_4760 (
        .din(new_Jinkela_wire_5687),
        .dout(new_Jinkela_wire_5688)
    );

    and_ii n_1663_ (
        .a(n_0929_),
        .b(n_0928_),
        .c(n_0930_)
    );

    bfr new_Jinkela_buffer_7328 (
        .din(new_Jinkela_wire_9097),
        .dout(new_Jinkela_wire_9098)
    );

    bfr new_Jinkela_buffer_7289 (
        .din(new_Jinkela_wire_9052),
        .dout(new_Jinkela_wire_9053)
    );

    spl2 new_Jinkela_splitter_344 (
        .a(new_Jinkela_wire_5632),
        .b(new_Jinkela_wire_5633),
        .c(new_Jinkela_wire_5634)
    );

    and_ii n_1664_ (
        .a(new_Jinkela_wire_7201),
        .b(new_Jinkela_wire_9751),
        .c(n_0931_)
    );

    and_bb n_1665_ (
        .a(new_Jinkela_wire_7200),
        .b(new_Jinkela_wire_9750),
        .c(n_0932_)
    );

    bfr new_Jinkela_buffer_4804 (
        .din(new_Jinkela_wire_5735),
        .dout(new_Jinkela_wire_5736)
    );

    bfr new_Jinkela_buffer_7290 (
        .din(new_Jinkela_wire_9053),
        .dout(new_Jinkela_wire_9054)
    );

    bfr new_Jinkela_buffer_4744 (
        .din(new_Jinkela_wire_5663),
        .dout(new_Jinkela_wire_5664)
    );

    and_ii n_1666_ (
        .a(n_0932_),
        .b(n_0931_),
        .c(n_0933_)
    );

    bfr new_Jinkela_buffer_7342 (
        .din(new_Jinkela_wire_9114),
        .dout(new_Jinkela_wire_9115)
    );

    bfr new_Jinkela_buffer_4745 (
        .din(new_Jinkela_wire_5664),
        .dout(new_Jinkela_wire_5665)
    );

    or_bi n_1667_ (
        .a(new_Jinkela_wire_2978),
        .b(new_Jinkela_wire_1905),
        .c(n_0934_)
    );

    bfr new_Jinkela_buffer_7329 (
        .din(new_Jinkela_wire_9098),
        .dout(new_Jinkela_wire_9099)
    );

    bfr new_Jinkela_buffer_7291 (
        .din(new_Jinkela_wire_9054),
        .dout(new_Jinkela_wire_9055)
    );

    bfr new_Jinkela_buffer_4761 (
        .din(new_Jinkela_wire_5688),
        .dout(new_Jinkela_wire_5689)
    );

    and_bi n_1668_ (
        .a(new_Jinkela_wire_2977),
        .b(new_Jinkela_wire_1906),
        .c(n_0935_)
    );

    bfr new_Jinkela_buffer_4746 (
        .din(new_Jinkela_wire_5665),
        .dout(new_Jinkela_wire_5666)
    );

    and_bi n_1669_ (
        .a(n_0934_),
        .b(n_0935_),
        .c(n_0936_)
    );

    bfr new_Jinkela_buffer_7292 (
        .din(new_Jinkela_wire_9055),
        .dout(new_Jinkela_wire_9056)
    );

    and_bi n_1670_ (
        .a(new_Jinkela_wire_1393),
        .b(new_Jinkela_wire_7243),
        .c(n_0937_)
    );

    bfr new_Jinkela_buffer_4869 (
        .din(new_Jinkela_wire_5805),
        .dout(new_Jinkela_wire_5806)
    );

    bfr new_Jinkela_buffer_7343 (
        .din(new_Jinkela_wire_9119),
        .dout(new_Jinkela_wire_9120)
    );

    bfr new_Jinkela_buffer_4747 (
        .din(new_Jinkela_wire_5666),
        .dout(new_Jinkela_wire_5667)
    );

    or_bb n_1671_ (
        .a(new_Jinkela_wire_600),
        .b(new_Jinkela_wire_1166),
        .c(n_0938_)
    );

    bfr new_Jinkela_buffer_7330 (
        .din(new_Jinkela_wire_9099),
        .dout(new_Jinkela_wire_9100)
    );

    bfr new_Jinkela_buffer_7293 (
        .din(new_Jinkela_wire_9056),
        .dout(new_Jinkela_wire_9057)
    );

    bfr new_Jinkela_buffer_4762 (
        .din(new_Jinkela_wire_5689),
        .dout(new_Jinkela_wire_5690)
    );

    and_bb n_1672_ (
        .a(new_Jinkela_wire_599),
        .b(new_Jinkela_wire_1165),
        .c(n_0939_)
    );

    bfr new_Jinkela_buffer_4748 (
        .din(new_Jinkela_wire_5667),
        .dout(new_Jinkela_wire_5668)
    );

    or_bb n_1673_ (
        .a(new_Jinkela_wire_7828),
        .b(new_Jinkela_wire_1394),
        .c(n_0940_)
    );

    spl3L new_Jinkela_splitter_715 (
        .a(n_0482_),
        .d(new_Jinkela_wire_9138),
        .b(new_Jinkela_wire_9139),
        .c(new_Jinkela_wire_9140)
    );

    bfr new_Jinkela_buffer_7294 (
        .din(new_Jinkela_wire_9057),
        .dout(new_Jinkela_wire_9058)
    );

    bfr new_Jinkela_buffer_4824 (
        .din(new_Jinkela_wire_5758),
        .dout(new_Jinkela_wire_5759)
    );

    and_bi n_1674_ (
        .a(new_Jinkela_wire_5155),
        .b(n_0940_),
        .c(n_0941_)
    );

    bfr new_Jinkela_buffer_4805 (
        .din(new_Jinkela_wire_5736),
        .dout(new_Jinkela_wire_5737)
    );

    spl2 new_Jinkela_splitter_711 (
        .a(new_Jinkela_wire_9115),
        .b(new_Jinkela_wire_9116),
        .c(new_Jinkela_wire_9117)
    );

    bfr new_Jinkela_buffer_4749 (
        .din(new_Jinkela_wire_5668),
        .dout(new_Jinkela_wire_5669)
    );

    and_ii n_1675_ (
        .a(n_0941_),
        .b(new_Jinkela_wire_4665),
        .c(n_0942_)
    );

    bfr new_Jinkela_buffer_7331 (
        .din(new_Jinkela_wire_9100),
        .dout(new_Jinkela_wire_9101)
    );

    bfr new_Jinkela_buffer_7295 (
        .din(new_Jinkela_wire_9058),
        .dout(new_Jinkela_wire_9059)
    );

    bfr new_Jinkela_buffer_4763 (
        .din(new_Jinkela_wire_5690),
        .dout(new_Jinkela_wire_5691)
    );

    and_ii n_1676_ (
        .a(new_Jinkela_wire_3770),
        .b(new_Jinkela_wire_5072),
        .c(n_0943_)
    );

    bfr new_Jinkela_buffer_4750 (
        .din(new_Jinkela_wire_5669),
        .dout(new_Jinkela_wire_5670)
    );

    and_bb n_1677_ (
        .a(new_Jinkela_wire_3769),
        .b(new_Jinkela_wire_5071),
        .c(n_0944_)
    );

    bfr new_Jinkela_buffer_7296 (
        .din(new_Jinkela_wire_9059),
        .dout(new_Jinkela_wire_9060)
    );

    and_ii n_1678_ (
        .a(n_0944_),
        .b(n_0943_),
        .c(n_0945_)
    );

    bfr new_Jinkela_buffer_4751 (
        .din(new_Jinkela_wire_5670),
        .dout(new_Jinkela_wire_5671)
    );

    or_bb n_1679_ (
        .a(new_Jinkela_wire_4969),
        .b(new_Jinkela_wire_6189),
        .c(n_0946_)
    );

    bfr new_Jinkela_buffer_7332 (
        .din(new_Jinkela_wire_9101),
        .dout(new_Jinkela_wire_9102)
    );

    bfr new_Jinkela_buffer_7297 (
        .din(new_Jinkela_wire_9060),
        .dout(new_Jinkela_wire_9061)
    );

    bfr new_Jinkela_buffer_4764 (
        .din(new_Jinkela_wire_5691),
        .dout(new_Jinkela_wire_5692)
    );

    and_bb n_1680_ (
        .a(new_Jinkela_wire_4968),
        .b(new_Jinkela_wire_6188),
        .c(n_0947_)
    );

    bfr new_Jinkela_buffer_4752 (
        .din(new_Jinkela_wire_5671),
        .dout(new_Jinkela_wire_5672)
    );

    and_bi n_1681_ (
        .a(n_0946_),
        .b(n_0947_),
        .c(n_0948_)
    );

    bfr new_Jinkela_buffer_7344 (
        .din(new_Jinkela_wire_9120),
        .dout(new_Jinkela_wire_9121)
    );

    bfr new_Jinkela_buffer_7298 (
        .din(new_Jinkela_wire_9061),
        .dout(new_Jinkela_wire_9062)
    );

    and_bb n_1682_ (
        .a(new_Jinkela_wire_1388),
        .b(new_Jinkela_wire_2240),
        .c(n_0949_)
    );

    bfr new_Jinkela_buffer_4806 (
        .din(new_Jinkela_wire_5737),
        .dout(new_Jinkela_wire_5738)
    );

    bfr new_Jinkela_buffer_4753 (
        .din(new_Jinkela_wire_5672),
        .dout(new_Jinkela_wire_5673)
    );

    and_ii n_1683_ (
        .a(new_Jinkela_wire_2590),
        .b(new_Jinkela_wire_1207),
        .c(n_0950_)
    );

    bfr new_Jinkela_buffer_7333 (
        .din(new_Jinkela_wire_9102),
        .dout(new_Jinkela_wire_9103)
    );

    bfr new_Jinkela_buffer_7299 (
        .din(new_Jinkela_wire_9062),
        .dout(new_Jinkela_wire_9063)
    );

    bfr new_Jinkela_buffer_4765 (
        .din(new_Jinkela_wire_5692),
        .dout(new_Jinkela_wire_5693)
    );

    and_ii n_1684_ (
        .a(new_Jinkela_wire_9297),
        .b(new_Jinkela_wire_9886),
        .c(n_0951_)
    );

    bfr new_Jinkela_buffer_4754 (
        .din(new_Jinkela_wire_5673),
        .dout(new_Jinkela_wire_5674)
    );

    and_bi n_1685_ (
        .a(new_Jinkela_wire_511),
        .b(new_Jinkela_wire_1277),
        .c(n_0952_)
    );

    bfr new_Jinkela_buffer_7300 (
        .din(new_Jinkela_wire_9063),
        .dout(new_Jinkela_wire_9064)
    );

    and_bi n_1686_ (
        .a(new_Jinkela_wire_1378),
        .b(new_Jinkela_wire_1101),
        .c(n_0953_)
    );

    spl3L new_Jinkela_splitter_359 (
        .a(n_0115_),
        .d(new_Jinkela_wire_5876),
        .b(new_Jinkela_wire_5877),
        .c(new_Jinkela_wire_5878)
    );

    bfr new_Jinkela_buffer_4755 (
        .din(new_Jinkela_wire_5674),
        .dout(new_Jinkela_wire_5675)
    );

    and_ii n_1687_ (
        .a(n_0953_),
        .b(n_0952_),
        .c(n_0954_)
    );

    bfr new_Jinkela_buffer_7334 (
        .din(new_Jinkela_wire_9103),
        .dout(new_Jinkela_wire_9104)
    );

    bfr new_Jinkela_buffer_7301 (
        .din(new_Jinkela_wire_9064),
        .dout(new_Jinkela_wire_9065)
    );

    bfr new_Jinkela_buffer_4766 (
        .din(new_Jinkela_wire_5693),
        .dout(new_Jinkela_wire_5694)
    );

    and_bi n_1688_ (
        .a(new_Jinkela_wire_3935),
        .b(new_Jinkela_wire_8078),
        .c(n_0955_)
    );

    bfr new_Jinkela_buffer_4825 (
        .din(new_Jinkela_wire_5759),
        .dout(new_Jinkela_wire_5760)
    );

    and_bi n_1689_ (
        .a(new_Jinkela_wire_8077),
        .b(new_Jinkela_wire_3934),
        .c(n_0956_)
    );

    bfr new_Jinkela_buffer_4807 (
        .din(new_Jinkela_wire_5738),
        .dout(new_Jinkela_wire_5739)
    );

    bfr new_Jinkela_buffer_7302 (
        .din(new_Jinkela_wire_9065),
        .dout(new_Jinkela_wire_9066)
    );

    bfr new_Jinkela_buffer_4767 (
        .din(new_Jinkela_wire_5694),
        .dout(new_Jinkela_wire_5695)
    );

    and_ii n_1690_ (
        .a(n_0956_),
        .b(n_0955_),
        .c(n_0957_)
    );

    spl2 new_Jinkela_splitter_716 (
        .a(n_0105_),
        .b(new_Jinkela_wire_9141),
        .c(new_Jinkela_wire_9142)
    );

    and_bi n_1691_ (
        .a(new_Jinkela_wire_1989),
        .b(new_Jinkela_wire_1271),
        .c(n_0958_)
    );

    bfr new_Jinkela_buffer_7335 (
        .din(new_Jinkela_wire_9104),
        .dout(new_Jinkela_wire_9105)
    );

    bfr new_Jinkela_buffer_7303 (
        .din(new_Jinkela_wire_9066),
        .dout(new_Jinkela_wire_9067)
    );

    bfr new_Jinkela_buffer_4768 (
        .din(new_Jinkela_wire_5695),
        .dout(new_Jinkela_wire_5696)
    );

    and_bi n_1692_ (
        .a(new_Jinkela_wire_1266),
        .b(new_Jinkela_wire_883),
        .c(n_0959_)
    );

    bfr new_Jinkela_buffer_4933 (
        .din(new_Jinkela_wire_5872),
        .dout(new_Jinkela_wire_5873)
    );

    and_ii n_1693_ (
        .a(n_0959_),
        .b(n_0958_),
        .c(n_0960_)
    );

    bfr new_Jinkela_buffer_4808 (
        .din(new_Jinkela_wire_5739),
        .dout(new_Jinkela_wire_5740)
    );

    bfr new_Jinkela_buffer_7345 (
        .din(new_Jinkela_wire_9121),
        .dout(new_Jinkela_wire_9122)
    );

    bfr new_Jinkela_buffer_7304 (
        .din(new_Jinkela_wire_9067),
        .dout(new_Jinkela_wire_9068)
    );

    bfr new_Jinkela_buffer_4769 (
        .din(new_Jinkela_wire_5696),
        .dout(new_Jinkela_wire_5697)
    );

    and_bi n_1694_ (
        .a(new_Jinkela_wire_1977),
        .b(new_Jinkela_wire_1347),
        .c(n_0961_)
    );

    bfr new_Jinkela_buffer_864 (
        .din(new_Jinkela_wire_929),
        .dout(new_Jinkela_wire_930)
    );

    bfr new_Jinkela_buffer_1021 (
        .din(new_Jinkela_wire_1095),
        .dout(new_Jinkela_wire_1096)
    );

    bfr new_Jinkela_buffer_865 (
        .din(new_Jinkela_wire_930),
        .dout(new_Jinkela_wire_931)
    );

    bfr new_Jinkela_buffer_905 (
        .din(new_Jinkela_wire_975),
        .dout(new_Jinkela_wire_976)
    );

    bfr new_Jinkela_buffer_866 (
        .din(new_Jinkela_wire_931),
        .dout(new_Jinkela_wire_932)
    );

    bfr new_Jinkela_buffer_957 (
        .din(new_Jinkela_wire_1031),
        .dout(new_Jinkela_wire_1032)
    );

    bfr new_Jinkela_buffer_867 (
        .din(new_Jinkela_wire_932),
        .dout(new_Jinkela_wire_933)
    );

    bfr new_Jinkela_buffer_906 (
        .din(new_Jinkela_wire_976),
        .dout(new_Jinkela_wire_977)
    );

    bfr new_Jinkela_buffer_868 (
        .din(new_Jinkela_wire_933),
        .dout(new_Jinkela_wire_934)
    );

    spl3L new_Jinkela_splitter_35 (
        .a(N18),
        .d(new_Jinkela_wire_1167),
        .b(new_Jinkela_wire_1221),
        .c(new_Jinkela_wire_1306)
    );

    bfr new_Jinkela_buffer_1024 (
        .din(new_Jinkela_wire_1098),
        .dout(new_Jinkela_wire_1099)
    );

    bfr new_Jinkela_buffer_869 (
        .din(new_Jinkela_wire_934),
        .dout(new_Jinkela_wire_935)
    );

    bfr new_Jinkela_buffer_907 (
        .din(new_Jinkela_wire_977),
        .dout(new_Jinkela_wire_978)
    );

    bfr new_Jinkela_buffer_870 (
        .din(new_Jinkela_wire_935),
        .dout(new_Jinkela_wire_936)
    );

    bfr new_Jinkela_buffer_958 (
        .din(new_Jinkela_wire_1032),
        .dout(new_Jinkela_wire_1033)
    );

    bfr new_Jinkela_buffer_871 (
        .din(new_Jinkela_wire_936),
        .dout(new_Jinkela_wire_937)
    );

    bfr new_Jinkela_buffer_908 (
        .din(new_Jinkela_wire_978),
        .dout(new_Jinkela_wire_979)
    );

    bfr new_Jinkela_buffer_872 (
        .din(new_Jinkela_wire_937),
        .dout(new_Jinkela_wire_938)
    );

    bfr new_Jinkela_buffer_1022 (
        .din(new_Jinkela_wire_1096),
        .dout(new_Jinkela_wire_1097)
    );

    bfr new_Jinkela_buffer_873 (
        .din(new_Jinkela_wire_938),
        .dout(new_Jinkela_wire_939)
    );

    bfr new_Jinkela_buffer_909 (
        .din(new_Jinkela_wire_979),
        .dout(new_Jinkela_wire_980)
    );

    bfr new_Jinkela_buffer_874 (
        .din(new_Jinkela_wire_939),
        .dout(new_Jinkela_wire_940)
    );

    bfr new_Jinkela_buffer_959 (
        .din(new_Jinkela_wire_1033),
        .dout(new_Jinkela_wire_1034)
    );

    bfr new_Jinkela_buffer_875 (
        .din(new_Jinkela_wire_940),
        .dout(new_Jinkela_wire_941)
    );

    bfr new_Jinkela_buffer_910 (
        .din(new_Jinkela_wire_980),
        .dout(new_Jinkela_wire_981)
    );

    bfr new_Jinkela_buffer_876 (
        .din(new_Jinkela_wire_941),
        .dout(new_Jinkela_wire_942)
    );

    bfr new_Jinkela_buffer_877 (
        .din(new_Jinkela_wire_942),
        .dout(new_Jinkela_wire_943)
    );

    bfr new_Jinkela_buffer_911 (
        .din(new_Jinkela_wire_981),
        .dout(new_Jinkela_wire_982)
    );

    bfr new_Jinkela_buffer_878 (
        .din(new_Jinkela_wire_943),
        .dout(new_Jinkela_wire_944)
    );

    bfr new_Jinkela_buffer_960 (
        .din(new_Jinkela_wire_1034),
        .dout(new_Jinkela_wire_1035)
    );

    bfr new_Jinkela_buffer_879 (
        .din(new_Jinkela_wire_944),
        .dout(new_Jinkela_wire_945)
    );

    bfr new_Jinkela_buffer_912 (
        .din(new_Jinkela_wire_982),
        .dout(new_Jinkela_wire_983)
    );

    bfr new_Jinkela_buffer_880 (
        .din(new_Jinkela_wire_945),
        .dout(new_Jinkela_wire_946)
    );

    bfr new_Jinkela_buffer_1025 (
        .din(new_Jinkela_wire_1099),
        .dout(new_Jinkela_wire_1100)
    );

    bfr new_Jinkela_buffer_881 (
        .din(new_Jinkela_wire_946),
        .dout(new_Jinkela_wire_947)
    );

    bfr new_Jinkela_buffer_913 (
        .din(new_Jinkela_wire_983),
        .dout(new_Jinkela_wire_984)
    );

    bfr new_Jinkela_buffer_882 (
        .din(new_Jinkela_wire_947),
        .dout(new_Jinkela_wire_948)
    );

    bfr new_Jinkela_buffer_961 (
        .din(new_Jinkela_wire_1035),
        .dout(new_Jinkela_wire_1036)
    );

    bfr new_Jinkela_buffer_914 (
        .din(new_Jinkela_wire_984),
        .dout(new_Jinkela_wire_985)
    );

    bfr new_Jinkela_buffer_1088 (
        .din(N179),
        .dout(new_Jinkela_wire_1395)
    );

    bfr new_Jinkela_buffer_915 (
        .din(new_Jinkela_wire_985),
        .dout(new_Jinkela_wire_986)
    );

    bfr new_Jinkela_buffer_962 (
        .din(new_Jinkela_wire_1036),
        .dout(new_Jinkela_wire_1037)
    );

    bfr new_Jinkela_buffer_6423 (
        .din(new_Jinkela_wire_7847),
        .dout(new_Jinkela_wire_7848)
    );

    bfr new_Jinkela_buffer_3123 (
        .din(new_Jinkela_wire_3559),
        .dout(new_Jinkela_wire_3560)
    );

    bfr new_Jinkela_buffer_2155 (
        .din(new_Jinkela_wire_2529),
        .dout(new_Jinkela_wire_2530)
    );

    bfr new_Jinkela_buffer_3059 (
        .din(new_Jinkela_wire_3488),
        .dout(new_Jinkela_wire_3489)
    );

    bfr new_Jinkela_buffer_7336 (
        .din(new_Jinkela_wire_9105),
        .dout(new_Jinkela_wire_9106)
    );

    bfr new_Jinkela_buffer_7305 (
        .din(new_Jinkela_wire_9068),
        .dout(new_Jinkela_wire_9069)
    );

    bfr new_Jinkela_buffer_2212 (
        .din(new_Jinkela_wire_2598),
        .dout(new_Jinkela_wire_2599)
    );

    bfr new_Jinkela_buffer_2198 (
        .din(new_Jinkela_wire_2578),
        .dout(new_Jinkela_wire_2579)
    );

    bfr new_Jinkela_buffer_3121 (
        .din(new_Jinkela_wire_3557),
        .dout(new_Jinkela_wire_3558)
    );

    bfr new_Jinkela_buffer_2156 (
        .din(new_Jinkela_wire_2530),
        .dout(new_Jinkela_wire_2531)
    );

    bfr new_Jinkela_buffer_3060 (
        .din(new_Jinkela_wire_3489),
        .dout(new_Jinkela_wire_3490)
    );

    bfr new_Jinkela_buffer_6426 (
        .din(new_Jinkela_wire_7852),
        .dout(new_Jinkela_wire_7853)
    );

    bfr new_Jinkela_buffer_7306 (
        .din(new_Jinkela_wire_9069),
        .dout(new_Jinkela_wire_9070)
    );

    spl2 new_Jinkela_splitter_566 (
        .a(n_0406_),
        .b(new_Jinkela_wire_7921),
        .c(new_Jinkela_wire_7922)
    );

    bfr new_Jinkela_buffer_2157 (
        .din(new_Jinkela_wire_2531),
        .dout(new_Jinkela_wire_2532)
    );

    bfr new_Jinkela_buffer_3061 (
        .din(new_Jinkela_wire_3490),
        .dout(new_Jinkela_wire_3491)
    );

    bfr new_Jinkela_buffer_6427 (
        .din(new_Jinkela_wire_7853),
        .dout(new_Jinkela_wire_7854)
    );

    bfr new_Jinkela_buffer_7357 (
        .din(new_net_9),
        .dout(new_Jinkela_wire_9143)
    );

    spl2 new_Jinkela_splitter_567 (
        .a(n_0268_),
        .b(new_Jinkela_wire_7923),
        .c(new_Jinkela_wire_7924)
    );

    bfr new_Jinkela_buffer_2199 (
        .din(new_Jinkela_wire_2579),
        .dout(new_Jinkela_wire_2580)
    );

    bfr new_Jinkela_buffer_3126 (
        .din(new_Jinkela_wire_3564),
        .dout(new_Jinkela_wire_3565)
    );

    bfr new_Jinkela_buffer_6488 (
        .din(new_Jinkela_wire_7916),
        .dout(new_Jinkela_wire_7917)
    );

    bfr new_Jinkela_buffer_7337 (
        .din(new_Jinkela_wire_9106),
        .dout(new_Jinkela_wire_9107)
    );

    bfr new_Jinkela_buffer_3124 (
        .din(new_Jinkela_wire_3560),
        .dout(new_Jinkela_wire_3561)
    );

    bfr new_Jinkela_buffer_2158 (
        .din(new_Jinkela_wire_2532),
        .dout(new_Jinkela_wire_2533)
    );

    bfr new_Jinkela_buffer_3062 (
        .din(new_Jinkela_wire_3491),
        .dout(new_Jinkela_wire_3492)
    );

    bfr new_Jinkela_buffer_6428 (
        .din(new_Jinkela_wire_7854),
        .dout(new_Jinkela_wire_7855)
    );

    bfr new_Jinkela_buffer_7346 (
        .din(new_Jinkela_wire_9122),
        .dout(new_Jinkela_wire_9123)
    );

    bfr new_Jinkela_buffer_7308 (
        .din(new_Jinkela_wire_9071),
        .dout(new_Jinkela_wire_9072)
    );

    bfr new_Jinkela_buffer_2344 (
        .din(N313),
        .dout(new_Jinkela_wire_2736)
    );

    spl2 new_Jinkela_splitter_568 (
        .a(n_0889_),
        .b(new_Jinkela_wire_7927),
        .c(new_Jinkela_wire_7928)
    );

    bfr new_Jinkela_buffer_2159 (
        .din(new_Jinkela_wire_2533),
        .dout(new_Jinkela_wire_2534)
    );

    bfr new_Jinkela_buffer_3063 (
        .din(new_Jinkela_wire_3492),
        .dout(new_Jinkela_wire_3493)
    );

    bfr new_Jinkela_buffer_6429 (
        .din(new_Jinkela_wire_7855),
        .dout(new_Jinkela_wire_7856)
    );

    bfr new_Jinkela_buffer_7338 (
        .din(new_Jinkela_wire_9107),
        .dout(new_Jinkela_wire_9108)
    );

    bfr new_Jinkela_buffer_7309 (
        .din(new_Jinkela_wire_9072),
        .dout(new_Jinkela_wire_9073)
    );

    bfr new_Jinkela_buffer_2213 (
        .din(new_Jinkela_wire_2599),
        .dout(new_Jinkela_wire_2600)
    );

    bfr new_Jinkela_buffer_2200 (
        .din(new_Jinkela_wire_2580),
        .dout(new_Jinkela_wire_2581)
    );

    bfr new_Jinkela_buffer_6489 (
        .din(new_Jinkela_wire_7917),
        .dout(new_Jinkela_wire_7918)
    );

    bfr new_Jinkela_buffer_3125 (
        .din(new_Jinkela_wire_3561),
        .dout(new_Jinkela_wire_3562)
    );

    bfr new_Jinkela_buffer_2160 (
        .din(new_Jinkela_wire_2534),
        .dout(new_Jinkela_wire_2535)
    );

    bfr new_Jinkela_buffer_3064 (
        .din(new_Jinkela_wire_3493),
        .dout(new_Jinkela_wire_3494)
    );

    bfr new_Jinkela_buffer_6430 (
        .din(new_Jinkela_wire_7856),
        .dout(new_Jinkela_wire_7857)
    );

    bfr new_Jinkela_buffer_7310 (
        .din(new_Jinkela_wire_9073),
        .dout(new_Jinkela_wire_9074)
    );

    bfr new_Jinkela_buffer_3139 (
        .din(n_0885_),
        .dout(new_Jinkela_wire_3578)
    );

    bfr new_Jinkela_buffer_2161 (
        .din(new_Jinkela_wire_2535),
        .dout(new_Jinkela_wire_2536)
    );

    bfr new_Jinkela_buffer_3065 (
        .din(new_Jinkela_wire_3494),
        .dout(new_Jinkela_wire_3495)
    );

    bfr new_Jinkela_buffer_6431 (
        .din(new_Jinkela_wire_7857),
        .dout(new_Jinkela_wire_7858)
    );

    bfr new_Jinkela_buffer_7360 (
        .din(n_0195_),
        .dout(new_Jinkela_wire_9148)
    );

    bfr new_Jinkela_buffer_6490 (
        .din(new_Jinkela_wire_7924),
        .dout(new_Jinkela_wire_7925)
    );

    bfr new_Jinkela_buffer_2278 (
        .din(new_Jinkela_wire_2664),
        .dout(new_Jinkela_wire_2665)
    );

    bfr new_Jinkela_buffer_2341 (
        .din(new_Jinkela_wire_2732),
        .dout(new_Jinkela_wire_2733)
    );

    spl2 new_Jinkela_splitter_565 (
        .a(new_Jinkela_wire_7918),
        .b(new_Jinkela_wire_7919),
        .c(new_Jinkela_wire_7920)
    );

    bfr new_Jinkela_buffer_7339 (
        .din(new_Jinkela_wire_9108),
        .dout(new_Jinkela_wire_9109)
    );

    bfr new_Jinkela_buffer_7311 (
        .din(new_Jinkela_wire_9074),
        .dout(new_Jinkela_wire_9075)
    );

    spl4L new_Jinkela_splitter_150 (
        .a(n_1153_),
        .d(new_Jinkela_wire_3579),
        .b(new_Jinkela_wire_3580),
        .e(new_Jinkela_wire_3581),
        .c(new_Jinkela_wire_3582)
    );

    bfr new_Jinkela_buffer_2162 (
        .din(new_Jinkela_wire_2536),
        .dout(new_Jinkela_wire_2537)
    );

    bfr new_Jinkela_buffer_3066 (
        .din(new_Jinkela_wire_3495),
        .dout(new_Jinkela_wire_3496)
    );

    bfr new_Jinkela_buffer_6432 (
        .din(new_Jinkela_wire_7858),
        .dout(new_Jinkela_wire_7859)
    );

    bfr new_Jinkela_buffer_7347 (
        .din(new_Jinkela_wire_9123),
        .dout(new_Jinkela_wire_9124)
    );

    bfr new_Jinkela_buffer_7312 (
        .din(new_Jinkela_wire_9075),
        .dout(new_Jinkela_wire_9076)
    );

    bfr new_Jinkela_buffer_2214 (
        .din(new_Jinkela_wire_2600),
        .dout(new_Jinkela_wire_2601)
    );

    bfr new_Jinkela_buffer_3127 (
        .din(new_Jinkela_wire_3565),
        .dout(new_Jinkela_wire_3566)
    );

    bfr new_Jinkela_buffer_2163 (
        .din(new_Jinkela_wire_2537),
        .dout(new_Jinkela_wire_2538)
    );

    bfr new_Jinkela_buffer_3067 (
        .din(new_Jinkela_wire_3496),
        .dout(new_Jinkela_wire_3497)
    );

    bfr new_Jinkela_buffer_6433 (
        .din(new_Jinkela_wire_7859),
        .dout(new_Jinkela_wire_7860)
    );

    bfr new_Jinkela_buffer_7359 (
        .din(n_0455_),
        .dout(new_Jinkela_wire_9147)
    );

    bfr new_Jinkela_buffer_7313 (
        .din(new_Jinkela_wire_9076),
        .dout(new_Jinkela_wire_9077)
    );

    bfr new_Jinkela_buffer_6788 (
        .din(n_0876_),
        .dout(new_Jinkela_wire_8383)
    );

    bfr new_Jinkela_buffer_2277 (
        .din(new_Jinkela_wire_2663),
        .dout(new_Jinkela_wire_2664)
    );

    spl3L new_Jinkela_splitter_151 (
        .a(n_1066_),
        .d(new_Jinkela_wire_3583),
        .b(new_Jinkela_wire_3584),
        .c(new_Jinkela_wire_3585)
    );

    spl2 new_Jinkela_splitter_152 (
        .a(new_Jinkela_wire_3585),
        .b(new_Jinkela_wire_3586),
        .c(new_Jinkela_wire_3587)
    );

    bfr new_Jinkela_buffer_2164 (
        .din(new_Jinkela_wire_2538),
        .dout(new_Jinkela_wire_2539)
    );

    bfr new_Jinkela_buffer_3068 (
        .din(new_Jinkela_wire_3497),
        .dout(new_Jinkela_wire_3498)
    );

    bfr new_Jinkela_buffer_6434 (
        .din(new_Jinkela_wire_7860),
        .dout(new_Jinkela_wire_7861)
    );

    bfr new_Jinkela_buffer_2215 (
        .din(new_Jinkela_wire_2601),
        .dout(new_Jinkela_wire_2602)
    );

    bfr new_Jinkela_buffer_3128 (
        .din(new_Jinkela_wire_3566),
        .dout(new_Jinkela_wire_3567)
    );

    bfr new_Jinkela_buffer_6491 (
        .din(new_Jinkela_wire_7925),
        .dout(new_Jinkela_wire_7926)
    );

    bfr new_Jinkela_buffer_7348 (
        .din(new_Jinkela_wire_9124),
        .dout(new_Jinkela_wire_9125)
    );

    bfr new_Jinkela_buffer_2165 (
        .din(new_Jinkela_wire_2539),
        .dout(new_Jinkela_wire_2540)
    );

    bfr new_Jinkela_buffer_3069 (
        .din(new_Jinkela_wire_3498),
        .dout(new_Jinkela_wire_3499)
    );

    bfr new_Jinkela_buffer_6435 (
        .din(new_Jinkela_wire_7861),
        .dout(new_Jinkela_wire_7862)
    );

    bfr new_Jinkela_buffer_7315 (
        .din(new_Jinkela_wire_9078),
        .dout(new_Jinkela_wire_9079)
    );

    spl2 new_Jinkela_splitter_129 (
        .a(new_Jinkela_wire_2665),
        .b(new_Jinkela_wire_2666),
        .c(new_Jinkela_wire_2667)
    );

    bfr new_Jinkela_buffer_6494 (
        .din(n_1150_),
        .dout(new_Jinkela_wire_7934)
    );

    bfr new_Jinkela_buffer_2166 (
        .din(new_Jinkela_wire_2540),
        .dout(new_Jinkela_wire_2541)
    );

    bfr new_Jinkela_buffer_3070 (
        .din(new_Jinkela_wire_3499),
        .dout(new_Jinkela_wire_3500)
    );

    bfr new_Jinkela_buffer_6436 (
        .din(new_Jinkela_wire_7862),
        .dout(new_Jinkela_wire_7863)
    );

    bfr new_Jinkela_buffer_6492 (
        .din(n_0798_),
        .dout(new_Jinkela_wire_7932)
    );

    bfr new_Jinkela_buffer_2216 (
        .din(new_Jinkela_wire_2602),
        .dout(new_Jinkela_wire_2603)
    );

    bfr new_Jinkela_buffer_3129 (
        .din(new_Jinkela_wire_3567),
        .dout(new_Jinkela_wire_3568)
    );

    bfr new_Jinkela_buffer_6493 (
        .din(new_Jinkela_wire_7932),
        .dout(new_Jinkela_wire_7933)
    );

    bfr new_Jinkela_buffer_7349 (
        .din(new_Jinkela_wire_9125),
        .dout(new_Jinkela_wire_9126)
    );

    bfr new_Jinkela_buffer_7316 (
        .din(new_Jinkela_wire_9079),
        .dout(new_Jinkela_wire_9080)
    );

    bfr new_Jinkela_buffer_2167 (
        .din(new_Jinkela_wire_2541),
        .dout(new_Jinkela_wire_2542)
    );

    bfr new_Jinkela_buffer_3071 (
        .din(new_Jinkela_wire_3500),
        .dout(new_Jinkela_wire_3501)
    );

    bfr new_Jinkela_buffer_6437 (
        .din(new_Jinkela_wire_7863),
        .dout(new_Jinkela_wire_7864)
    );

    bfr new_Jinkela_buffer_7361 (
        .din(n_0334_),
        .dout(new_Jinkela_wire_9149)
    );

    bfr new_Jinkela_buffer_7317 (
        .din(new_Jinkela_wire_9080),
        .dout(new_Jinkela_wire_9081)
    );

    spl2 new_Jinkela_splitter_570 (
        .a(n_0022_),
        .b(new_Jinkela_wire_7935),
        .c(new_Jinkela_wire_7936)
    );

    bfr new_Jinkela_buffer_2279 (
        .din(new_Jinkela_wire_2667),
        .dout(new_Jinkela_wire_2668)
    );

    bfr new_Jinkela_buffer_2168 (
        .din(new_Jinkela_wire_2542),
        .dout(new_Jinkela_wire_2543)
    );

    bfr new_Jinkela_buffer_3072 (
        .din(new_Jinkela_wire_3501),
        .dout(new_Jinkela_wire_3502)
    );

    bfr new_Jinkela_buffer_6438 (
        .din(new_Jinkela_wire_7864),
        .dout(new_Jinkela_wire_7865)
    );

    spl2 new_Jinkela_splitter_717 (
        .a(new_Jinkela_wire_9144),
        .b(new_Jinkela_wire_9145),
        .c(new_Jinkela_wire_9146)
    );

    bfr new_Jinkela_buffer_2217 (
        .din(new_Jinkela_wire_2603),
        .dout(new_Jinkela_wire_2604)
    );

    bfr new_Jinkela_buffer_3130 (
        .din(new_Jinkela_wire_3568),
        .dout(new_Jinkela_wire_3569)
    );

    bfr new_Jinkela_buffer_6495 (
        .din(new_net_2491),
        .dout(new_Jinkela_wire_7937)
    );

    bfr new_Jinkela_buffer_7318 (
        .din(new_Jinkela_wire_9081),
        .dout(new_Jinkela_wire_9082)
    );

    bfr new_Jinkela_buffer_2169 (
        .din(new_Jinkela_wire_2543),
        .dout(new_Jinkela_wire_2544)
    );

    bfr new_Jinkela_buffer_3073 (
        .din(new_Jinkela_wire_3502),
        .dout(new_Jinkela_wire_3503)
    );

    bfr new_Jinkela_buffer_6439 (
        .din(new_Jinkela_wire_7865),
        .dout(new_Jinkela_wire_7866)
    );

    bfr new_Jinkela_buffer_6537 (
        .din(n_1084_),
        .dout(new_Jinkela_wire_7985)
    );

    bfr new_Jinkela_buffer_2408 (
        .din(N83),
        .dout(new_Jinkela_wire_2805)
    );

    spl2 new_Jinkela_splitter_153 (
        .a(n_0301_),
        .b(new_Jinkela_wire_3588),
        .c(new_Jinkela_wire_3589)
    );

    bfr new_Jinkela_buffer_6496 (
        .din(new_Jinkela_wire_7937),
        .dout(new_Jinkela_wire_7938)
    );

    bfr new_Jinkela_buffer_7319 (
        .din(new_Jinkela_wire_9082),
        .dout(new_Jinkela_wire_9083)
    );

    bfr new_Jinkela_buffer_3141 (
        .din(new_Jinkela_wire_3590),
        .dout(new_Jinkela_wire_3591)
    );

    bfr new_Jinkela_buffer_2170 (
        .din(new_Jinkela_wire_2544),
        .dout(new_Jinkela_wire_2545)
    );

    bfr new_Jinkela_buffer_3074 (
        .din(new_Jinkela_wire_3503),
        .dout(new_Jinkela_wire_3504)
    );

    bfr new_Jinkela_buffer_6440 (
        .din(new_Jinkela_wire_7866),
        .dout(new_Jinkela_wire_7867)
    );

    spl2 new_Jinkela_splitter_720 (
        .a(n_0124_),
        .b(new_Jinkela_wire_9155),
        .c(new_Jinkela_wire_9156)
    );

    bfr new_Jinkela_buffer_7351 (
        .din(new_Jinkela_wire_9127),
        .dout(new_Jinkela_wire_9128)
    );

    bfr new_Jinkela_buffer_7320 (
        .din(new_Jinkela_wire_9083),
        .dout(new_Jinkela_wire_9084)
    );

    bfr new_Jinkela_buffer_2218 (
        .din(new_Jinkela_wire_2604),
        .dout(new_Jinkela_wire_2605)
    );

    bfr new_Jinkela_buffer_3131 (
        .din(new_Jinkela_wire_3569),
        .dout(new_Jinkela_wire_3570)
    );

    bfr new_Jinkela_buffer_2171 (
        .din(new_Jinkela_wire_2545),
        .dout(new_Jinkela_wire_2546)
    );

    bfr new_Jinkela_buffer_3075 (
        .din(new_Jinkela_wire_3504),
        .dout(new_Jinkela_wire_3505)
    );

    bfr new_Jinkela_buffer_6441 (
        .din(new_Jinkela_wire_7867),
        .dout(new_Jinkela_wire_7868)
    );

    bfr new_Jinkela_buffer_7362 (
        .din(n_0322_),
        .dout(new_Jinkela_wire_9157)
    );

    bfr new_Jinkela_buffer_7321 (
        .din(new_Jinkela_wire_9084),
        .dout(new_Jinkela_wire_9085)
    );

    spl2 new_Jinkela_splitter_571 (
        .a(n_0057_),
        .b(new_Jinkela_wire_7951),
        .c(new_Jinkela_wire_7953)
    );

    bfr new_Jinkela_buffer_2342 (
        .din(new_Jinkela_wire_2733),
        .dout(new_Jinkela_wire_2734)
    );

    bfr new_Jinkela_buffer_3140 (
        .din(n_1149_),
        .dout(new_Jinkela_wire_3590)
    );

    bfr new_Jinkela_buffer_2172 (
        .din(new_Jinkela_wire_2546),
        .dout(new_Jinkela_wire_2547)
    );

    bfr new_Jinkela_buffer_3076 (
        .din(new_Jinkela_wire_3505),
        .dout(new_Jinkela_wire_3506)
    );

    bfr new_Jinkela_buffer_6442 (
        .din(new_Jinkela_wire_7868),
        .dout(new_Jinkela_wire_7869)
    );

    bfr new_Jinkela_buffer_7352 (
        .din(new_Jinkela_wire_9128),
        .dout(new_Jinkela_wire_9129)
    );

    bfr new_Jinkela_buffer_7322 (
        .din(new_Jinkela_wire_9085),
        .dout(new_Jinkela_wire_9086)
    );

    bfr new_Jinkela_buffer_2219 (
        .din(new_Jinkela_wire_2605),
        .dout(new_Jinkela_wire_2606)
    );

    bfr new_Jinkela_buffer_3132 (
        .din(new_Jinkela_wire_3570),
        .dout(new_Jinkela_wire_3571)
    );

    bfr new_Jinkela_buffer_6497 (
        .din(new_Jinkela_wire_7938),
        .dout(new_Jinkela_wire_7939)
    );

    bfr new_Jinkela_buffer_3077 (
        .din(new_Jinkela_wire_3506),
        .dout(new_Jinkela_wire_3507)
    );

    bfr new_Jinkela_buffer_6443 (
        .din(new_Jinkela_wire_7869),
        .dout(new_Jinkela_wire_7870)
    );

    spl3L new_Jinkela_splitter_718 (
        .a(n_0918_),
        .d(new_Jinkela_wire_9150),
        .b(new_Jinkela_wire_9151),
        .c(new_Jinkela_wire_9152)
    );

    spl2 new_Jinkela_splitter_707 (
        .a(new_Jinkela_wire_9086),
        .b(new_Jinkela_wire_9087),
        .c(new_Jinkela_wire_9088)
    );

    bfr new_Jinkela_buffer_2220 (
        .din(new_Jinkela_wire_2606),
        .dout(new_Jinkela_wire_2607)
    );

    spl2 new_Jinkela_splitter_155 (
        .a(new_net_0),
        .b(new_Jinkela_wire_3610),
        .c(new_Jinkela_wire_3611)
    );

    bfr new_Jinkela_buffer_2280 (
        .din(new_Jinkela_wire_2668),
        .dout(new_Jinkela_wire_2669)
    );

    bfr new_Jinkela_buffer_3078 (
        .din(new_Jinkela_wire_3507),
        .dout(new_Jinkela_wire_3508)
    );

    bfr new_Jinkela_buffer_6444 (
        .din(new_Jinkela_wire_7870),
        .dout(new_Jinkela_wire_7871)
    );

    spl4L new_Jinkela_splitter_572 (
        .a(new_Jinkela_wire_7953),
        .d(new_Jinkela_wire_7954),
        .b(new_Jinkela_wire_7955),
        .e(new_Jinkela_wire_7956),
        .c(new_Jinkela_wire_7957)
    );

    bfr new_Jinkela_buffer_2221 (
        .din(new_Jinkela_wire_2607),
        .dout(new_Jinkela_wire_2608)
    );

    bfr new_Jinkela_buffer_3133 (
        .din(new_Jinkela_wire_3571),
        .dout(new_Jinkela_wire_3572)
    );

    bfr new_Jinkela_buffer_7353 (
        .din(new_Jinkela_wire_9129),
        .dout(new_Jinkela_wire_9130)
    );

    bfr new_Jinkela_buffer_2343 (
        .din(new_Jinkela_wire_2734),
        .dout(new_Jinkela_wire_2735)
    );

    bfr new_Jinkela_buffer_3079 (
        .din(new_Jinkela_wire_3508),
        .dout(new_Jinkela_wire_3509)
    );

    bfr new_Jinkela_buffer_6445 (
        .din(new_Jinkela_wire_7871),
        .dout(new_Jinkela_wire_7872)
    );

    spl2 new_Jinkela_splitter_719 (
        .a(new_Jinkela_wire_9152),
        .b(new_Jinkela_wire_9153),
        .c(new_Jinkela_wire_9154)
    );

    bfr new_Jinkela_buffer_7354 (
        .din(new_Jinkela_wire_9130),
        .dout(new_Jinkela_wire_9131)
    );

    bfr new_Jinkela_buffer_6498 (
        .din(new_Jinkela_wire_7939),
        .dout(new_Jinkela_wire_7940)
    );

    bfr new_Jinkela_buffer_2222 (
        .din(new_Jinkela_wire_2608),
        .dout(new_Jinkela_wire_2609)
    );

    spl3L new_Jinkela_splitter_154 (
        .a(n_0010_),
        .d(new_Jinkela_wire_3593),
        .b(new_Jinkela_wire_3594),
        .c(new_Jinkela_wire_3595)
    );

    bfr new_Jinkela_buffer_3967 (
        .din(n_0636_),
        .dout(new_Jinkela_wire_4656)
    );

    bfr new_Jinkela_buffer_3915 (
        .din(new_Jinkela_wire_4585),
        .dout(new_Jinkela_wire_4586)
    );

    bfr new_Jinkela_buffer_3963 (
        .din(new_Jinkela_wire_4639),
        .dout(new_Jinkela_wire_4640)
    );

    bfr new_Jinkela_buffer_3916 (
        .din(new_Jinkela_wire_4586),
        .dout(new_Jinkela_wire_4587)
    );

    spl2 new_Jinkela_splitter_255 (
        .a(n_0715_),
        .b(new_Jinkela_wire_4663),
        .c(new_Jinkela_wire_4664)
    );

    bfr new_Jinkela_buffer_3917 (
        .din(new_Jinkela_wire_4587),
        .dout(new_Jinkela_wire_4588)
    );

    bfr new_Jinkela_buffer_3964 (
        .din(new_Jinkela_wire_4640),
        .dout(new_Jinkela_wire_4641)
    );

    bfr new_Jinkela_buffer_3918 (
        .din(new_Jinkela_wire_4588),
        .dout(new_Jinkela_wire_4589)
    );

    bfr new_Jinkela_buffer_3919 (
        .din(new_Jinkela_wire_4589),
        .dout(new_Jinkela_wire_4590)
    );

    spl2 new_Jinkela_splitter_254 (
        .a(n_0710_),
        .b(new_Jinkela_wire_4661),
        .c(new_Jinkela_wire_4662)
    );

    bfr new_Jinkela_buffer_3965 (
        .din(new_Jinkela_wire_4641),
        .dout(new_Jinkela_wire_4642)
    );

    bfr new_Jinkela_buffer_3920 (
        .din(new_Jinkela_wire_4590),
        .dout(new_Jinkela_wire_4591)
    );

    bfr new_Jinkela_buffer_3968 (
        .din(new_Jinkela_wire_4656),
        .dout(new_Jinkela_wire_4657)
    );

    bfr new_Jinkela_buffer_3921 (
        .din(new_Jinkela_wire_4591),
        .dout(new_Jinkela_wire_4592)
    );

    bfr new_Jinkela_buffer_3970 (
        .din(n_0937_),
        .dout(new_Jinkela_wire_4665)
    );

    bfr new_Jinkela_buffer_3922 (
        .din(new_Jinkela_wire_4592),
        .dout(new_Jinkela_wire_4593)
    );

    bfr new_Jinkela_buffer_3969 (
        .din(new_Jinkela_wire_4657),
        .dout(new_Jinkela_wire_4658)
    );

    bfr new_Jinkela_buffer_3923 (
        .din(new_Jinkela_wire_4593),
        .dout(new_Jinkela_wire_4594)
    );

    spl2 new_Jinkela_splitter_256 (
        .a(n_0168_),
        .b(new_Jinkela_wire_4680),
        .c(new_Jinkela_wire_4681)
    );

    bfr new_Jinkela_buffer_3924 (
        .din(new_Jinkela_wire_4594),
        .dout(new_Jinkela_wire_4595)
    );

    spl2 new_Jinkela_splitter_253 (
        .a(new_Jinkela_wire_4658),
        .b(new_Jinkela_wire_4659),
        .c(new_Jinkela_wire_4660)
    );

    bfr new_Jinkela_buffer_3925 (
        .din(new_Jinkela_wire_4595),
        .dout(new_Jinkela_wire_4596)
    );

    bfr new_Jinkela_buffer_3926 (
        .din(new_Jinkela_wire_4596),
        .dout(new_Jinkela_wire_4597)
    );

    bfr new_Jinkela_buffer_3972 (
        .din(new_Jinkela_wire_4666),
        .dout(new_Jinkela_wire_4667)
    );

    bfr new_Jinkela_buffer_3927 (
        .din(new_Jinkela_wire_4597),
        .dout(new_Jinkela_wire_4598)
    );

    bfr new_Jinkela_buffer_3971 (
        .din(n_0544_),
        .dout(new_Jinkela_wire_4666)
    );

    bfr new_Jinkela_buffer_3928 (
        .din(new_Jinkela_wire_4598),
        .dout(new_Jinkela_wire_4599)
    );

    bfr new_Jinkela_buffer_4039 (
        .din(new_net_2568),
        .dout(new_Jinkela_wire_4738)
    );

    bfr new_Jinkela_buffer_3929 (
        .din(new_Jinkela_wire_4599),
        .dout(new_Jinkela_wire_4600)
    );

    bfr new_Jinkela_buffer_3973 (
        .din(new_Jinkela_wire_4667),
        .dout(new_Jinkela_wire_4668)
    );

    bfr new_Jinkela_buffer_3930 (
        .din(new_Jinkela_wire_4600),
        .dout(new_Jinkela_wire_4601)
    );

    spl2 new_Jinkela_splitter_258 (
        .a(n_1362_),
        .b(new_Jinkela_wire_4781),
        .c(new_Jinkela_wire_4782)
    );

    bfr new_Jinkela_buffer_3931 (
        .din(new_Jinkela_wire_4601),
        .dout(new_Jinkela_wire_4602)
    );

    bfr new_Jinkela_buffer_3974 (
        .din(new_Jinkela_wire_4668),
        .dout(new_Jinkela_wire_4669)
    );

    bfr new_Jinkela_buffer_3932 (
        .din(new_Jinkela_wire_4602),
        .dout(new_Jinkela_wire_4603)
    );

    bfr new_Jinkela_buffer_3985 (
        .din(new_Jinkela_wire_4681),
        .dout(new_Jinkela_wire_4682)
    );

    bfr new_Jinkela_buffer_4082 (
        .din(new_net_2533),
        .dout(new_Jinkela_wire_4783)
    );

    bfr new_Jinkela_buffer_3933 (
        .din(new_Jinkela_wire_4603),
        .dout(new_Jinkela_wire_4604)
    );

    bfr new_Jinkela_buffer_3975 (
        .din(new_Jinkela_wire_4669),
        .dout(new_Jinkela_wire_4670)
    );

    bfr new_Jinkela_buffer_3934 (
        .din(new_Jinkela_wire_4604),
        .dout(new_Jinkela_wire_4605)
    );

    bfr new_Jinkela_buffer_4040 (
        .din(new_Jinkela_wire_4738),
        .dout(new_Jinkela_wire_4739)
    );

    bfr new_Jinkela_buffer_3935 (
        .din(new_Jinkela_wire_4605),
        .dout(new_Jinkela_wire_4606)
    );

    bfr new_Jinkela_buffer_5634 (
        .din(new_Jinkela_wire_6754),
        .dout(new_Jinkela_wire_6755)
    );

    bfr new_Jinkela_buffer_5614 (
        .din(new_Jinkela_wire_6728),
        .dout(new_Jinkela_wire_6729)
    );

    spl3L new_Jinkela_splitter_443 (
        .a(n_0030_),
        .d(new_Jinkela_wire_6799),
        .b(new_Jinkela_wire_6800),
        .c(new_Jinkela_wire_6801)
    );

    bfr new_Jinkela_buffer_5615 (
        .din(new_Jinkela_wire_6729),
        .dout(new_Jinkela_wire_6730)
    );

    bfr new_Jinkela_buffer_5635 (
        .din(new_Jinkela_wire_6755),
        .dout(new_Jinkela_wire_6756)
    );

    bfr new_Jinkela_buffer_5616 (
        .din(new_Jinkela_wire_6730),
        .dout(new_Jinkela_wire_6731)
    );

    bfr new_Jinkela_buffer_5648 (
        .din(new_Jinkela_wire_6772),
        .dout(new_Jinkela_wire_6773)
    );

    bfr new_Jinkela_buffer_5617 (
        .din(new_Jinkela_wire_6731),
        .dout(new_Jinkela_wire_6732)
    );

    bfr new_Jinkela_buffer_5636 (
        .din(new_Jinkela_wire_6756),
        .dout(new_Jinkela_wire_6757)
    );

    bfr new_Jinkela_buffer_5618 (
        .din(new_Jinkela_wire_6732),
        .dout(new_Jinkela_wire_6733)
    );

    spl4L new_Jinkela_splitter_441 (
        .a(n_0040_),
        .d(new_Jinkela_wire_6792),
        .b(new_Jinkela_wire_6793),
        .e(new_Jinkela_wire_6794),
        .c(new_Jinkela_wire_6795)
    );

    bfr new_Jinkela_buffer_5657 (
        .din(n_0417_),
        .dout(new_Jinkela_wire_6791)
    );

    bfr new_Jinkela_buffer_5619 (
        .din(new_Jinkela_wire_6733),
        .dout(new_Jinkela_wire_6734)
    );

    bfr new_Jinkela_buffer_5637 (
        .din(new_Jinkela_wire_6757),
        .dout(new_Jinkela_wire_6758)
    );

    bfr new_Jinkela_buffer_5620 (
        .din(new_Jinkela_wire_6734),
        .dout(new_Jinkela_wire_6735)
    );

    bfr new_Jinkela_buffer_5649 (
        .din(new_Jinkela_wire_6773),
        .dout(new_Jinkela_wire_6774)
    );

    bfr new_Jinkela_buffer_5621 (
        .din(new_Jinkela_wire_6735),
        .dout(new_Jinkela_wire_6736)
    );

    bfr new_Jinkela_buffer_5638 (
        .din(new_Jinkela_wire_6758),
        .dout(new_Jinkela_wire_6759)
    );

    bfr new_Jinkela_buffer_5622 (
        .din(new_Jinkela_wire_6736),
        .dout(new_Jinkela_wire_6737)
    );

    bfr new_Jinkela_buffer_5658 (
        .din(new_Jinkela_wire_6795),
        .dout(new_Jinkela_wire_6796)
    );

    spl2 new_Jinkela_splitter_444 (
        .a(n_0264_),
        .b(new_Jinkela_wire_6804),
        .c(new_Jinkela_wire_6805)
    );

    bfr new_Jinkela_buffer_5623 (
        .din(new_Jinkela_wire_6737),
        .dout(new_Jinkela_wire_6738)
    );

    bfr new_Jinkela_buffer_5639 (
        .din(new_Jinkela_wire_6759),
        .dout(new_Jinkela_wire_6760)
    );

    bfr new_Jinkela_buffer_5624 (
        .din(new_Jinkela_wire_6738),
        .dout(new_Jinkela_wire_6739)
    );

    bfr new_Jinkela_buffer_5650 (
        .din(new_Jinkela_wire_6774),
        .dout(new_Jinkela_wire_6775)
    );

    bfr new_Jinkela_buffer_5625 (
        .din(new_Jinkela_wire_6739),
        .dout(new_Jinkela_wire_6740)
    );

    bfr new_Jinkela_buffer_5640 (
        .din(new_Jinkela_wire_6760),
        .dout(new_Jinkela_wire_6761)
    );

    bfr new_Jinkela_buffer_5626 (
        .din(new_Jinkela_wire_6740),
        .dout(new_Jinkela_wire_6741)
    );

    bfr new_Jinkela_buffer_5641 (
        .din(new_Jinkela_wire_6761),
        .dout(new_Jinkela_wire_6762)
    );

    bfr new_Jinkela_buffer_5651 (
        .din(new_Jinkela_wire_6775),
        .dout(new_Jinkela_wire_6776)
    );

    bfr new_Jinkela_buffer_5642 (
        .din(new_Jinkela_wire_6762),
        .dout(new_Jinkela_wire_6763)
    );

    bfr new_Jinkela_buffer_5643 (
        .din(new_Jinkela_wire_6763),
        .dout(new_Jinkela_wire_6764)
    );

    bfr new_Jinkela_buffer_5652 (
        .din(new_Jinkela_wire_6776),
        .dout(new_Jinkela_wire_6777)
    );

    spl2 new_Jinkela_splitter_435 (
        .a(new_Jinkela_wire_6764),
        .b(new_Jinkela_wire_6765),
        .c(new_Jinkela_wire_6766)
    );

    bfr new_Jinkela_buffer_5653 (
        .din(new_Jinkela_wire_6777),
        .dout(new_Jinkela_wire_6778)
    );

    spl3L new_Jinkela_splitter_445 (
        .a(n_1301_),
        .d(new_Jinkela_wire_6806),
        .b(new_Jinkela_wire_6807),
        .c(new_Jinkela_wire_6808)
    );

    bfr new_Jinkela_buffer_5659 (
        .din(new_Jinkela_wire_6801),
        .dout(new_Jinkela_wire_6802)
    );

    spl2 new_Jinkela_splitter_442 (
        .a(new_Jinkela_wire_6796),
        .b(new_Jinkela_wire_6797),
        .c(new_Jinkela_wire_6798)
    );

    spl2 new_Jinkela_splitter_437 (
        .a(new_Jinkela_wire_6778),
        .b(new_Jinkela_wire_6779),
        .c(new_Jinkela_wire_6780)
    );

    bfr new_Jinkela_buffer_5654 (
        .din(new_Jinkela_wire_6780),
        .dout(new_Jinkela_wire_6781)
    );

    bfr new_Jinkela_buffer_5666 (
        .din(n_0247_),
        .dout(new_Jinkela_wire_6814)
    );

    bfr new_Jinkela_buffer_5660 (
        .din(new_Jinkela_wire_6802),
        .dout(new_Jinkela_wire_6803)
    );

    bfr new_Jinkela_buffer_5655 (
        .din(new_Jinkela_wire_6781),
        .dout(new_Jinkela_wire_6782)
    );

    and_bi n_1695_ (
        .a(new_Jinkela_wire_1245),
        .b(new_Jinkela_wire_2739),
        .c(n_0962_)
    );

    or_bb n_2409_ (
        .a(new_Jinkela_wire_3711),
        .b(new_Jinkela_wire_6805),
        .c(n_0284_)
    );

    bfr new_Jinkela_buffer_4870 (
        .din(new_Jinkela_wire_5806),
        .dout(new_Jinkela_wire_5807)
    );

    bfr new_Jinkela_buffer_4770 (
        .din(new_Jinkela_wire_5697),
        .dout(new_Jinkela_wire_5698)
    );

    and_ii n_1696_ (
        .a(n_0962_),
        .b(n_0961_),
        .c(n_0963_)
    );

    and_bb n_2410_ (
        .a(new_Jinkela_wire_6821),
        .b(new_Jinkela_wire_6708),
        .c(n_0285_)
    );

    bfr new_Jinkela_buffer_4826 (
        .din(new_Jinkela_wire_5760),
        .dout(new_Jinkela_wire_5761)
    );

    and_ii n_1697_ (
        .a(new_Jinkela_wire_4008),
        .b(new_Jinkela_wire_6784),
        .c(n_0964_)
    );

    or_bb n_2411_ (
        .a(new_Jinkela_wire_5234),
        .b(new_Jinkela_wire_5637),
        .c(n_0286_)
    );

    bfr new_Jinkela_buffer_4809 (
        .din(new_Jinkela_wire_5740),
        .dout(new_Jinkela_wire_5741)
    );

    bfr new_Jinkela_buffer_4771 (
        .din(new_Jinkela_wire_5698),
        .dout(new_Jinkela_wire_5699)
    );

    and_bb n_1698_ (
        .a(new_Jinkela_wire_4007),
        .b(new_Jinkela_wire_6783),
        .c(n_0965_)
    );

    and_bi n_2412_ (
        .a(new_Jinkela_wire_3842),
        .b(new_Jinkela_wire_10485),
        .c(n_0287_)
    );

    and_ii n_1699_ (
        .a(n_0965_),
        .b(n_0964_),
        .c(n_0966_)
    );

    and_bi n_2413_ (
        .a(new_Jinkela_wire_10135),
        .b(new_Jinkela_wire_7926),
        .c(n_0288_)
    );

    bfr new_Jinkela_buffer_4772 (
        .din(new_Jinkela_wire_5699),
        .dout(new_Jinkela_wire_5700)
    );

    and_bi n_1700_ (
        .a(new_Jinkela_wire_6514),
        .b(new_Jinkela_wire_5558),
        .c(n_0967_)
    );

    or_bb n_2414_ (
        .a(new_Jinkela_wire_9542),
        .b(n_0287_),
        .c(n_0289_)
    );

    and_bi n_1701_ (
        .a(new_Jinkela_wire_5557),
        .b(new_Jinkela_wire_6513),
        .c(n_0968_)
    );

    or_bb n_2415_ (
        .a(new_Jinkela_wire_6902),
        .b(n_0285_),
        .c(n_0290_)
    );

    bfr new_Jinkela_buffer_4810 (
        .din(new_Jinkela_wire_5741),
        .dout(new_Jinkela_wire_5742)
    );

    bfr new_Jinkela_buffer_4773 (
        .din(new_Jinkela_wire_5700),
        .dout(new_Jinkela_wire_5701)
    );

    or_bb n_1702_ (
        .a(n_0968_),
        .b(n_0967_),
        .c(n_0969_)
    );

    and_bi n_2416_ (
        .a(n_0284_),
        .b(new_Jinkela_wire_3850),
        .c(n_0291_)
    );

    and_bi n_1703_ (
        .a(new_Jinkela_wire_95),
        .b(new_Jinkela_wire_1170),
        .c(n_0970_)
    );

    and_bi n_2417_ (
        .a(new_Jinkela_wire_6312),
        .b(new_Jinkela_wire_7095),
        .c(n_0292_)
    );

    bfr new_Jinkela_buffer_4774 (
        .din(new_Jinkela_wire_5701),
        .dout(new_Jinkela_wire_5702)
    );

    and_bi n_1704_ (
        .a(new_Jinkela_wire_1317),
        .b(new_Jinkela_wire_2169),
        .c(n_0971_)
    );

    and_bi n_2418_ (
        .a(new_Jinkela_wire_9473),
        .b(new_Jinkela_wire_9546),
        .c(n_0293_)
    );

    bfr new_Jinkela_buffer_4827 (
        .din(new_Jinkela_wire_5761),
        .dout(new_Jinkela_wire_5762)
    );

    and_ii n_1705_ (
        .a(n_0971_),
        .b(n_0970_),
        .c(n_0972_)
    );

    or_bb n_2419_ (
        .a(n_0293_),
        .b(n_0292_),
        .c(n_0294_)
    );

    bfr new_Jinkela_buffer_4811 (
        .din(new_Jinkela_wire_5742),
        .dout(new_Jinkela_wire_5743)
    );

    bfr new_Jinkela_buffer_4775 (
        .din(new_Jinkela_wire_5702),
        .dout(new_Jinkela_wire_5703)
    );

    and_bi n_1706_ (
        .a(new_Jinkela_wire_3201),
        .b(new_Jinkela_wire_1279),
        .c(n_0973_)
    );

    and_bi n_2420_ (
        .a(new_Jinkela_wire_7096),
        .b(new_Jinkela_wire_6313),
        .c(n_0295_)
    );

    and_bi n_1707_ (
        .a(new_Jinkela_wire_1182),
        .b(new_Jinkela_wire_695),
        .c(n_0974_)
    );

    and_bi n_2421_ (
        .a(new_Jinkela_wire_9547),
        .b(new_Jinkela_wire_9474),
        .c(n_0296_)
    );

    bfr new_Jinkela_buffer_4776 (
        .din(new_Jinkela_wire_5703),
        .dout(new_Jinkela_wire_5704)
    );

    and_ii n_1708_ (
        .a(n_0974_),
        .b(n_0973_),
        .c(n_0975_)
    );

    and_ii n_2422_ (
        .a(new_Jinkela_wire_6013),
        .b(new_Jinkela_wire_9485),
        .c(n_0297_)
    );

    and_bi n_1709_ (
        .a(new_Jinkela_wire_6399),
        .b(new_Jinkela_wire_6009),
        .c(n_0976_)
    );

    and_bi n_2423_ (
        .a(n_0297_),
        .b(new_Jinkela_wire_4015),
        .c(n_0298_)
    );

    bfr new_Jinkela_buffer_4812 (
        .din(new_Jinkela_wire_5743),
        .dout(new_Jinkela_wire_5744)
    );

    bfr new_Jinkela_buffer_4777 (
        .din(new_Jinkela_wire_5704),
        .dout(new_Jinkela_wire_5705)
    );

    and_bi n_1710_ (
        .a(new_Jinkela_wire_6008),
        .b(new_Jinkela_wire_6398),
        .c(n_0977_)
    );

    and_bi n_2424_ (
        .a(new_Jinkela_wire_4085),
        .b(new_Jinkela_wire_8400),
        .c(n_0299_)
    );

    and_ii n_1711_ (
        .a(n_0977_),
        .b(n_0976_),
        .c(n_0978_)
    );

    and_bi n_2425_ (
        .a(new_Jinkela_wire_10562),
        .b(new_Jinkela_wire_7250),
        .c(n_0300_)
    );

    bfr new_Jinkela_buffer_4871 (
        .din(new_Jinkela_wire_5807),
        .dout(new_Jinkela_wire_5808)
    );

    bfr new_Jinkela_buffer_4778 (
        .din(new_Jinkela_wire_5705),
        .dout(new_Jinkela_wire_5706)
    );

    and_bi n_1712_ (
        .a(new_Jinkela_wire_3358),
        .b(new_Jinkela_wire_1188),
        .c(n_0979_)
    );

    and_ii n_2426_ (
        .a(n_0300_),
        .b(n_0299_),
        .c(n_0301_)
    );

    bfr new_Jinkela_buffer_4828 (
        .din(new_Jinkela_wire_5762),
        .dout(new_Jinkela_wire_5763)
    );

    and_bi n_1713_ (
        .a(new_Jinkela_wire_1352),
        .b(new_Jinkela_wire_1475),
        .c(n_0980_)
    );

    and_bi n_2427_ (
        .a(new_Jinkela_wire_8399),
        .b(new_Jinkela_wire_4086),
        .c(n_0302_)
    );

    bfr new_Jinkela_buffer_4813 (
        .din(new_Jinkela_wire_5744),
        .dout(new_Jinkela_wire_5745)
    );

    bfr new_Jinkela_buffer_4779 (
        .din(new_Jinkela_wire_5706),
        .dout(new_Jinkela_wire_5707)
    );

    and_ii n_1714_ (
        .a(n_0980_),
        .b(n_0979_),
        .c(n_0981_)
    );

    and_bi n_2428_ (
        .a(new_Jinkela_wire_7249),
        .b(new_Jinkela_wire_10561),
        .c(n_0303_)
    );

    and_ii n_2429_ (
        .a(new_Jinkela_wire_6247),
        .b(new_Jinkela_wire_8850),
        .c(n_0304_)
    );

    and_bi n_1715_ (
        .a(new_Jinkela_wire_8302),
        .b(new_Jinkela_wire_8933),
        .c(n_0982_)
    );

    bfr new_Jinkela_buffer_4780 (
        .din(new_Jinkela_wire_5707),
        .dout(new_Jinkela_wire_5708)
    );

    and_bi n_1716_ (
        .a(new_Jinkela_wire_8932),
        .b(new_Jinkela_wire_8301),
        .c(n_0983_)
    );

    and_bb n_2430_ (
        .a(n_0304_),
        .b(new_Jinkela_wire_3589),
        .c(n_0305_)
    );

    or_bb n_1717_ (
        .a(n_0983_),
        .b(n_0982_),
        .c(n_0984_)
    );

    or_ii n_2431_ (
        .a(new_Jinkela_wire_7542),
        .b(new_Jinkela_wire_4859),
        .c(n_0306_)
    );

    bfr new_Jinkela_buffer_4814 (
        .din(new_Jinkela_wire_5745),
        .dout(new_Jinkela_wire_5746)
    );

    bfr new_Jinkela_buffer_4781 (
        .din(new_Jinkela_wire_5708),
        .dout(new_Jinkela_wire_5709)
    );

    and_bi n_1718_ (
        .a(new_Jinkela_wire_3120),
        .b(new_Jinkela_wire_1205),
        .c(n_0985_)
    );

    or_bb n_2432_ (
        .a(new_Jinkela_wire_5411),
        .b(n_0291_),
        .c(n_0307_)
    );

    and_bi n_1719_ (
        .a(new_Jinkela_wire_1225),
        .b(new_Jinkela_wire_275),
        .c(n_0986_)
    );

    or_bb n_2433_ (
        .a(new_Jinkela_wire_8852),
        .b(new_Jinkela_wire_3588),
        .c(n_0308_)
    );

    bfr new_Jinkela_buffer_4782 (
        .din(new_Jinkela_wire_5709),
        .dout(new_Jinkela_wire_5710)
    );

    and_bi n_2434_ (
        .a(new_Jinkela_wire_4858),
        .b(new_Jinkela_wire_5281),
        .c(n_0309_)
    );

    and_ii n_1720_ (
        .a(n_0986_),
        .b(n_0985_),
        .c(n_0987_)
    );

    bfr new_Jinkela_buffer_4829 (
        .din(new_Jinkela_wire_5763),
        .dout(new_Jinkela_wire_5764)
    );

    and_bi n_1721_ (
        .a(new_Jinkela_wire_1903),
        .b(new_Jinkela_wire_1202),
        .c(n_0988_)
    );

    and_bi n_2435_ (
        .a(new_Jinkela_wire_4014),
        .b(new_Jinkela_wire_6015),
        .c(n_0310_)
    );

    bfr new_Jinkela_buffer_4815 (
        .din(new_Jinkela_wire_5746),
        .dout(new_Jinkela_wire_5747)
    );

    bfr new_Jinkela_buffer_4783 (
        .din(new_Jinkela_wire_5710),
        .dout(new_Jinkela_wire_5711)
    );

    and_bi n_1722_ (
        .a(new_Jinkela_wire_1351),
        .b(new_Jinkela_wire_3275),
        .c(n_0989_)
    );

    or_bb n_2436_ (
        .a(new_Jinkela_wire_5501),
        .b(n_0309_),
        .c(n_0311_)
    );

    and_ii n_1723_ (
        .a(n_0989_),
        .b(n_0988_),
        .c(n_0990_)
    );

    and_bi n_2437_ (
        .a(n_0307_),
        .b(new_Jinkela_wire_7199),
        .c(n_0312_)
    );

    bfr new_Jinkela_buffer_4784 (
        .din(new_Jinkela_wire_5711),
        .dout(new_Jinkela_wire_5712)
    );

    and_bi n_1724_ (
        .a(new_Jinkela_wire_1782),
        .b(new_Jinkela_wire_1377),
        .c(n_0991_)
    );

    and_bi n_2438_ (
        .a(new_Jinkela_wire_7203),
        .b(new_Jinkela_wire_7843),
        .c(n_0313_)
    );

    bfr new_Jinkela_buffer_4934 (
        .din(n_1234_),
        .dout(new_Jinkela_wire_5882)
    );

    and_bi n_1725_ (
        .a(new_Jinkela_wire_1374),
        .b(new_Jinkela_wire_3053),
        .c(n_0992_)
    );

    and_bb n_2439_ (
        .a(new_Jinkela_wire_9601),
        .b(new_Jinkela_wire_9153),
        .c(n_0314_)
    );

    bfr new_Jinkela_buffer_4816 (
        .din(new_Jinkela_wire_5747),
        .dout(new_Jinkela_wire_5748)
    );

    bfr new_Jinkela_buffer_4785 (
        .din(new_Jinkela_wire_5712),
        .dout(new_Jinkela_wire_5713)
    );

    and_ii n_1726_ (
        .a(n_0992_),
        .b(n_0991_),
        .c(n_0993_)
    );

    and_ii n_2440_ (
        .a(new_Jinkela_wire_9602),
        .b(new_Jinkela_wire_9154),
        .c(n_0315_)
    );

    and_ii n_1727_ (
        .a(new_Jinkela_wire_9537),
        .b(new_Jinkela_wire_8286),
        .c(n_0994_)
    );

    or_bb n_2441_ (
        .a(new_Jinkela_wire_6707),
        .b(new_Jinkela_wire_8571),
        .c(n_0316_)
    );

    bfr new_Jinkela_buffer_4872 (
        .din(new_Jinkela_wire_5808),
        .dout(new_Jinkela_wire_5809)
    );

    bfr new_Jinkela_buffer_4786 (
        .din(new_Jinkela_wire_5713),
        .dout(new_Jinkela_wire_5714)
    );

    and_bb n_1728_ (
        .a(new_Jinkela_wire_9536),
        .b(new_Jinkela_wire_8285),
        .c(n_0995_)
    );

    and_bi n_2442_ (
        .a(new_Jinkela_wire_7308),
        .b(new_Jinkela_wire_10559),
        .c(n_0317_)
    );

    bfr new_Jinkela_buffer_4830 (
        .din(new_Jinkela_wire_5764),
        .dout(new_Jinkela_wire_5765)
    );

    or_bb n_1729_ (
        .a(n_0995_),
        .b(n_0994_),
        .c(n_0996_)
    );

    and_bi n_2443_ (
        .a(new_Jinkela_wire_10560),
        .b(new_Jinkela_wire_7307),
        .c(n_0318_)
    );

    bfr new_Jinkela_buffer_4817 (
        .din(new_Jinkela_wire_5748),
        .dout(new_Jinkela_wire_5749)
    );

    bfr new_Jinkela_buffer_4787 (
        .din(new_Jinkela_wire_5714),
        .dout(new_Jinkela_wire_5715)
    );

    or_bb n_1730_ (
        .a(new_Jinkela_wire_5011),
        .b(new_Jinkela_wire_8198),
        .c(n_0997_)
    );

    or_bb n_2444_ (
        .a(new_Jinkela_wire_5730),
        .b(new_Jinkela_wire_3727),
        .c(n_0319_)
    );

    or_ii n_1731_ (
        .a(new_Jinkela_wire_5010),
        .b(new_Jinkela_wire_8197),
        .c(n_0998_)
    );

    or_bb n_2445_ (
        .a(n_0319_),
        .b(n_0316_),
        .c(n_0320_)
    );

    bfr new_Jinkela_buffer_4788 (
        .din(new_Jinkela_wire_5715),
        .dout(new_Jinkela_wire_5716)
    );

    and_bb n_1732_ (
        .a(n_0998_),
        .b(n_0997_),
        .c(n_0999_)
    );

    and_ii n_2446_ (
        .a(n_0320_),
        .b(new_Jinkela_wire_8395),
        .c(n_0321_)
    );

    and_bi n_1733_ (
        .a(new_Jinkela_wire_7460),
        .b(new_Jinkela_wire_10418),
        .c(n_1000_)
    );

    and_ii n_2447_ (
        .a(new_Jinkela_wire_8766),
        .b(new_Jinkela_wire_9466),
        .c(n_0322_)
    );

    bfr new_Jinkela_buffer_4818 (
        .din(new_Jinkela_wire_5749),
        .dout(new_Jinkela_wire_5750)
    );

    bfr new_Jinkela_buffer_4789 (
        .din(new_Jinkela_wire_5716),
        .dout(new_Jinkela_wire_5717)
    );

    and_bi n_1734_ (
        .a(new_Jinkela_wire_10417),
        .b(new_Jinkela_wire_7459),
        .c(n_1001_)
    );

    and_bi n_2448_ (
        .a(new_Jinkela_wire_7744),
        .b(new_Jinkela_wire_9753),
        .c(n_0323_)
    );

    or_bb n_2449_ (
        .a(n_0323_),
        .b(new_Jinkela_wire_9157),
        .c(n_0324_)
    );

    and_ii n_1735_ (
        .a(n_1001_),
        .b(n_1000_),
        .c(n_1002_)
    );

    spl3L new_Jinkela_splitter_360 (
        .a(n_0000_),
        .d(new_Jinkela_wire_5879),
        .b(new_Jinkela_wire_5880),
        .c(new_Jinkela_wire_5881)
    );

    bfr new_Jinkela_buffer_4790 (
        .din(new_Jinkela_wire_5717),
        .dout(new_Jinkela_wire_5718)
    );

    and_bb n_2450_ (
        .a(new_Jinkela_wire_8763),
        .b(new_Jinkela_wire_9467),
        .c(n_0325_)
    );

    or_bb n_1736_ (
        .a(new_Jinkela_wire_8297),
        .b(new_Jinkela_wire_4431),
        .c(n_1003_)
    );

    bfr new_Jinkela_buffer_6509 (
        .din(new_Jinkela_wire_7951),
        .dout(new_Jinkela_wire_7952)
    );

    bfr new_Jinkela_buffer_3976 (
        .din(new_Jinkela_wire_4670),
        .dout(new_Jinkela_wire_4671)
    );

    bfr new_Jinkela_buffer_6446 (
        .din(new_Jinkela_wire_7872),
        .dout(new_Jinkela_wire_7873)
    );

    bfr new_Jinkela_buffer_3936 (
        .din(new_Jinkela_wire_4606),
        .dout(new_Jinkela_wire_4607)
    );

    spl2 new_Jinkela_splitter_574 (
        .a(n_0118_),
        .b(new_Jinkela_wire_7990),
        .c(new_Jinkela_wire_7991)
    );

    bfr new_Jinkela_buffer_6499 (
        .din(new_Jinkela_wire_7940),
        .dout(new_Jinkela_wire_7941)
    );

    bfr new_Jinkela_buffer_3986 (
        .din(new_Jinkela_wire_4682),
        .dout(new_Jinkela_wire_4683)
    );

    bfr new_Jinkela_buffer_6447 (
        .din(new_Jinkela_wire_7873),
        .dout(new_Jinkela_wire_7874)
    );

    bfr new_Jinkela_buffer_3937 (
        .din(new_Jinkela_wire_4607),
        .dout(new_Jinkela_wire_4608)
    );

    bfr new_Jinkela_buffer_3977 (
        .din(new_Jinkela_wire_4671),
        .dout(new_Jinkela_wire_4672)
    );

    bfr new_Jinkela_buffer_6448 (
        .din(new_Jinkela_wire_7874),
        .dout(new_Jinkela_wire_7875)
    );

    bfr new_Jinkela_buffer_3938 (
        .din(new_Jinkela_wire_4608),
        .dout(new_Jinkela_wire_4609)
    );

    bfr new_Jinkela_buffer_6500 (
        .din(new_Jinkela_wire_7941),
        .dout(new_Jinkela_wire_7942)
    );

    spl2 new_Jinkela_splitter_260 (
        .a(n_0166_),
        .b(new_Jinkela_wire_4854),
        .c(new_Jinkela_wire_4855)
    );

    bfr new_Jinkela_buffer_6449 (
        .din(new_Jinkela_wire_7875),
        .dout(new_Jinkela_wire_7876)
    );

    bfr new_Jinkela_buffer_3939 (
        .din(new_Jinkela_wire_4609),
        .dout(new_Jinkela_wire_4610)
    );

    bfr new_Jinkela_buffer_6510 (
        .din(new_Jinkela_wire_7957),
        .dout(new_Jinkela_wire_7958)
    );

    bfr new_Jinkela_buffer_3978 (
        .din(new_Jinkela_wire_4672),
        .dout(new_Jinkela_wire_4673)
    );

    bfr new_Jinkela_buffer_6450 (
        .din(new_Jinkela_wire_7876),
        .dout(new_Jinkela_wire_7877)
    );

    bfr new_Jinkela_buffer_3940 (
        .din(new_Jinkela_wire_4610),
        .dout(new_Jinkela_wire_4611)
    );

    bfr new_Jinkela_buffer_6501 (
        .din(new_Jinkela_wire_7942),
        .dout(new_Jinkela_wire_7943)
    );

    bfr new_Jinkela_buffer_3987 (
        .din(new_Jinkela_wire_4683),
        .dout(new_Jinkela_wire_4684)
    );

    bfr new_Jinkela_buffer_6451 (
        .din(new_Jinkela_wire_7877),
        .dout(new_Jinkela_wire_7878)
    );

    bfr new_Jinkela_buffer_3941 (
        .din(new_Jinkela_wire_4611),
        .dout(new_Jinkela_wire_4612)
    );

    bfr new_Jinkela_buffer_3979 (
        .din(new_Jinkela_wire_4673),
        .dout(new_Jinkela_wire_4674)
    );

    bfr new_Jinkela_buffer_6452 (
        .din(new_Jinkela_wire_7878),
        .dout(new_Jinkela_wire_7879)
    );

    bfr new_Jinkela_buffer_3942 (
        .din(new_Jinkela_wire_4612),
        .dout(new_Jinkela_wire_4613)
    );

    bfr new_Jinkela_buffer_6538 (
        .din(new_Jinkela_wire_7985),
        .dout(new_Jinkela_wire_7986)
    );

    bfr new_Jinkela_buffer_6502 (
        .din(new_Jinkela_wire_7943),
        .dout(new_Jinkela_wire_7944)
    );

    bfr new_Jinkela_buffer_4041 (
        .din(new_Jinkela_wire_4739),
        .dout(new_Jinkela_wire_4740)
    );

    bfr new_Jinkela_buffer_6453 (
        .din(new_Jinkela_wire_7879),
        .dout(new_Jinkela_wire_7880)
    );

    bfr new_Jinkela_buffer_3943 (
        .din(new_Jinkela_wire_4613),
        .dout(new_Jinkela_wire_4614)
    );

    bfr new_Jinkela_buffer_3980 (
        .din(new_Jinkela_wire_4674),
        .dout(new_Jinkela_wire_4675)
    );

    bfr new_Jinkela_buffer_6454 (
        .din(new_Jinkela_wire_7880),
        .dout(new_Jinkela_wire_7881)
    );

    bfr new_Jinkela_buffer_3944 (
        .din(new_Jinkela_wire_4614),
        .dout(new_Jinkela_wire_4615)
    );

    bfr new_Jinkela_buffer_6503 (
        .din(new_Jinkela_wire_7944),
        .dout(new_Jinkela_wire_7945)
    );

    bfr new_Jinkela_buffer_3988 (
        .din(new_Jinkela_wire_4684),
        .dout(new_Jinkela_wire_4685)
    );

    bfr new_Jinkela_buffer_6455 (
        .din(new_Jinkela_wire_7881),
        .dout(new_Jinkela_wire_7882)
    );

    bfr new_Jinkela_buffer_3945 (
        .din(new_Jinkela_wire_4615),
        .dout(new_Jinkela_wire_4616)
    );

    bfr new_Jinkela_buffer_6511 (
        .din(new_Jinkela_wire_7958),
        .dout(new_Jinkela_wire_7959)
    );

    bfr new_Jinkela_buffer_3981 (
        .din(new_Jinkela_wire_4675),
        .dout(new_Jinkela_wire_4676)
    );

    bfr new_Jinkela_buffer_6456 (
        .din(new_Jinkela_wire_7882),
        .dout(new_Jinkela_wire_7883)
    );

    bfr new_Jinkela_buffer_3946 (
        .din(new_Jinkela_wire_4616),
        .dout(new_Jinkela_wire_4617)
    );

    bfr new_Jinkela_buffer_6504 (
        .din(new_Jinkela_wire_7945),
        .dout(new_Jinkela_wire_7946)
    );

    bfr new_Jinkela_buffer_4083 (
        .din(new_Jinkela_wire_4783),
        .dout(new_Jinkela_wire_4784)
    );

    bfr new_Jinkela_buffer_6457 (
        .din(new_Jinkela_wire_7883),
        .dout(new_Jinkela_wire_7884)
    );

    bfr new_Jinkela_buffer_3947 (
        .din(new_Jinkela_wire_4617),
        .dout(new_Jinkela_wire_4618)
    );

    bfr new_Jinkela_buffer_6539 (
        .din(new_Jinkela_wire_7986),
        .dout(new_Jinkela_wire_7987)
    );

    bfr new_Jinkela_buffer_3982 (
        .din(new_Jinkela_wire_4676),
        .dout(new_Jinkela_wire_4677)
    );

    bfr new_Jinkela_buffer_6458 (
        .din(new_Jinkela_wire_7884),
        .dout(new_Jinkela_wire_7885)
    );

    bfr new_Jinkela_buffer_3948 (
        .din(new_Jinkela_wire_4618),
        .dout(new_Jinkela_wire_4619)
    );

    spl3L new_Jinkela_splitter_575 (
        .a(n_0694_),
        .d(new_Jinkela_wire_7992),
        .b(new_Jinkela_wire_7993),
        .c(new_Jinkela_wire_7994)
    );

    bfr new_Jinkela_buffer_6505 (
        .din(new_Jinkela_wire_7946),
        .dout(new_Jinkela_wire_7947)
    );

    bfr new_Jinkela_buffer_3989 (
        .din(new_Jinkela_wire_4685),
        .dout(new_Jinkela_wire_4686)
    );

    bfr new_Jinkela_buffer_6459 (
        .din(new_Jinkela_wire_7885),
        .dout(new_Jinkela_wire_7886)
    );

    bfr new_Jinkela_buffer_3949 (
        .din(new_Jinkela_wire_4619),
        .dout(new_Jinkela_wire_4620)
    );

    bfr new_Jinkela_buffer_6512 (
        .din(new_Jinkela_wire_7959),
        .dout(new_Jinkela_wire_7960)
    );

    bfr new_Jinkela_buffer_3983 (
        .din(new_Jinkela_wire_4677),
        .dout(new_Jinkela_wire_4678)
    );

    bfr new_Jinkela_buffer_6460 (
        .din(new_Jinkela_wire_7886),
        .dout(new_Jinkela_wire_7887)
    );

    bfr new_Jinkela_buffer_3950 (
        .din(new_Jinkela_wire_4620),
        .dout(new_Jinkela_wire_4621)
    );

    bfr new_Jinkela_buffer_6506 (
        .din(new_Jinkela_wire_7947),
        .dout(new_Jinkela_wire_7948)
    );

    bfr new_Jinkela_buffer_4042 (
        .din(new_Jinkela_wire_4740),
        .dout(new_Jinkela_wire_4741)
    );

    bfr new_Jinkela_buffer_6461 (
        .din(new_Jinkela_wire_7887),
        .dout(new_Jinkela_wire_7888)
    );

    bfr new_Jinkela_buffer_3951 (
        .din(new_Jinkela_wire_4621),
        .dout(new_Jinkela_wire_4622)
    );

    bfr new_Jinkela_buffer_7307 (
        .din(new_Jinkela_wire_9070),
        .dout(new_Jinkela_wire_9071)
    );

    bfr new_Jinkela_buffer_3984 (
        .din(new_Jinkela_wire_4678),
        .dout(new_Jinkela_wire_4679)
    );

    bfr new_Jinkela_buffer_6462 (
        .din(new_Jinkela_wire_7888),
        .dout(new_Jinkela_wire_7889)
    );

    bfr new_Jinkela_buffer_3952 (
        .din(new_Jinkela_wire_4622),
        .dout(new_Jinkela_wire_4623)
    );

    bfr new_Jinkela_buffer_6540 (
        .din(n_1247_),
        .dout(new_Jinkela_wire_7997)
    );

    bfr new_Jinkela_buffer_6507 (
        .din(new_Jinkela_wire_7948),
        .dout(new_Jinkela_wire_7949)
    );

    bfr new_Jinkela_buffer_3990 (
        .din(new_Jinkela_wire_4686),
        .dout(new_Jinkela_wire_4687)
    );

    bfr new_Jinkela_buffer_6463 (
        .din(new_Jinkela_wire_7889),
        .dout(new_Jinkela_wire_7890)
    );

    bfr new_Jinkela_buffer_3953 (
        .din(new_Jinkela_wire_4623),
        .dout(new_Jinkela_wire_4624)
    );

    bfr new_Jinkela_buffer_6513 (
        .din(new_Jinkela_wire_7960),
        .dout(new_Jinkela_wire_7961)
    );

    bfr new_Jinkela_buffer_4117 (
        .din(new_net_7),
        .dout(new_Jinkela_wire_4818)
    );

    bfr new_Jinkela_buffer_6464 (
        .din(new_Jinkela_wire_7890),
        .dout(new_Jinkela_wire_7891)
    );

    bfr new_Jinkela_buffer_3954 (
        .din(new_Jinkela_wire_4624),
        .dout(new_Jinkela_wire_4625)
    );

    bfr new_Jinkela_buffer_6508 (
        .din(new_Jinkela_wire_7949),
        .dout(new_Jinkela_wire_7950)
    );

    bfr new_Jinkela_buffer_3991 (
        .din(new_Jinkela_wire_4687),
        .dout(new_Jinkela_wire_4688)
    );

    bfr new_Jinkela_buffer_6465 (
        .din(new_Jinkela_wire_7891),
        .dout(new_Jinkela_wire_7892)
    );

    bfr new_Jinkela_buffer_3955 (
        .din(new_Jinkela_wire_4625),
        .dout(new_Jinkela_wire_4626)
    );

    spl2 new_Jinkela_splitter_576 (
        .a(n_0158_),
        .b(new_Jinkela_wire_7995),
        .c(new_Jinkela_wire_7996)
    );

    bfr new_Jinkela_buffer_4043 (
        .din(new_Jinkela_wire_4741),
        .dout(new_Jinkela_wire_4742)
    );

    bfr new_Jinkela_buffer_6466 (
        .din(new_Jinkela_wire_7892),
        .dout(new_Jinkela_wire_7893)
    );

    bfr new_Jinkela_buffer_3992 (
        .din(new_Jinkela_wire_4688),
        .dout(new_Jinkela_wire_4689)
    );

    spl2 new_Jinkela_splitter_573 (
        .a(new_Jinkela_wire_7987),
        .b(new_Jinkela_wire_7988),
        .c(new_Jinkela_wire_7989)
    );

    bfr new_Jinkela_buffer_916 (
        .din(new_Jinkela_wire_986),
        .dout(new_Jinkela_wire_987)
    );

    bfr new_Jinkela_buffer_7355 (
        .din(new_Jinkela_wire_9131),
        .dout(new_Jinkela_wire_9132)
    );

    spl2 new_Jinkela_splitter_33 (
        .a(new_Jinkela_wire_1100),
        .b(new_Jinkela_wire_1101),
        .c(new_Jinkela_wire_1102)
    );

    spl3L new_Jinkela_splitter_723 (
        .a(n_0025_),
        .d(new_Jinkela_wire_9200),
        .b(new_Jinkela_wire_9201),
        .c(new_Jinkela_wire_9202)
    );

    bfr new_Jinkela_buffer_917 (
        .din(new_Jinkela_wire_987),
        .dout(new_Jinkela_wire_988)
    );

    spl2 new_Jinkela_splitter_713 (
        .a(new_Jinkela_wire_9132),
        .b(new_Jinkela_wire_9133),
        .c(new_Jinkela_wire_9134)
    );

    bfr new_Jinkela_buffer_963 (
        .din(new_Jinkela_wire_1037),
        .dout(new_Jinkela_wire_1038)
    );

    bfr new_Jinkela_buffer_918 (
        .din(new_Jinkela_wire_988),
        .dout(new_Jinkela_wire_989)
    );

    bfr new_Jinkela_buffer_7363 (
        .din(new_Jinkela_wire_9161),
        .dout(new_Jinkela_wire_9162)
    );

    spl4L new_Jinkela_splitter_721 (
        .a(n_0037_),
        .d(new_Jinkela_wire_9158),
        .b(new_Jinkela_wire_9159),
        .e(new_Jinkela_wire_9160),
        .c(new_Jinkela_wire_9161)
    );

    bfr new_Jinkela_buffer_1026 (
        .din(new_Jinkela_wire_1102),
        .dout(new_Jinkela_wire_1103)
    );

    bfr new_Jinkela_buffer_919 (
        .din(new_Jinkela_wire_989),
        .dout(new_Jinkela_wire_990)
    );

    spl2 new_Jinkela_splitter_726 (
        .a(n_0675_),
        .b(new_Jinkela_wire_9250),
        .c(new_Jinkela_wire_9251)
    );

    spl4L new_Jinkela_splitter_725 (
        .a(n_0824_),
        .d(new_Jinkela_wire_9246),
        .b(new_Jinkela_wire_9247),
        .e(new_Jinkela_wire_9248),
        .c(new_Jinkela_wire_9249)
    );

    bfr new_Jinkela_buffer_964 (
        .din(new_Jinkela_wire_1038),
        .dout(new_Jinkela_wire_1039)
    );

    spl2 new_Jinkela_splitter_722 (
        .a(new_Jinkela_wire_9162),
        .b(new_Jinkela_wire_9163),
        .c(new_Jinkela_wire_9164)
    );

    bfr new_Jinkela_buffer_920 (
        .din(new_Jinkela_wire_990),
        .dout(new_Jinkela_wire_991)
    );

    bfr new_Jinkela_buffer_7364 (
        .din(new_Jinkela_wire_9164),
        .dout(new_Jinkela_wire_9165)
    );

    bfr new_Jinkela_buffer_1090 (
        .din(new_Jinkela_wire_1396),
        .dout(new_Jinkela_wire_1397)
    );

    bfr new_Jinkela_buffer_921 (
        .din(new_Jinkela_wire_991),
        .dout(new_Jinkela_wire_992)
    );

    bfr new_Jinkela_buffer_7399 (
        .din(new_Jinkela_wire_9202),
        .dout(new_Jinkela_wire_9203)
    );

    spl2 new_Jinkela_splitter_729 (
        .a(n_0232_),
        .b(new_Jinkela_wire_9291),
        .c(new_Jinkela_wire_9292)
    );

    bfr new_Jinkela_buffer_965 (
        .din(new_Jinkela_wire_1039),
        .dout(new_Jinkela_wire_1040)
    );

    bfr new_Jinkela_buffer_7365 (
        .din(new_Jinkela_wire_9165),
        .dout(new_Jinkela_wire_9166)
    );

    bfr new_Jinkela_buffer_922 (
        .din(new_Jinkela_wire_992),
        .dout(new_Jinkela_wire_993)
    );

    bfr new_Jinkela_buffer_7400 (
        .din(new_Jinkela_wire_9203),
        .dout(new_Jinkela_wire_9204)
    );

    bfr new_Jinkela_buffer_1089 (
        .din(new_Jinkela_wire_1395),
        .dout(new_Jinkela_wire_1396)
    );

    bfr new_Jinkela_buffer_1160 (
        .din(N328),
        .dout(new_Jinkela_wire_1472)
    );

    bfr new_Jinkela_buffer_7366 (
        .din(new_Jinkela_wire_9166),
        .dout(new_Jinkela_wire_9167)
    );

    bfr new_Jinkela_buffer_923 (
        .din(new_Jinkela_wire_993),
        .dout(new_Jinkela_wire_994)
    );

    bfr new_Jinkela_buffer_966 (
        .din(new_Jinkela_wire_1040),
        .dout(new_Jinkela_wire_1041)
    );

    spl3L new_Jinkela_splitter_727 (
        .a(n_0061_),
        .d(new_Jinkela_wire_9252),
        .b(new_Jinkela_wire_9253),
        .c(new_Jinkela_wire_9254)
    );

    bfr new_Jinkela_buffer_7367 (
        .din(new_Jinkela_wire_9167),
        .dout(new_Jinkela_wire_9168)
    );

    bfr new_Jinkela_buffer_924 (
        .din(new_Jinkela_wire_994),
        .dout(new_Jinkela_wire_995)
    );

    bfr new_Jinkela_buffer_7401 (
        .din(new_Jinkela_wire_9204),
        .dout(new_Jinkela_wire_9205)
    );

    bfr new_Jinkela_buffer_1027 (
        .din(new_Jinkela_wire_1103),
        .dout(new_Jinkela_wire_1104)
    );

    bfr new_Jinkela_buffer_7368 (
        .din(new_Jinkela_wire_9168),
        .dout(new_Jinkela_wire_9169)
    );

    bfr new_Jinkela_buffer_925 (
        .din(new_Jinkela_wire_995),
        .dout(new_Jinkela_wire_996)
    );

    bfr new_Jinkela_buffer_7440 (
        .din(new_Jinkela_wire_9254),
        .dout(new_Jinkela_wire_9255)
    );

    bfr new_Jinkela_buffer_967 (
        .din(new_Jinkela_wire_1041),
        .dout(new_Jinkela_wire_1042)
    );

    spl2 new_Jinkela_splitter_731 (
        .a(n_0735_),
        .b(new_Jinkela_wire_9298),
        .c(new_Jinkela_wire_9299)
    );

    bfr new_Jinkela_buffer_7369 (
        .din(new_Jinkela_wire_9169),
        .dout(new_Jinkela_wire_9170)
    );

    bfr new_Jinkela_buffer_926 (
        .din(new_Jinkela_wire_996),
        .dout(new_Jinkela_wire_997)
    );

    bfr new_Jinkela_buffer_7402 (
        .din(new_Jinkela_wire_9205),
        .dout(new_Jinkela_wire_9206)
    );

    bfr new_Jinkela_buffer_1096 (
        .din(N280),
        .dout(new_Jinkela_wire_1403)
    );

    bfr new_Jinkela_buffer_7370 (
        .din(new_Jinkela_wire_9170),
        .dout(new_Jinkela_wire_9171)
    );

    bfr new_Jinkela_buffer_927 (
        .din(new_Jinkela_wire_997),
        .dout(new_Jinkela_wire_998)
    );

    spl2 new_Jinkela_splitter_730 (
        .a(n_0950_),
        .b(new_Jinkela_wire_9296),
        .c(new_Jinkela_wire_9297)
    );

    bfr new_Jinkela_buffer_968 (
        .din(new_Jinkela_wire_1042),
        .dout(new_Jinkela_wire_1043)
    );

    bfr new_Jinkela_buffer_7371 (
        .din(new_Jinkela_wire_9171),
        .dout(new_Jinkela_wire_9172)
    );

    bfr new_Jinkela_buffer_928 (
        .din(new_Jinkela_wire_998),
        .dout(new_Jinkela_wire_999)
    );

    bfr new_Jinkela_buffer_7403 (
        .din(new_Jinkela_wire_9206),
        .dout(new_Jinkela_wire_9207)
    );

    bfr new_Jinkela_buffer_1093 (
        .din(new_Jinkela_wire_1399),
        .dout(new_Jinkela_wire_1400)
    );

    bfr new_Jinkela_buffer_1028 (
        .din(new_Jinkela_wire_1104),
        .dout(new_Jinkela_wire_1105)
    );

    bfr new_Jinkela_buffer_7372 (
        .din(new_Jinkela_wire_9172),
        .dout(new_Jinkela_wire_9173)
    );

    bfr new_Jinkela_buffer_929 (
        .din(new_Jinkela_wire_999),
        .dout(new_Jinkela_wire_1000)
    );

    bfr new_Jinkela_buffer_7474 (
        .din(new_Jinkela_wire_9292),
        .dout(new_Jinkela_wire_9293)
    );

    bfr new_Jinkela_buffer_969 (
        .din(new_Jinkela_wire_1043),
        .dout(new_Jinkela_wire_1044)
    );

    bfr new_Jinkela_buffer_7373 (
        .din(new_Jinkela_wire_9173),
        .dout(new_Jinkela_wire_9174)
    );

    bfr new_Jinkela_buffer_930 (
        .din(new_Jinkela_wire_1000),
        .dout(new_Jinkela_wire_1001)
    );

    bfr new_Jinkela_buffer_7404 (
        .din(new_Jinkela_wire_9207),
        .dout(new_Jinkela_wire_9208)
    );

    bfr new_Jinkela_buffer_7374 (
        .din(new_Jinkela_wire_9174),
        .dout(new_Jinkela_wire_9175)
    );

    bfr new_Jinkela_buffer_931 (
        .din(new_Jinkela_wire_1001),
        .dout(new_Jinkela_wire_1002)
    );

    bfr new_Jinkela_buffer_7441 (
        .din(new_Jinkela_wire_9255),
        .dout(new_Jinkela_wire_9256)
    );

    bfr new_Jinkela_buffer_970 (
        .din(new_Jinkela_wire_1044),
        .dout(new_Jinkela_wire_1045)
    );

    bfr new_Jinkela_buffer_7375 (
        .din(new_Jinkela_wire_9175),
        .dout(new_Jinkela_wire_9176)
    );

    bfr new_Jinkela_buffer_932 (
        .din(new_Jinkela_wire_1002),
        .dout(new_Jinkela_wire_1003)
    );

    bfr new_Jinkela_buffer_7405 (
        .din(new_Jinkela_wire_9208),
        .dout(new_Jinkela_wire_9209)
    );

    bfr new_Jinkela_buffer_1029 (
        .din(new_Jinkela_wire_1105),
        .dout(new_Jinkela_wire_1106)
    );

    bfr new_Jinkela_buffer_7376 (
        .din(new_Jinkela_wire_9176),
        .dout(new_Jinkela_wire_9177)
    );

    bfr new_Jinkela_buffer_933 (
        .din(new_Jinkela_wire_1003),
        .dout(new_Jinkela_wire_1004)
    );

    bfr new_Jinkela_buffer_971 (
        .din(new_Jinkela_wire_1045),
        .dout(new_Jinkela_wire_1046)
    );

    bfr new_Jinkela_buffer_7377 (
        .din(new_Jinkela_wire_9177),
        .dout(new_Jinkela_wire_9178)
    );

    bfr new_Jinkela_buffer_934 (
        .din(new_Jinkela_wire_1004),
        .dout(new_Jinkela_wire_1005)
    );

    bfr new_Jinkela_buffer_7406 (
        .din(new_Jinkela_wire_9209),
        .dout(new_Jinkela_wire_9210)
    );

    bfr new_Jinkela_buffer_1092 (
        .din(N141),
        .dout(new_Jinkela_wire_1399)
    );

    bfr new_Jinkela_buffer_7378 (
        .din(new_Jinkela_wire_9178),
        .dout(new_Jinkela_wire_9179)
    );

    bfr new_Jinkela_buffer_935 (
        .din(new_Jinkela_wire_1005),
        .dout(new_Jinkela_wire_1006)
    );

    bfr new_Jinkela_buffer_7442 (
        .din(new_Jinkela_wire_9256),
        .dout(new_Jinkela_wire_9257)
    );

    bfr new_Jinkela_buffer_972 (
        .din(new_Jinkela_wire_1046),
        .dout(new_Jinkela_wire_1047)
    );

    bfr new_Jinkela_buffer_7379 (
        .din(new_Jinkela_wire_9179),
        .dout(new_Jinkela_wire_9180)
    );

    bfr new_Jinkela_buffer_936 (
        .din(new_Jinkela_wire_1006),
        .dout(new_Jinkela_wire_1007)
    );

    bfr new_Jinkela_buffer_7407 (
        .din(new_Jinkela_wire_9210),
        .dout(new_Jinkela_wire_9211)
    );

    bfr new_Jinkela_buffer_1091 (
        .din(new_Jinkela_wire_1397),
        .dout(new_Jinkela_wire_1398)
    );

    bfr new_Jinkela_buffer_1030 (
        .din(new_Jinkela_wire_1106),
        .dout(new_Jinkela_wire_1107)
    );

    bfr new_Jinkela_buffer_7380 (
        .din(new_Jinkela_wire_9180),
        .dout(new_Jinkela_wire_9181)
    );

    bfr new_Jinkela_buffer_7358 (
        .din(new_Jinkela_wire_9143),
        .dout(new_Jinkela_wire_9144)
    );

    bfr new_Jinkela_buffer_7314 (
        .din(new_Jinkela_wire_9077),
        .dout(new_Jinkela_wire_9078)
    );

    bfr new_Jinkela_buffer_4831 (
        .din(new_Jinkela_wire_5765),
        .dout(new_Jinkela_wire_5766)
    );

    bfr new_Jinkela_buffer_4819 (
        .din(new_Jinkela_wire_5750),
        .dout(new_Jinkela_wire_5751)
    );

    bfr new_Jinkela_buffer_7475 (
        .din(new_Jinkela_wire_9293),
        .dout(new_Jinkela_wire_9294)
    );

    bfr new_Jinkela_buffer_4791 (
        .din(new_Jinkela_wire_5718),
        .dout(new_Jinkela_wire_5719)
    );

    bfr new_Jinkela_buffer_7381 (
        .din(new_Jinkela_wire_9181),
        .dout(new_Jinkela_wire_9182)
    );

    bfr new_Jinkela_buffer_7408 (
        .din(new_Jinkela_wire_9211),
        .dout(new_Jinkela_wire_9212)
    );

    bfr new_Jinkela_buffer_4792 (
        .din(new_Jinkela_wire_5719),
        .dout(new_Jinkela_wire_5720)
    );

    bfr new_Jinkela_buffer_7382 (
        .din(new_Jinkela_wire_9182),
        .dout(new_Jinkela_wire_9183)
    );

    spl2 new_Jinkela_splitter_361 (
        .a(n_0099_),
        .b(new_Jinkela_wire_5883),
        .c(new_Jinkela_wire_5884)
    );

    bfr new_Jinkela_buffer_4820 (
        .din(new_Jinkela_wire_5751),
        .dout(new_Jinkela_wire_5752)
    );

    bfr new_Jinkela_buffer_7443 (
        .din(new_Jinkela_wire_9257),
        .dout(new_Jinkela_wire_9258)
    );

    bfr new_Jinkela_buffer_4793 (
        .din(new_Jinkela_wire_5720),
        .dout(new_Jinkela_wire_5721)
    );

    bfr new_Jinkela_buffer_7383 (
        .din(new_Jinkela_wire_9183),
        .dout(new_Jinkela_wire_9184)
    );

    bfr new_Jinkela_buffer_4873 (
        .din(new_Jinkela_wire_5809),
        .dout(new_Jinkela_wire_5810)
    );

    bfr new_Jinkela_buffer_7409 (
        .din(new_Jinkela_wire_9212),
        .dout(new_Jinkela_wire_9213)
    );

    bfr new_Jinkela_buffer_4794 (
        .din(new_Jinkela_wire_5721),
        .dout(new_Jinkela_wire_5722)
    );

    bfr new_Jinkela_buffer_7384 (
        .din(new_Jinkela_wire_9184),
        .dout(new_Jinkela_wire_9185)
    );

    bfr new_Jinkela_buffer_4832 (
        .din(new_Jinkela_wire_5766),
        .dout(new_Jinkela_wire_5767)
    );

    bfr new_Jinkela_buffer_4821 (
        .din(new_Jinkela_wire_5752),
        .dout(new_Jinkela_wire_5753)
    );

    spl2 new_Jinkela_splitter_732 (
        .a(n_0884_),
        .b(new_Jinkela_wire_9300),
        .c(new_Jinkela_wire_9301)
    );

    bfr new_Jinkela_buffer_4795 (
        .din(new_Jinkela_wire_5722),
        .dout(new_Jinkela_wire_5723)
    );

    bfr new_Jinkela_buffer_7385 (
        .din(new_Jinkela_wire_9185),
        .dout(new_Jinkela_wire_9186)
    );

    bfr new_Jinkela_buffer_7410 (
        .din(new_Jinkela_wire_9213),
        .dout(new_Jinkela_wire_9214)
    );

    bfr new_Jinkela_buffer_4796 (
        .din(new_Jinkela_wire_5723),
        .dout(new_Jinkela_wire_5724)
    );

    bfr new_Jinkela_buffer_7386 (
        .din(new_Jinkela_wire_9186),
        .dout(new_Jinkela_wire_9187)
    );

    bfr new_Jinkela_buffer_7350 (
        .din(new_Jinkela_wire_9126),
        .dout(new_Jinkela_wire_9127)
    );

    bfr new_Jinkela_buffer_4822 (
        .din(new_Jinkela_wire_5753),
        .dout(new_Jinkela_wire_5754)
    );

    bfr new_Jinkela_buffer_7444 (
        .din(new_Jinkela_wire_9258),
        .dout(new_Jinkela_wire_9259)
    );

    bfr new_Jinkela_buffer_4797 (
        .din(new_Jinkela_wire_5724),
        .dout(new_Jinkela_wire_5725)
    );

    bfr new_Jinkela_buffer_7387 (
        .din(new_Jinkela_wire_9187),
        .dout(new_Jinkela_wire_9188)
    );

    bfr new_Jinkela_buffer_7411 (
        .din(new_Jinkela_wire_9214),
        .dout(new_Jinkela_wire_9215)
    );

    bfr new_Jinkela_buffer_4798 (
        .din(new_Jinkela_wire_5725),
        .dout(new_Jinkela_wire_5726)
    );

    bfr new_Jinkela_buffer_7388 (
        .din(new_Jinkela_wire_9188),
        .dout(new_Jinkela_wire_9189)
    );

    bfr new_Jinkela_buffer_4833 (
        .din(new_Jinkela_wire_5767),
        .dout(new_Jinkela_wire_5768)
    );

    bfr new_Jinkela_buffer_7476 (
        .din(new_Jinkela_wire_9294),
        .dout(new_Jinkela_wire_9295)
    );

    bfr new_Jinkela_buffer_4799 (
        .din(new_Jinkela_wire_5726),
        .dout(new_Jinkela_wire_5727)
    );

    bfr new_Jinkela_buffer_7389 (
        .din(new_Jinkela_wire_9189),
        .dout(new_Jinkela_wire_9190)
    );

    bfr new_Jinkela_buffer_4874 (
        .din(new_Jinkela_wire_5810),
        .dout(new_Jinkela_wire_5811)
    );

    bfr new_Jinkela_buffer_7412 (
        .din(new_Jinkela_wire_9215),
        .dout(new_Jinkela_wire_9216)
    );

    spl2 new_Jinkela_splitter_353 (
        .a(new_Jinkela_wire_5727),
        .b(new_Jinkela_wire_5728),
        .c(new_Jinkela_wire_5729)
    );

    bfr new_Jinkela_buffer_7390 (
        .din(new_Jinkela_wire_9190),
        .dout(new_Jinkela_wire_9191)
    );

    bfr new_Jinkela_buffer_4943 (
        .din(new_net_2574),
        .dout(new_Jinkela_wire_5893)
    );

    bfr new_Jinkela_buffer_7445 (
        .din(new_Jinkela_wire_9259),
        .dout(new_Jinkela_wire_9260)
    );

    bfr new_Jinkela_buffer_4834 (
        .din(new_Jinkela_wire_5768),
        .dout(new_Jinkela_wire_5769)
    );

    bfr new_Jinkela_buffer_7391 (
        .din(new_Jinkela_wire_9191),
        .dout(new_Jinkela_wire_9192)
    );

    bfr new_Jinkela_buffer_4835 (
        .din(new_Jinkela_wire_5769),
        .dout(new_Jinkela_wire_5770)
    );

    bfr new_Jinkela_buffer_7413 (
        .din(new_Jinkela_wire_9216),
        .dout(new_Jinkela_wire_9217)
    );

    bfr new_Jinkela_buffer_4935 (
        .din(new_Jinkela_wire_5884),
        .dout(new_Jinkela_wire_5885)
    );

    bfr new_Jinkela_buffer_4875 (
        .din(new_Jinkela_wire_5811),
        .dout(new_Jinkela_wire_5812)
    );

    bfr new_Jinkela_buffer_7392 (
        .din(new_Jinkela_wire_9192),
        .dout(new_Jinkela_wire_9193)
    );

    bfr new_Jinkela_buffer_4836 (
        .din(new_Jinkela_wire_5770),
        .dout(new_Jinkela_wire_5771)
    );

    bfr new_Jinkela_buffer_7393 (
        .din(new_Jinkela_wire_9193),
        .dout(new_Jinkela_wire_9194)
    );

    bfr new_Jinkela_buffer_4837 (
        .din(new_Jinkela_wire_5771),
        .dout(new_Jinkela_wire_5772)
    );

    bfr new_Jinkela_buffer_7414 (
        .din(new_Jinkela_wire_9217),
        .dout(new_Jinkela_wire_9218)
    );

    bfr new_Jinkela_buffer_4876 (
        .din(new_Jinkela_wire_5812),
        .dout(new_Jinkela_wire_5813)
    );

    bfr new_Jinkela_buffer_7394 (
        .din(new_Jinkela_wire_9194),
        .dout(new_Jinkela_wire_9195)
    );

    bfr new_Jinkela_buffer_4838 (
        .din(new_Jinkela_wire_5772),
        .dout(new_Jinkela_wire_5773)
    );

    bfr new_Jinkela_buffer_7446 (
        .din(new_Jinkela_wire_9260),
        .dout(new_Jinkela_wire_9261)
    );

    bfr new_Jinkela_buffer_7395 (
        .din(new_Jinkela_wire_9195),
        .dout(new_Jinkela_wire_9196)
    );

    bfr new_Jinkela_buffer_4839 (
        .din(new_Jinkela_wire_5773),
        .dout(new_Jinkela_wire_5774)
    );

    bfr new_Jinkela_buffer_7415 (
        .din(new_Jinkela_wire_9218),
        .dout(new_Jinkela_wire_9219)
    );

    spl2 new_Jinkela_splitter_362 (
        .a(n_1333_),
        .b(new_Jinkela_wire_5918),
        .c(new_Jinkela_wire_5919)
    );

    bfr new_Jinkela_buffer_4877 (
        .din(new_Jinkela_wire_5813),
        .dout(new_Jinkela_wire_5814)
    );

    bfr new_Jinkela_buffer_7396 (
        .din(new_Jinkela_wire_9196),
        .dout(new_Jinkela_wire_9197)
    );

    bfr new_Jinkela_buffer_4840 (
        .din(new_Jinkela_wire_5774),
        .dout(new_Jinkela_wire_5775)
    );

    spl2 new_Jinkela_splitter_733 (
        .a(n_0830_),
        .b(new_Jinkela_wire_9302),
        .c(new_Jinkela_wire_9303)
    );

    spl3L new_Jinkela_splitter_736 (
        .a(n_1295_),
        .d(new_Jinkela_wire_9341),
        .b(new_Jinkela_wire_9342),
        .c(new_Jinkela_wire_9343)
    );

    bfr new_Jinkela_buffer_4973 (
        .din(n_0671_),
        .dout(new_Jinkela_wire_5927)
    );

    bfr new_Jinkela_buffer_7397 (
        .din(new_Jinkela_wire_9197),
        .dout(new_Jinkela_wire_9198)
    );

    bfr new_Jinkela_buffer_4841 (
        .din(new_Jinkela_wire_5775),
        .dout(new_Jinkela_wire_5776)
    );

    bfr new_Jinkela_buffer_7416 (
        .din(new_Jinkela_wire_9219),
        .dout(new_Jinkela_wire_9220)
    );

    bfr new_Jinkela_buffer_4944 (
        .din(new_Jinkela_wire_5893),
        .dout(new_Jinkela_wire_5894)
    );

    bfr new_Jinkela_buffer_4878 (
        .din(new_Jinkela_wire_5814),
        .dout(new_Jinkela_wire_5815)
    );

    bfr new_Jinkela_buffer_7398 (
        .din(new_Jinkela_wire_9198),
        .dout(new_Jinkela_wire_9199)
    );

    bfr new_Jinkela_buffer_4842 (
        .din(new_Jinkela_wire_5776),
        .dout(new_Jinkela_wire_5777)
    );

    bfr new_Jinkela_buffer_7447 (
        .din(new_Jinkela_wire_9261),
        .dout(new_Jinkela_wire_9262)
    );

    bfr new_Jinkela_buffer_4936 (
        .din(new_Jinkela_wire_5885),
        .dout(new_Jinkela_wire_5886)
    );

    bfr new_Jinkela_buffer_7417 (
        .din(new_Jinkela_wire_9220),
        .dout(new_Jinkela_wire_9221)
    );

    bfr new_Jinkela_buffer_4843 (
        .din(new_Jinkela_wire_5777),
        .dout(new_Jinkela_wire_5778)
    );

    bfr new_Jinkela_buffer_7477 (
        .din(new_net_2525),
        .dout(new_Jinkela_wire_9304)
    );

    spl2 new_Jinkela_splitter_734 (
        .a(n_0078_),
        .b(new_Jinkela_wire_9336),
        .c(new_Jinkela_wire_9337)
    );

    bfr new_Jinkela_buffer_4879 (
        .din(new_Jinkela_wire_5815),
        .dout(new_Jinkela_wire_5816)
    );

    bfr new_Jinkela_buffer_7418 (
        .din(new_Jinkela_wire_9221),
        .dout(new_Jinkela_wire_9222)
    );

    bfr new_Jinkela_buffer_4844 (
        .din(new_Jinkela_wire_5778),
        .dout(new_Jinkela_wire_5779)
    );

    bfr new_Jinkela_buffer_7448 (
        .din(new_Jinkela_wire_9262),
        .dout(new_Jinkela_wire_9263)
    );

    bfr new_Jinkela_buffer_7419 (
        .din(new_Jinkela_wire_9222),
        .dout(new_Jinkela_wire_9223)
    );

    bfr new_Jinkela_buffer_2281 (
        .din(new_Jinkela_wire_2669),
        .dout(new_Jinkela_wire_2670)
    );

    bfr new_Jinkela_buffer_5661 (
        .din(new_Jinkela_wire_6808),
        .dout(new_Jinkela_wire_6809)
    );

    spl2 new_Jinkela_splitter_446 (
        .a(n_0280_),
        .b(new_Jinkela_wire_6815),
        .c(new_Jinkela_wire_6816)
    );

    bfr new_Jinkela_buffer_2223 (
        .din(new_Jinkela_wire_2609),
        .dout(new_Jinkela_wire_2610)
    );

    spl3L new_Jinkela_splitter_447 (
        .a(n_0038_),
        .d(new_Jinkela_wire_6822),
        .b(new_Jinkela_wire_6823),
        .c(new_Jinkela_wire_6824)
    );

    bfr new_Jinkela_buffer_2416 (
        .din(N177),
        .dout(new_Jinkela_wire_2813)
    );

    bfr new_Jinkela_buffer_5667 (
        .din(new_Jinkela_wire_6816),
        .dout(new_Jinkela_wire_6817)
    );

    bfr new_Jinkela_buffer_2224 (
        .din(new_Jinkela_wire_2610),
        .dout(new_Jinkela_wire_2611)
    );

    bfr new_Jinkela_buffer_5662 (
        .din(new_Jinkela_wire_6809),
        .dout(new_Jinkela_wire_6810)
    );

    spl3L new_Jinkela_splitter_130 (
        .a(new_Jinkela_wire_2670),
        .d(new_Jinkela_wire_2671),
        .b(new_Jinkela_wire_2672),
        .c(new_Jinkela_wire_2673)
    );

    bfr new_Jinkela_buffer_2225 (
        .din(new_Jinkela_wire_2611),
        .dout(new_Jinkela_wire_2612)
    );

    bfr new_Jinkela_buffer_5663 (
        .din(new_Jinkela_wire_6810),
        .dout(new_Jinkela_wire_6811)
    );

    bfr new_Jinkela_buffer_2346 (
        .din(new_Jinkela_wire_2737),
        .dout(new_Jinkela_wire_2738)
    );

    bfr new_Jinkela_buffer_2409 (
        .din(new_Jinkela_wire_2805),
        .dout(new_Jinkela_wire_2806)
    );

    spl2 new_Jinkela_splitter_448 (
        .a(n_0684_),
        .b(new_Jinkela_wire_6825),
        .c(new_Jinkela_wire_6826)
    );

    bfr new_Jinkela_buffer_2226 (
        .din(new_Jinkela_wire_2612),
        .dout(new_Jinkela_wire_2613)
    );

    bfr new_Jinkela_buffer_5664 (
        .din(new_Jinkela_wire_6811),
        .dout(new_Jinkela_wire_6812)
    );

    bfr new_Jinkela_buffer_2282 (
        .din(new_Jinkela_wire_2673),
        .dout(new_Jinkela_wire_2674)
    );

    bfr new_Jinkela_buffer_5675 (
        .din(n_1122_),
        .dout(new_Jinkela_wire_6830)
    );

    bfr new_Jinkela_buffer_2227 (
        .din(new_Jinkela_wire_2613),
        .dout(new_Jinkela_wire_2614)
    );

    bfr new_Jinkela_buffer_5665 (
        .din(new_Jinkela_wire_6812),
        .dout(new_Jinkela_wire_6813)
    );

    bfr new_Jinkela_buffer_2345 (
        .din(new_Jinkela_wire_2736),
        .dout(new_Jinkela_wire_2737)
    );

    bfr new_Jinkela_buffer_5668 (
        .din(new_Jinkela_wire_6817),
        .dout(new_Jinkela_wire_6818)
    );

    bfr new_Jinkela_buffer_2228 (
        .din(new_Jinkela_wire_2614),
        .dout(new_Jinkela_wire_2615)
    );

    bfr new_Jinkela_buffer_5672 (
        .din(new_Jinkela_wire_6826),
        .dout(new_Jinkela_wire_6827)
    );

    bfr new_Jinkela_buffer_2283 (
        .din(new_Jinkela_wire_2674),
        .dout(new_Jinkela_wire_2675)
    );

    bfr new_Jinkela_buffer_5669 (
        .din(new_Jinkela_wire_6818),
        .dout(new_Jinkela_wire_6819)
    );

    bfr new_Jinkela_buffer_2229 (
        .din(new_Jinkela_wire_2615),
        .dout(new_Jinkela_wire_2616)
    );

    bfr new_Jinkela_buffer_5677 (
        .din(n_1193_),
        .dout(new_Jinkela_wire_6834)
    );

    spl2 new_Jinkela_splitter_131 (
        .a(new_Jinkela_wire_2738),
        .b(new_Jinkela_wire_2739),
        .c(new_Jinkela_wire_2740)
    );

    bfr new_Jinkela_buffer_5670 (
        .din(new_Jinkela_wire_6819),
        .dout(new_Jinkela_wire_6820)
    );

    bfr new_Jinkela_buffer_2230 (
        .din(new_Jinkela_wire_2616),
        .dout(new_Jinkela_wire_2617)
    );

    spl4L new_Jinkela_splitter_451 (
        .a(n_0827_),
        .d(new_Jinkela_wire_6839),
        .b(new_Jinkela_wire_6840),
        .e(new_Jinkela_wire_6841),
        .c(new_Jinkela_wire_6842)
    );

    bfr new_Jinkela_buffer_2284 (
        .din(new_Jinkela_wire_2675),
        .dout(new_Jinkela_wire_2676)
    );

    bfr new_Jinkela_buffer_5671 (
        .din(new_Jinkela_wire_6820),
        .dout(new_Jinkela_wire_6821)
    );

    bfr new_Jinkela_buffer_2231 (
        .din(new_Jinkela_wire_2617),
        .dout(new_Jinkela_wire_2618)
    );

    bfr new_Jinkela_buffer_5673 (
        .din(new_Jinkela_wire_6827),
        .dout(new_Jinkela_wire_6828)
    );

    bfr new_Jinkela_buffer_2347 (
        .din(new_Jinkela_wire_2740),
        .dout(new_Jinkela_wire_2741)
    );

    bfr new_Jinkela_buffer_5676 (
        .din(new_Jinkela_wire_6830),
        .dout(new_Jinkela_wire_6831)
    );

    bfr new_Jinkela_buffer_2232 (
        .din(new_Jinkela_wire_2618),
        .dout(new_Jinkela_wire_2619)
    );

    bfr new_Jinkela_buffer_5674 (
        .din(new_Jinkela_wire_6828),
        .dout(new_Jinkela_wire_6829)
    );

    bfr new_Jinkela_buffer_2285 (
        .din(new_Jinkela_wire_2676),
        .dout(new_Jinkela_wire_2677)
    );

    bfr new_Jinkela_buffer_5716 (
        .din(new_Jinkela_wire_6888),
        .dout(new_Jinkela_wire_6889)
    );

    bfr new_Jinkela_buffer_2233 (
        .din(new_Jinkela_wire_2619),
        .dout(new_Jinkela_wire_2620)
    );

    spl2 new_Jinkela_splitter_449 (
        .a(new_Jinkela_wire_6831),
        .b(new_Jinkela_wire_6832),
        .c(new_Jinkela_wire_6833)
    );

    bfr new_Jinkela_buffer_5718 (
        .din(new_Jinkela_wire_6892),
        .dout(new_Jinkela_wire_6893)
    );

    spl3L new_Jinkela_splitter_452 (
        .a(n_0360_),
        .d(new_Jinkela_wire_6843),
        .b(new_Jinkela_wire_6844),
        .c(new_Jinkela_wire_6845)
    );

    bfr new_Jinkela_buffer_2234 (
        .din(new_Jinkela_wire_2620),
        .dout(new_Jinkela_wire_2621)
    );

    bfr new_Jinkela_buffer_5678 (
        .din(new_Jinkela_wire_6834),
        .dout(new_Jinkela_wire_6835)
    );

    bfr new_Jinkela_buffer_2286 (
        .din(new_Jinkela_wire_2677),
        .dout(new_Jinkela_wire_2678)
    );

    bfr new_Jinkela_buffer_5679 (
        .din(new_Jinkela_wire_6835),
        .dout(new_Jinkela_wire_6836)
    );

    bfr new_Jinkela_buffer_2235 (
        .din(new_Jinkela_wire_2621),
        .dout(new_Jinkela_wire_2622)
    );

    bfr new_Jinkela_buffer_5720 (
        .din(n_1341_),
        .dout(new_Jinkela_wire_6895)
    );

    bfr new_Jinkela_buffer_2410 (
        .din(new_Jinkela_wire_2806),
        .dout(new_Jinkela_wire_2807)
    );

    spl2 new_Jinkela_splitter_450 (
        .a(new_Jinkela_wire_6836),
        .b(new_Jinkela_wire_6837),
        .c(new_Jinkela_wire_6838)
    );

    bfr new_Jinkela_buffer_2236 (
        .din(new_Jinkela_wire_2622),
        .dout(new_Jinkela_wire_2623)
    );

    spl2 new_Jinkela_splitter_456 (
        .a(n_1123_),
        .b(new_Jinkela_wire_6891),
        .c(new_Jinkela_wire_6892)
    );

    bfr new_Jinkela_buffer_2287 (
        .din(new_Jinkela_wire_2678),
        .dout(new_Jinkela_wire_2679)
    );

    spl2 new_Jinkela_splitter_455 (
        .a(n_1133_),
        .b(new_Jinkela_wire_6887),
        .c(new_Jinkela_wire_6888)
    );

    bfr new_Jinkela_buffer_2237 (
        .din(new_Jinkela_wire_2623),
        .dout(new_Jinkela_wire_2624)
    );

    bfr new_Jinkela_buffer_5681 (
        .din(new_Jinkela_wire_6846),
        .dout(new_Jinkela_wire_6847)
    );

    bfr new_Jinkela_buffer_2413 (
        .din(new_Jinkela_wire_2809),
        .dout(new_Jinkela_wire_2810)
    );

    bfr new_Jinkela_buffer_5680 (
        .din(new_Jinkela_wire_6845),
        .dout(new_Jinkela_wire_6846)
    );

    bfr new_Jinkela_buffer_5682 (
        .din(new_Jinkela_wire_6847),
        .dout(new_Jinkela_wire_6848)
    );

    bfr new_Jinkela_buffer_2238 (
        .din(new_Jinkela_wire_2624),
        .dout(new_Jinkela_wire_2625)
    );

    bfr new_Jinkela_buffer_2288 (
        .din(new_Jinkela_wire_2679),
        .dout(new_Jinkela_wire_2680)
    );

    bfr new_Jinkela_buffer_2239 (
        .din(new_Jinkela_wire_2625),
        .dout(new_Jinkela_wire_2626)
    );

    bfr new_Jinkela_buffer_5717 (
        .din(new_Jinkela_wire_6889),
        .dout(new_Jinkela_wire_6890)
    );

    bfr new_Jinkela_buffer_2348 (
        .din(new_Jinkela_wire_2741),
        .dout(new_Jinkela_wire_2742)
    );

    spl3L new_Jinkela_splitter_453 (
        .a(new_Jinkela_wire_6848),
        .d(new_Jinkela_wire_6849),
        .b(new_Jinkela_wire_6850),
        .c(new_Jinkela_wire_6851)
    );

    bfr new_Jinkela_buffer_2240 (
        .din(new_Jinkela_wire_2626),
        .dout(new_Jinkela_wire_2627)
    );

    bfr new_Jinkela_buffer_5725 (
        .din(n_0289_),
        .dout(new_Jinkela_wire_6902)
    );

    bfr new_Jinkela_buffer_2289 (
        .din(new_Jinkela_wire_2680),
        .dout(new_Jinkela_wire_2681)
    );

    bfr new_Jinkela_buffer_5683 (
        .din(new_Jinkela_wire_6851),
        .dout(new_Jinkela_wire_6852)
    );

    bfr new_Jinkela_buffer_2241 (
        .din(new_Jinkela_wire_2627),
        .dout(new_Jinkela_wire_2628)
    );

    bfr new_Jinkela_buffer_5726 (
        .din(n_0153_),
        .dout(new_Jinkela_wire_6903)
    );

    bfr new_Jinkela_buffer_2411 (
        .din(new_Jinkela_wire_2807),
        .dout(new_Jinkela_wire_2808)
    );

    bfr new_Jinkela_buffer_5684 (
        .din(new_Jinkela_wire_6852),
        .dout(new_Jinkela_wire_6853)
    );

    bfr new_Jinkela_buffer_2242 (
        .din(new_Jinkela_wire_2628),
        .dout(new_Jinkela_wire_2629)
    );

    bfr new_Jinkela_buffer_5719 (
        .din(new_Jinkela_wire_6893),
        .dout(new_Jinkela_wire_6894)
    );

    bfr new_Jinkela_buffer_2290 (
        .din(new_Jinkela_wire_2681),
        .dout(new_Jinkela_wire_2682)
    );

    bfr new_Jinkela_buffer_5685 (
        .din(new_Jinkela_wire_6853),
        .dout(new_Jinkela_wire_6854)
    );

    bfr new_Jinkela_buffer_2243 (
        .din(new_Jinkela_wire_2629),
        .dout(new_Jinkela_wire_2630)
    );

    bfr new_Jinkela_buffer_5721 (
        .din(new_Jinkela_wire_6895),
        .dout(new_Jinkela_wire_6896)
    );

    bfr new_Jinkela_buffer_937 (
        .din(new_Jinkela_wire_1007),
        .dout(new_Jinkela_wire_1008)
    );

    spl2 new_Jinkela_splitter_156 (
        .a(n_0342_),
        .b(new_Jinkela_wire_3675),
        .c(new_Jinkela_wire_3676)
    );

    bfr new_Jinkela_buffer_6514 (
        .din(new_Jinkela_wire_7961),
        .dout(new_Jinkela_wire_7962)
    );

    bfr new_Jinkela_buffer_3134 (
        .din(new_Jinkela_wire_3572),
        .dout(new_Jinkela_wire_3573)
    );

    bfr new_Jinkela_buffer_6467 (
        .din(new_Jinkela_wire_7893),
        .dout(new_Jinkela_wire_7894)
    );

    bfr new_Jinkela_buffer_973 (
        .din(new_Jinkela_wire_1047),
        .dout(new_Jinkela_wire_1048)
    );

    bfr new_Jinkela_buffer_3143 (
        .din(new_Jinkela_wire_3595),
        .dout(new_Jinkela_wire_3596)
    );

    bfr new_Jinkela_buffer_938 (
        .din(new_Jinkela_wire_1008),
        .dout(new_Jinkela_wire_1009)
    );

    bfr new_Jinkela_buffer_3142 (
        .din(new_Jinkela_wire_3591),
        .dout(new_Jinkela_wire_3592)
    );

    bfr new_Jinkela_buffer_3135 (
        .din(new_Jinkela_wire_3573),
        .dout(new_Jinkela_wire_3574)
    );

    bfr new_Jinkela_buffer_6468 (
        .din(new_Jinkela_wire_7894),
        .dout(new_Jinkela_wire_7895)
    );

    spl3L new_Jinkela_splitter_577 (
        .a(n_1012_),
        .d(new_Jinkela_wire_7998),
        .b(new_Jinkela_wire_7999),
        .c(new_Jinkela_wire_8000)
    );

    bfr new_Jinkela_buffer_939 (
        .din(new_Jinkela_wire_1009),
        .dout(new_Jinkela_wire_1010)
    );

    bfr new_Jinkela_buffer_3157 (
        .din(new_Jinkela_wire_3611),
        .dout(new_Jinkela_wire_3612)
    );

    bfr new_Jinkela_buffer_6515 (
        .din(new_Jinkela_wire_7962),
        .dout(new_Jinkela_wire_7963)
    );

    bfr new_Jinkela_buffer_3136 (
        .din(new_Jinkela_wire_3574),
        .dout(new_Jinkela_wire_3575)
    );

    bfr new_Jinkela_buffer_6469 (
        .din(new_Jinkela_wire_7895),
        .dout(new_Jinkela_wire_7896)
    );

    bfr new_Jinkela_buffer_974 (
        .din(new_Jinkela_wire_1048),
        .dout(new_Jinkela_wire_1049)
    );

    bfr new_Jinkela_buffer_940 (
        .din(new_Jinkela_wire_1010),
        .dout(new_Jinkela_wire_1011)
    );

    bfr new_Jinkela_buffer_6546 (
        .din(n_0379_),
        .dout(new_Jinkela_wire_8010)
    );

    bfr new_Jinkela_buffer_3137 (
        .din(new_Jinkela_wire_3575),
        .dout(new_Jinkela_wire_3576)
    );

    bfr new_Jinkela_buffer_6470 (
        .din(new_Jinkela_wire_7896),
        .dout(new_Jinkela_wire_7897)
    );

    bfr new_Jinkela_buffer_1094 (
        .din(new_Jinkela_wire_1400),
        .dout(new_Jinkela_wire_1401)
    );

    bfr new_Jinkela_buffer_1031 (
        .din(new_Jinkela_wire_1107),
        .dout(new_Jinkela_wire_1108)
    );

    bfr new_Jinkela_buffer_941 (
        .din(new_Jinkela_wire_1011),
        .dout(new_Jinkela_wire_1012)
    );

    bfr new_Jinkela_buffer_6516 (
        .din(new_Jinkela_wire_7963),
        .dout(new_Jinkela_wire_7964)
    );

    bfr new_Jinkela_buffer_3144 (
        .din(new_Jinkela_wire_3596),
        .dout(new_Jinkela_wire_3597)
    );

    bfr new_Jinkela_buffer_6471 (
        .din(new_Jinkela_wire_7897),
        .dout(new_Jinkela_wire_7898)
    );

    bfr new_Jinkela_buffer_975 (
        .din(new_Jinkela_wire_1049),
        .dout(new_Jinkela_wire_1050)
    );

    spl2 new_Jinkela_splitter_157 (
        .a(n_1336_),
        .b(new_Jinkela_wire_3677),
        .c(new_Jinkela_wire_3678)
    );

    bfr new_Jinkela_buffer_942 (
        .din(new_Jinkela_wire_1012),
        .dout(new_Jinkela_wire_1013)
    );

    bfr new_Jinkela_buffer_6541 (
        .din(n_1297_),
        .dout(new_Jinkela_wire_8003)
    );

    bfr new_Jinkela_buffer_3145 (
        .din(new_Jinkela_wire_3597),
        .dout(new_Jinkela_wire_3598)
    );

    bfr new_Jinkela_buffer_6472 (
        .din(new_Jinkela_wire_7898),
        .dout(new_Jinkela_wire_7899)
    );

    bfr new_Jinkela_buffer_943 (
        .din(new_Jinkela_wire_1013),
        .dout(new_Jinkela_wire_1014)
    );

    bfr new_Jinkela_buffer_6517 (
        .din(new_Jinkela_wire_7964),
        .dout(new_Jinkela_wire_7965)
    );

    bfr new_Jinkela_buffer_3146 (
        .din(new_Jinkela_wire_3598),
        .dout(new_Jinkela_wire_3599)
    );

    bfr new_Jinkela_buffer_6473 (
        .din(new_Jinkela_wire_7899),
        .dout(new_Jinkela_wire_7900)
    );

    bfr new_Jinkela_buffer_976 (
        .din(new_Jinkela_wire_1050),
        .dout(new_Jinkela_wire_1051)
    );

    bfr new_Jinkela_buffer_3158 (
        .din(new_Jinkela_wire_3612),
        .dout(new_Jinkela_wire_3613)
    );

    bfr new_Jinkela_buffer_944 (
        .din(new_Jinkela_wire_1014),
        .dout(new_Jinkela_wire_1015)
    );

    bfr new_Jinkela_buffer_3147 (
        .din(new_Jinkela_wire_3599),
        .dout(new_Jinkela_wire_3600)
    );

    bfr new_Jinkela_buffer_6474 (
        .din(new_Jinkela_wire_7900),
        .dout(new_Jinkela_wire_7901)
    );

    bfr new_Jinkela_buffer_1032 (
        .din(new_Jinkela_wire_1108),
        .dout(new_Jinkela_wire_1109)
    );

    bfr new_Jinkela_buffer_945 (
        .din(new_Jinkela_wire_1015),
        .dout(new_Jinkela_wire_1016)
    );

    spl4L new_Jinkela_splitter_159 (
        .a(n_1275_),
        .d(new_Jinkela_wire_3694),
        .b(new_Jinkela_wire_3695),
        .e(new_Jinkela_wire_3696),
        .c(new_Jinkela_wire_3697)
    );

    bfr new_Jinkela_buffer_6518 (
        .din(new_Jinkela_wire_7965),
        .dout(new_Jinkela_wire_7966)
    );

    bfr new_Jinkela_buffer_3148 (
        .din(new_Jinkela_wire_3600),
        .dout(new_Jinkela_wire_3601)
    );

    bfr new_Jinkela_buffer_6475 (
        .din(new_Jinkela_wire_7901),
        .dout(new_Jinkela_wire_7902)
    );

    bfr new_Jinkela_buffer_977 (
        .din(new_Jinkela_wire_1051),
        .dout(new_Jinkela_wire_1052)
    );

    bfr new_Jinkela_buffer_3159 (
        .din(new_Jinkela_wire_3613),
        .dout(new_Jinkela_wire_3614)
    );

    bfr new_Jinkela_buffer_946 (
        .din(new_Jinkela_wire_1016),
        .dout(new_Jinkela_wire_1017)
    );

    spl2 new_Jinkela_splitter_578 (
        .a(new_Jinkela_wire_8000),
        .b(new_Jinkela_wire_8001),
        .c(new_Jinkela_wire_8002)
    );

    bfr new_Jinkela_buffer_3149 (
        .din(new_Jinkela_wire_3601),
        .dout(new_Jinkela_wire_3602)
    );

    bfr new_Jinkela_buffer_6476 (
        .din(new_Jinkela_wire_7902),
        .dout(new_Jinkela_wire_7903)
    );

    bfr new_Jinkela_buffer_1224 (
        .din(new_Jinkela_wire_1542),
        .dout(new_Jinkela_wire_1543)
    );

    bfr new_Jinkela_buffer_3220 (
        .din(new_Jinkela_wire_3678),
        .dout(new_Jinkela_wire_3679)
    );

    bfr new_Jinkela_buffer_978 (
        .din(new_Jinkela_wire_1052),
        .dout(new_Jinkela_wire_1053)
    );

    spl2 new_Jinkela_splitter_160 (
        .a(n_0561_),
        .b(new_Jinkela_wire_3698),
        .c(new_Jinkela_wire_3699)
    );

    bfr new_Jinkela_buffer_6519 (
        .din(new_Jinkela_wire_7966),
        .dout(new_Jinkela_wire_7967)
    );

    bfr new_Jinkela_buffer_3150 (
        .din(new_Jinkela_wire_3602),
        .dout(new_Jinkela_wire_3603)
    );

    bfr new_Jinkela_buffer_6477 (
        .din(new_Jinkela_wire_7903),
        .dout(new_Jinkela_wire_7904)
    );

    bfr new_Jinkela_buffer_1288 (
        .din(N134),
        .dout(new_Jinkela_wire_1609)
    );

    bfr new_Jinkela_buffer_1033 (
        .din(new_Jinkela_wire_1109),
        .dout(new_Jinkela_wire_1110)
    );

    bfr new_Jinkela_buffer_3160 (
        .din(new_Jinkela_wire_3614),
        .dout(new_Jinkela_wire_3615)
    );

    bfr new_Jinkela_buffer_979 (
        .din(new_Jinkela_wire_1053),
        .dout(new_Jinkela_wire_1054)
    );

    bfr new_Jinkela_buffer_3151 (
        .din(new_Jinkela_wire_3603),
        .dout(new_Jinkela_wire_3604)
    );

    bfr new_Jinkela_buffer_6478 (
        .din(new_Jinkela_wire_7904),
        .dout(new_Jinkela_wire_7905)
    );

    bfr new_Jinkela_buffer_980 (
        .din(new_Jinkela_wire_1054),
        .dout(new_Jinkela_wire_1055)
    );

    bfr new_Jinkela_buffer_3233 (
        .din(n_0875_),
        .dout(new_Jinkela_wire_3700)
    );

    bfr new_Jinkela_buffer_6520 (
        .din(new_Jinkela_wire_7967),
        .dout(new_Jinkela_wire_7968)
    );

    bfr new_Jinkela_buffer_3152 (
        .din(new_Jinkela_wire_3604),
        .dout(new_Jinkela_wire_3605)
    );

    bfr new_Jinkela_buffer_6479 (
        .din(new_Jinkela_wire_7905),
        .dout(new_Jinkela_wire_7906)
    );

    bfr new_Jinkela_buffer_1034 (
        .din(new_Jinkela_wire_1110),
        .dout(new_Jinkela_wire_1111)
    );

    bfr new_Jinkela_buffer_3161 (
        .din(new_Jinkela_wire_3615),
        .dout(new_Jinkela_wire_3616)
    );

    bfr new_Jinkela_buffer_981 (
        .din(new_Jinkela_wire_1055),
        .dout(new_Jinkela_wire_1056)
    );

    bfr new_Jinkela_buffer_3153 (
        .din(new_Jinkela_wire_3605),
        .dout(new_Jinkela_wire_3606)
    );

    bfr new_Jinkela_buffer_6480 (
        .din(new_Jinkela_wire_7906),
        .dout(new_Jinkela_wire_7907)
    );

    bfr new_Jinkela_buffer_1095 (
        .din(new_Jinkela_wire_1401),
        .dout(new_Jinkela_wire_1402)
    );

    bfr new_Jinkela_buffer_3236 (
        .din(n_0283_),
        .dout(new_Jinkela_wire_3705)
    );

    bfr new_Jinkela_buffer_6542 (
        .din(new_Jinkela_wire_8003),
        .dout(new_Jinkela_wire_8004)
    );

    bfr new_Jinkela_buffer_982 (
        .din(new_Jinkela_wire_1056),
        .dout(new_Jinkela_wire_1057)
    );

    bfr new_Jinkela_buffer_3221 (
        .din(new_Jinkela_wire_3679),
        .dout(new_Jinkela_wire_3680)
    );

    bfr new_Jinkela_buffer_6521 (
        .din(new_Jinkela_wire_7968),
        .dout(new_Jinkela_wire_7969)
    );

    bfr new_Jinkela_buffer_3154 (
        .din(new_Jinkela_wire_3606),
        .dout(new_Jinkela_wire_3607)
    );

    bfr new_Jinkela_buffer_6481 (
        .din(new_Jinkela_wire_7907),
        .dout(new_Jinkela_wire_7908)
    );

    bfr new_Jinkela_buffer_1035 (
        .din(new_Jinkela_wire_1111),
        .dout(new_Jinkela_wire_1112)
    );

    bfr new_Jinkela_buffer_3162 (
        .din(new_Jinkela_wire_3616),
        .dout(new_Jinkela_wire_3617)
    );

    bfr new_Jinkela_buffer_983 (
        .din(new_Jinkela_wire_1057),
        .dout(new_Jinkela_wire_1058)
    );

    bfr new_Jinkela_buffer_3155 (
        .din(new_Jinkela_wire_3607),
        .dout(new_Jinkela_wire_3608)
    );

    bfr new_Jinkela_buffer_6482 (
        .din(new_Jinkela_wire_7908),
        .dout(new_Jinkela_wire_7909)
    );

    bfr new_Jinkela_buffer_1098 (
        .din(new_Jinkela_wire_1404),
        .dout(new_Jinkela_wire_1405)
    );

    bfr new_Jinkela_buffer_6543 (
        .din(new_Jinkela_wire_8004),
        .dout(new_Jinkela_wire_8005)
    );

    bfr new_Jinkela_buffer_984 (
        .din(new_Jinkela_wire_1058),
        .dout(new_Jinkela_wire_1059)
    );

    bfr new_Jinkela_buffer_6522 (
        .din(new_Jinkela_wire_7969),
        .dout(new_Jinkela_wire_7970)
    );

    bfr new_Jinkela_buffer_3156 (
        .din(new_Jinkela_wire_3608),
        .dout(new_Jinkela_wire_3609)
    );

    bfr new_Jinkela_buffer_6483 (
        .din(new_Jinkela_wire_7909),
        .dout(new_Jinkela_wire_7910)
    );

    bfr new_Jinkela_buffer_1036 (
        .din(new_Jinkela_wire_1112),
        .dout(new_Jinkela_wire_1113)
    );

    bfr new_Jinkela_buffer_3163 (
        .din(new_Jinkela_wire_3617),
        .dout(new_Jinkela_wire_3618)
    );

    bfr new_Jinkela_buffer_985 (
        .din(new_Jinkela_wire_1059),
        .dout(new_Jinkela_wire_1060)
    );

    bfr new_Jinkela_buffer_6547 (
        .din(new_Jinkela_wire_8010),
        .dout(new_Jinkela_wire_8011)
    );

    bfr new_Jinkela_buffer_3222 (
        .din(new_Jinkela_wire_3680),
        .dout(new_Jinkela_wire_3681)
    );

    bfr new_Jinkela_buffer_6484 (
        .din(new_Jinkela_wire_7910),
        .dout(new_Jinkela_wire_7911)
    );

    spl4L new_Jinkela_splitter_162 (
        .a(n_1201_),
        .d(new_Jinkela_wire_3712),
        .b(new_Jinkela_wire_3713),
        .e(new_Jinkela_wire_3714),
        .c(new_Jinkela_wire_3715)
    );

    spl2 new_Jinkela_splitter_98 (
        .a(N358),
        .b(new_Jinkela_wire_1541),
        .c(new_Jinkela_wire_1542)
    );

    bfr new_Jinkela_buffer_3164 (
        .din(new_Jinkela_wire_3618),
        .dout(new_Jinkela_wire_3619)
    );

    spl3L new_Jinkela_splitter_581 (
        .a(n_0017_),
        .d(new_Jinkela_wire_8071),
        .b(new_Jinkela_wire_8072),
        .c(new_Jinkela_wire_8073)
    );

    bfr new_Jinkela_buffer_986 (
        .din(new_Jinkela_wire_1060),
        .dout(new_Jinkela_wire_1061)
    );

    bfr new_Jinkela_buffer_6523 (
        .din(new_Jinkela_wire_7970),
        .dout(new_Jinkela_wire_7971)
    );

    bfr new_Jinkela_buffer_6485 (
        .din(new_Jinkela_wire_7911),
        .dout(new_Jinkela_wire_7912)
    );

    bfr new_Jinkela_buffer_1097 (
        .din(new_Jinkela_wire_1403),
        .dout(new_Jinkela_wire_1404)
    );

    bfr new_Jinkela_buffer_1037 (
        .din(new_Jinkela_wire_1113),
        .dout(new_Jinkela_wire_1114)
    );

    bfr new_Jinkela_buffer_3165 (
        .din(new_Jinkela_wire_3619),
        .dout(new_Jinkela_wire_3620)
    );

    bfr new_Jinkela_buffer_987 (
        .din(new_Jinkela_wire_1061),
        .dout(new_Jinkela_wire_1062)
    );

    spl2 new_Jinkela_splitter_582 (
        .a(n_1039_),
        .b(new_Jinkela_wire_8074),
        .c(new_Jinkela_wire_8075)
    );

    bfr new_Jinkela_buffer_6486 (
        .din(new_Jinkela_wire_7912),
        .dout(new_Jinkela_wire_7913)
    );

    bfr new_Jinkela_buffer_3223 (
        .din(new_Jinkela_wire_3681),
        .dout(new_Jinkela_wire_3682)
    );

    bfr new_Jinkela_buffer_3166 (
        .din(new_Jinkela_wire_3620),
        .dout(new_Jinkela_wire_3621)
    );

    bfr new_Jinkela_buffer_6544 (
        .din(new_Jinkela_wire_8005),
        .dout(new_Jinkela_wire_8006)
    );

    bfr new_Jinkela_buffer_988 (
        .din(new_Jinkela_wire_1062),
        .dout(new_Jinkela_wire_1063)
    );

    bfr new_Jinkela_buffer_6524 (
        .din(new_Jinkela_wire_7971),
        .dout(new_Jinkela_wire_7972)
    );

    spl2 new_Jinkela_splitter_564 (
        .a(new_Jinkela_wire_7913),
        .b(new_Jinkela_wire_7914),
        .c(new_Jinkela_wire_7915)
    );

    bfr new_Jinkela_buffer_1161 (
        .din(new_Jinkela_wire_1472),
        .dout(new_Jinkela_wire_1473)
    );

    bfr new_Jinkela_buffer_3234 (
        .din(new_Jinkela_wire_3700),
        .dout(new_Jinkela_wire_3701)
    );

    bfr new_Jinkela_buffer_1038 (
        .din(new_Jinkela_wire_1114),
        .dout(new_Jinkela_wire_1115)
    );

    bfr new_Jinkela_buffer_3167 (
        .din(new_Jinkela_wire_3621),
        .dout(new_Jinkela_wire_3622)
    );

    bfr new_Jinkela_buffer_8415 (
        .din(new_Jinkela_wire_10580),
        .dout(new_Jinkela_wire_10581)
    );

    bfr new_Jinkela_buffer_8416 (
        .din(new_Jinkela_wire_10581),
        .dout(new_Jinkela_wire_10582)
    );

    bfr new_Jinkela_buffer_8417 (
        .din(new_Jinkela_wire_10582),
        .dout(new_Jinkela_wire_10583)
    );

    bfr new_Jinkela_buffer_8418 (
        .din(new_Jinkela_wire_10583),
        .dout(new_Jinkela_wire_10584)
    );

    bfr new_Jinkela_buffer_8419 (
        .din(new_Jinkela_wire_10584),
        .dout(new_Jinkela_wire_10585)
    );

    bfr new_Jinkela_buffer_8420 (
        .din(new_Jinkela_wire_10585),
        .dout(new_Jinkela_wire_10586)
    );

    spl3L new_Jinkela_splitter_569 (
        .a(n_0667_),
        .d(new_Jinkela_wire_7929),
        .b(new_Jinkela_wire_7930),
        .c(new_Jinkela_wire_7931)
    );

    bfr new_Jinkela_buffer_8421 (
        .din(new_Jinkela_wire_10586),
        .dout(new_Jinkela_wire_10587)
    );

    bfr new_Jinkela_buffer_8422 (
        .din(new_Jinkela_wire_10587),
        .dout(new_Jinkela_wire_10588)
    );

    bfr new_Jinkela_buffer_8423 (
        .din(new_Jinkela_wire_10588),
        .dout(new_Jinkela_wire_10589)
    );

    bfr new_Jinkela_buffer_8424 (
        .din(new_Jinkela_wire_10589),
        .dout(new_Jinkela_wire_10590)
    );

    bfr new_Jinkela_buffer_8425 (
        .din(new_Jinkela_wire_10590),
        .dout(new_Jinkela_wire_10591)
    );

    bfr new_Jinkela_buffer_8426 (
        .din(new_Jinkela_wire_10591),
        .dout(new_Jinkela_wire_10592)
    );

    bfr new_Jinkela_buffer_8427 (
        .din(new_Jinkela_wire_10592),
        .dout(new_Jinkela_wire_10593)
    );

    bfr new_Jinkela_buffer_8428 (
        .din(new_Jinkela_wire_10593),
        .dout(new_Jinkela_wire_10594)
    );

    bfr new_Jinkela_buffer_8429 (
        .din(new_Jinkela_wire_10594),
        .dout(new_Jinkela_wire_10595)
    );

    bfr new_Jinkela_buffer_8430 (
        .din(new_Jinkela_wire_10595),
        .dout(new_Jinkela_wire_10596)
    );

    bfr new_Jinkela_buffer_8431 (
        .din(new_Jinkela_wire_10596),
        .dout(new_Jinkela_wire_10597)
    );

    bfr new_Jinkela_buffer_8432 (
        .din(new_Jinkela_wire_10597),
        .dout(new_Jinkela_wire_10598)
    );

    bfr new_Jinkela_buffer_8433 (
        .din(new_Jinkela_wire_10598),
        .dout(new_Jinkela_wire_10599)
    );

    bfr new_Jinkela_buffer_8434 (
        .din(new_Jinkela_wire_10599),
        .dout(new_Jinkela_wire_10600)
    );

    bfr new_Jinkela_buffer_8435 (
        .din(new_Jinkela_wire_10600),
        .dout(new_Jinkela_wire_10601)
    );

    and_bb n_1737_ (
        .a(new_Jinkela_wire_8296),
        .b(new_Jinkela_wire_4430),
        .c(n_1004_)
    );

    and_bi n_2451_ (
        .a(new_Jinkela_wire_7842),
        .b(new_Jinkela_wire_7204),
        .c(n_0326_)
    );

    and_bi n_1738_ (
        .a(n_1003_),
        .b(n_1004_),
        .c(n_1005_)
    );

    and_bi n_2452_ (
        .a(new_Jinkela_wire_9754),
        .b(new_Jinkela_wire_7745),
        .c(n_0327_)
    );

    or_bb n_1739_ (
        .a(n_1005_),
        .b(new_Jinkela_wire_10221),
        .c(n_1006_)
    );

    or_bb n_2453_ (
        .a(new_Jinkela_wire_8366),
        .b(new_Jinkela_wire_5063),
        .c(n_0328_)
    );

    and_bi n_1740_ (
        .a(new_Jinkela_wire_1686),
        .b(new_Jinkela_wire_1363),
        .c(n_1007_)
    );

    or_bb n_2454_ (
        .a(n_0328_),
        .b(new_Jinkela_wire_6187),
        .c(n_0329_)
    );

    and_bi n_1741_ (
        .a(new_Jinkela_wire_1276),
        .b(new_Jinkela_wire_2381),
        .c(n_1008_)
    );

    and_ii n_2455_ (
        .a(n_0329_),
        .b(new_Jinkela_wire_7836),
        .c(n_0330_)
    );

    and_ii n_1742_ (
        .a(n_1008_),
        .b(n_1007_),
        .c(n_1009_)
    );

    or_ii n_2456_ (
        .a(new_Jinkela_wire_8322),
        .b(new_Jinkela_wire_4863),
        .c(n_0331_)
    );

    and_bi n_1743_ (
        .a(new_Jinkela_wire_1786),
        .b(new_Jinkela_wire_1196),
        .c(n_1010_)
    );

    or_bb n_2457_ (
        .a(new_Jinkela_wire_3834),
        .b(n_0312_),
        .c(n_0332_)
    );

    and_bi n_1744_ (
        .a(new_Jinkela_wire_1269),
        .b(new_Jinkela_wire_515),
        .c(n_1011_)
    );

    or_bi n_2458_ (
        .a(new_Jinkela_wire_8368),
        .b(new_Jinkela_wire_7834),
        .c(n_0333_)
    );

    and_ii n_1745_ (
        .a(n_1011_),
        .b(n_1010_),
        .c(n_1012_)
    );

    and_bi n_2459_ (
        .a(n_0333_),
        .b(new_Jinkela_wire_5066),
        .c(n_0334_)
    );

    or_bb n_1746_ (
        .a(new_Jinkela_wire_7999),
        .b(new_Jinkela_wire_8271),
        .c(n_1013_)
    );

    and_bi n_2460_ (
        .a(new_Jinkela_wire_4862),
        .b(new_Jinkela_wire_9149),
        .c(n_0335_)
    );

    and_bb n_1747_ (
        .a(new_Jinkela_wire_7998),
        .b(new_Jinkela_wire_8270),
        .c(n_1014_)
    );

    and_bi n_2461_ (
        .a(new_Jinkela_wire_3523),
        .b(new_Jinkela_wire_5150),
        .c(n_0336_)
    );

    and_bi n_1748_ (
        .a(n_1013_),
        .b(n_1014_),
        .c(n_1015_)
    );

    and_bi n_2462_ (
        .a(new_Jinkela_wire_354),
        .b(n_0336_),
        .c(n_0337_)
    );

    and_bi n_1749_ (
        .a(new_Jinkela_wire_3193),
        .b(new_Jinkela_wire_1282),
        .c(n_1016_)
    );

    or_bb n_2463_ (
        .a(new_Jinkela_wire_3726),
        .b(new_Jinkela_wire_6706),
        .c(n_0338_)
    );

    and_bi n_1750_ (
        .a(new_Jinkela_wire_1189),
        .b(new_Jinkela_wire_804),
        .c(n_1017_)
    );

    and_bi n_2464_ (
        .a(n_0338_),
        .b(new_Jinkela_wire_8573),
        .c(n_0339_)
    );

    and_ii n_1751_ (
        .a(n_1017_),
        .b(n_1016_),
        .c(n_1018_)
    );

    or_bb n_2465_ (
        .a(n_0339_),
        .b(new_Jinkela_wire_9616),
        .c(n_0340_)
    );

    and_bi n_1752_ (
        .a(new_Jinkela_wire_2551),
        .b(new_Jinkela_wire_1209),
        .c(n_1019_)
    );

    or_bb n_2466_ (
        .a(new_Jinkela_wire_6249),
        .b(n_0335_),
        .c(n_0341_)
    );

    and_bi n_1753_ (
        .a(new_Jinkela_wire_1248),
        .b(new_Jinkela_wire_1022),
        .c(n_1020_)
    );

    and_bi n_2467_ (
        .a(n_0332_),
        .b(new_Jinkela_wire_5248),
        .c(n_0342_)
    );

    and_ii n_1754_ (
        .a(n_1020_),
        .b(n_1019_),
        .c(n_1021_)
    );

    and_bi n_2468_ (
        .a(new_Jinkela_wire_8436),
        .b(new_Jinkela_wire_3676),
        .c(new_net_7)
    );

    and_bi n_1755_ (
        .a(new_Jinkela_wire_3950),
        .b(new_Jinkela_wire_5283),
        .c(n_1022_)
    );

    inv n_2469_ (
        .din(new_Jinkela_wire_5880),
        .dout(n_0343_)
    );

    and_bi n_1756_ (
        .a(new_Jinkela_wire_5282),
        .b(new_Jinkela_wire_3949),
        .c(n_1023_)
    );

    or_bb n_2470_ (
        .a(new_Jinkela_wire_4050),
        .b(new_Jinkela_wire_3728),
        .c(n_0344_)
    );

    or_bi n_2471_ (
        .a(new_Jinkela_wire_7216),
        .b(new_Jinkela_wire_9708),
        .c(n_0345_)
    );

    and_ii n_1757_ (
        .a(n_1023_),
        .b(n_1022_),
        .c(n_1024_)
    );

    or_bi n_1758_ (
        .a(new_Jinkela_wire_9762),
        .b(new_Jinkela_wire_5001),
        .c(n_1025_)
    );

    and_bi n_2472_ (
        .a(n_0345_),
        .b(new_Jinkela_wire_6151),
        .c(n_0346_)
    );

    and_bi n_1759_ (
        .a(new_Jinkela_wire_9761),
        .b(new_Jinkela_wire_5000),
        .c(n_1026_)
    );

    or_ii n_2473_ (
        .a(new_Jinkela_wire_8442),
        .b(new_Jinkela_wire_6766),
        .c(n_0347_)
    );

    and_bi n_1760_ (
        .a(n_1025_),
        .b(n_1026_),
        .c(n_1027_)
    );

    or_bb n_2474_ (
        .a(new_Jinkela_wire_8441),
        .b(new_Jinkela_wire_6765),
        .c(n_0348_)
    );

    and_bi n_1761_ (
        .a(new_Jinkela_wire_1097),
        .b(new_Jinkela_wire_1321),
        .c(n_1028_)
    );

    or_ii n_2475_ (
        .a(n_0348_),
        .b(n_0347_),
        .c(new_net_2501)
    );

    and_bi n_2476_ (
        .a(new_Jinkela_wire_9706),
        .b(new_Jinkela_wire_9365),
        .c(n_0349_)
    );

    and_bi n_1762_ (
        .a(new_Jinkela_wire_1375),
        .b(new_Jinkela_wire_109),
        .c(n_1029_)
    );

    and_ii n_1763_ (
        .a(n_1029_),
        .b(n_1028_),
        .c(n_1030_)
    );

    or_ii n_2477_ (
        .a(new_Jinkela_wire_7068),
        .b(new_Jinkela_wire_10522),
        .c(n_0350_)
    );

    and_bi n_1764_ (
        .a(new_Jinkela_wire_344),
        .b(new_Jinkela_wire_1252),
        .c(n_1031_)
    );

    and_bi n_2478_ (
        .a(n_0350_),
        .b(new_Jinkela_wire_8532),
        .c(n_0351_)
    );

    and_bi n_1765_ (
        .a(new_Jinkela_wire_1295),
        .b(new_Jinkela_wire_204),
        .c(n_1032_)
    );

    and_bi n_2479_ (
        .a(new_Jinkela_wire_9376),
        .b(new_Jinkela_wire_4069),
        .c(n_0352_)
    );

    and_ii n_1766_ (
        .a(n_1032_),
        .b(n_1031_),
        .c(n_1033_)
    );

    and_bi n_2480_ (
        .a(new_Jinkela_wire_4068),
        .b(new_Jinkela_wire_9375),
        .c(n_0353_)
    );

    or_bb n_2481_ (
        .a(n_0353_),
        .b(n_0352_),
        .c(new_net_2515)
    );

    and_ii n_1767_ (
        .a(new_Jinkela_wire_6336),
        .b(new_Jinkela_wire_4516),
        .c(n_1034_)
    );

    and_bb n_1768_ (
        .a(new_Jinkela_wire_6335),
        .b(new_Jinkela_wire_4515),
        .c(n_1035_)
    );

    inv n_2482_ (
        .din(new_Jinkela_wire_10502),
        .dout(n_0354_)
    );

    and_ii n_1769_ (
        .a(n_1035_),
        .b(n_1034_),
        .c(n_1036_)
    );

    and_ii n_2483_ (
        .a(new_Jinkela_wire_7067),
        .b(new_Jinkela_wire_6427),
        .c(n_0355_)
    );

    or_bi n_1770_ (
        .a(new_Jinkela_wire_10379),
        .b(new_Jinkela_wire_5396),
        .c(n_1037_)
    );

    and_bi n_2484_ (
        .a(new_Jinkela_wire_9038),
        .b(new_Jinkela_wire_9640),
        .c(n_0356_)
    );

    and_bi n_1771_ (
        .a(new_Jinkela_wire_10378),
        .b(new_Jinkela_wire_5395),
        .c(n_1038_)
    );

    and_bi n_2485_ (
        .a(new_Jinkela_wire_9639),
        .b(new_Jinkela_wire_9037),
        .c(n_0357_)
    );

    or_bb n_2486_ (
        .a(n_0357_),
        .b(n_0356_),
        .c(new_net_2535)
    );

    and_bi n_1772_ (
        .a(n_1037_),
        .b(n_1038_),
        .c(n_1039_)
    );

    and_bi n_1773_ (
        .a(new_Jinkela_wire_1698),
        .b(new_Jinkela_wire_1177),
        .c(n_1040_)
    );

    and_bi n_2487_ (
        .a(new_Jinkela_wire_9707),
        .b(new_Jinkela_wire_9133),
        .c(n_0358_)
    );

    and_bi n_1774_ (
        .a(new_Jinkela_wire_1284),
        .b(new_Jinkela_wire_2310),
        .c(n_1041_)
    );

    and_bi n_2488_ (
        .a(new_Jinkela_wire_9134),
        .b(new_Jinkela_wire_9704),
        .c(n_0359_)
    );

    and_ii n_1775_ (
        .a(n_1041_),
        .b(n_1040_),
        .c(n_1042_)
    );

    or_bb n_2489_ (
        .a(n_0359_),
        .b(n_0358_),
        .c(new_net_2493)
    );

    and_bi n_1776_ (
        .a(new_Jinkela_wire_2975),
        .b(new_Jinkela_wire_1262),
        .c(n_1043_)
    );

    inv n_2490_ (
        .din(new_Jinkela_wire_6804),
        .dout(new_net_2570)
    );

    and_ii n_2491_ (
        .a(new_Jinkela_wire_5458),
        .b(new_Jinkela_wire_8767),
        .c(n_0360_)
    );

    and_bi n_1777_ (
        .a(new_Jinkela_wire_1230),
        .b(new_Jinkela_wire_1545),
        .c(n_1044_)
    );

    and_bi n_2492_ (
        .a(new_Jinkela_wire_4433),
        .b(new_Jinkela_wire_6886),
        .c(n_0361_)
    );

    and_ii n_1778_ (
        .a(n_1044_),
        .b(n_1043_),
        .c(n_1045_)
    );

    bfr new_Jinkela_buffer_2349 (
        .din(new_Jinkela_wire_2742),
        .dout(new_Jinkela_wire_2743)
    );

    bfr new_Jinkela_buffer_7478 (
        .din(new_Jinkela_wire_9304),
        .dout(new_Jinkela_wire_9305)
    );

    bfr new_Jinkela_buffer_2244 (
        .din(new_Jinkela_wire_2630),
        .dout(new_Jinkela_wire_2631)
    );

    bfr new_Jinkela_buffer_7420 (
        .din(new_Jinkela_wire_9223),
        .dout(new_Jinkela_wire_9224)
    );

    bfr new_Jinkela_buffer_2291 (
        .din(new_Jinkela_wire_2682),
        .dout(new_Jinkela_wire_2683)
    );

    bfr new_Jinkela_buffer_7449 (
        .din(new_Jinkela_wire_9263),
        .dout(new_Jinkela_wire_9264)
    );

    bfr new_Jinkela_buffer_2245 (
        .din(new_Jinkela_wire_2631),
        .dout(new_Jinkela_wire_2632)
    );

    bfr new_Jinkela_buffer_7421 (
        .din(new_Jinkela_wire_9224),
        .dout(new_Jinkela_wire_9225)
    );

    bfr new_Jinkela_buffer_2420 (
        .din(N251),
        .dout(new_Jinkela_wire_2817)
    );

    bfr new_Jinkela_buffer_2246 (
        .din(new_Jinkela_wire_2632),
        .dout(new_Jinkela_wire_2633)
    );

    bfr new_Jinkela_buffer_7509 (
        .din(new_Jinkela_wire_9337),
        .dout(new_Jinkela_wire_9338)
    );

    bfr new_Jinkela_buffer_7422 (
        .din(new_Jinkela_wire_9225),
        .dout(new_Jinkela_wire_9226)
    );

    bfr new_Jinkela_buffer_2292 (
        .din(new_Jinkela_wire_2683),
        .dout(new_Jinkela_wire_2684)
    );

    bfr new_Jinkela_buffer_7450 (
        .din(new_Jinkela_wire_9264),
        .dout(new_Jinkela_wire_9265)
    );

    bfr new_Jinkela_buffer_2247 (
        .din(new_Jinkela_wire_2633),
        .dout(new_Jinkela_wire_2634)
    );

    bfr new_Jinkela_buffer_7423 (
        .din(new_Jinkela_wire_9226),
        .dout(new_Jinkela_wire_9227)
    );

    spl3L new_Jinkela_splitter_132 (
        .a(new_Jinkela_wire_2743),
        .d(new_Jinkela_wire_2744),
        .b(new_Jinkela_wire_2745),
        .c(new_Jinkela_wire_2746)
    );

    bfr new_Jinkela_buffer_7479 (
        .din(new_Jinkela_wire_9305),
        .dout(new_Jinkela_wire_9306)
    );

    bfr new_Jinkela_buffer_2248 (
        .din(new_Jinkela_wire_2634),
        .dout(new_Jinkela_wire_2635)
    );

    bfr new_Jinkela_buffer_7424 (
        .din(new_Jinkela_wire_9227),
        .dout(new_Jinkela_wire_9228)
    );

    bfr new_Jinkela_buffer_2293 (
        .din(new_Jinkela_wire_2684),
        .dout(new_Jinkela_wire_2685)
    );

    bfr new_Jinkela_buffer_7451 (
        .din(new_Jinkela_wire_9265),
        .dout(new_Jinkela_wire_9266)
    );

    bfr new_Jinkela_buffer_2249 (
        .din(new_Jinkela_wire_2635),
        .dout(new_Jinkela_wire_2636)
    );

    bfr new_Jinkela_buffer_7425 (
        .din(new_Jinkela_wire_9228),
        .dout(new_Jinkela_wire_9229)
    );

    bfr new_Jinkela_buffer_2414 (
        .din(new_Jinkela_wire_2810),
        .dout(new_Jinkela_wire_2811)
    );

    bfr new_Jinkela_buffer_7510 (
        .din(n_0259_),
        .dout(new_Jinkela_wire_9344)
    );

    bfr new_Jinkela_buffer_2250 (
        .din(new_Jinkela_wire_2636),
        .dout(new_Jinkela_wire_2637)
    );

    bfr new_Jinkela_buffer_7426 (
        .din(new_Jinkela_wire_9229),
        .dout(new_Jinkela_wire_9230)
    );

    bfr new_Jinkela_buffer_2294 (
        .din(new_Jinkela_wire_2685),
        .dout(new_Jinkela_wire_2686)
    );

    bfr new_Jinkela_buffer_7452 (
        .din(new_Jinkela_wire_9266),
        .dout(new_Jinkela_wire_9267)
    );

    bfr new_Jinkela_buffer_2251 (
        .din(new_Jinkela_wire_2637),
        .dout(new_Jinkela_wire_2638)
    );

    bfr new_Jinkela_buffer_7427 (
        .din(new_Jinkela_wire_9230),
        .dout(new_Jinkela_wire_9231)
    );

    bfr new_Jinkela_buffer_2350 (
        .din(new_Jinkela_wire_2746),
        .dout(new_Jinkela_wire_2747)
    );

    bfr new_Jinkela_buffer_7480 (
        .din(new_Jinkela_wire_9306),
        .dout(new_Jinkela_wire_9307)
    );

    bfr new_Jinkela_buffer_2252 (
        .din(new_Jinkela_wire_2638),
        .dout(new_Jinkela_wire_2639)
    );

    bfr new_Jinkela_buffer_7428 (
        .din(new_Jinkela_wire_9231),
        .dout(new_Jinkela_wire_9232)
    );

    bfr new_Jinkela_buffer_2295 (
        .din(new_Jinkela_wire_2686),
        .dout(new_Jinkela_wire_2687)
    );

    bfr new_Jinkela_buffer_7453 (
        .din(new_Jinkela_wire_9267),
        .dout(new_Jinkela_wire_9268)
    );

    bfr new_Jinkela_buffer_2253 (
        .din(new_Jinkela_wire_2639),
        .dout(new_Jinkela_wire_2640)
    );

    bfr new_Jinkela_buffer_7429 (
        .din(new_Jinkela_wire_9232),
        .dout(new_Jinkela_wire_9233)
    );

    bfr new_Jinkela_buffer_2417 (
        .din(new_Jinkela_wire_2813),
        .dout(new_Jinkela_wire_2814)
    );

    bfr new_Jinkela_buffer_2254 (
        .din(new_Jinkela_wire_2640),
        .dout(new_Jinkela_wire_2641)
    );

    spl2 new_Jinkela_splitter_737 (
        .a(n_1369_),
        .b(new_Jinkela_wire_9345),
        .c(new_Jinkela_wire_9346)
    );

    bfr new_Jinkela_buffer_7430 (
        .din(new_Jinkela_wire_9233),
        .dout(new_Jinkela_wire_9234)
    );

    bfr new_Jinkela_buffer_2296 (
        .din(new_Jinkela_wire_2687),
        .dout(new_Jinkela_wire_2688)
    );

    bfr new_Jinkela_buffer_7454 (
        .din(new_Jinkela_wire_9268),
        .dout(new_Jinkela_wire_9269)
    );

    bfr new_Jinkela_buffer_2255 (
        .din(new_Jinkela_wire_2641),
        .dout(new_Jinkela_wire_2642)
    );

    bfr new_Jinkela_buffer_7431 (
        .din(new_Jinkela_wire_9234),
        .dout(new_Jinkela_wire_9235)
    );

    bfr new_Jinkela_buffer_2351 (
        .din(new_Jinkela_wire_2747),
        .dout(new_Jinkela_wire_2748)
    );

    bfr new_Jinkela_buffer_7481 (
        .din(new_Jinkela_wire_9307),
        .dout(new_Jinkela_wire_9308)
    );

    bfr new_Jinkela_buffer_2256 (
        .din(new_Jinkela_wire_2642),
        .dout(new_Jinkela_wire_2643)
    );

    bfr new_Jinkela_buffer_7432 (
        .din(new_Jinkela_wire_9235),
        .dout(new_Jinkela_wire_9236)
    );

    bfr new_Jinkela_buffer_2297 (
        .din(new_Jinkela_wire_2688),
        .dout(new_Jinkela_wire_2689)
    );

    bfr new_Jinkela_buffer_7455 (
        .din(new_Jinkela_wire_9269),
        .dout(new_Jinkela_wire_9270)
    );

    bfr new_Jinkela_buffer_2257 (
        .din(new_Jinkela_wire_2643),
        .dout(new_Jinkela_wire_2644)
    );

    bfr new_Jinkela_buffer_7433 (
        .din(new_Jinkela_wire_9236),
        .dout(new_Jinkela_wire_9237)
    );

    bfr new_Jinkela_buffer_2415 (
        .din(new_Jinkela_wire_2811),
        .dout(new_Jinkela_wire_2812)
    );

    bfr new_Jinkela_buffer_2258 (
        .din(new_Jinkela_wire_2644),
        .dout(new_Jinkela_wire_2645)
    );

    spl2 new_Jinkela_splitter_740 (
        .a(n_0771_),
        .b(new_Jinkela_wire_9366),
        .c(new_Jinkela_wire_9367)
    );

    bfr new_Jinkela_buffer_7434 (
        .din(new_Jinkela_wire_9237),
        .dout(new_Jinkela_wire_9238)
    );

    bfr new_Jinkela_buffer_2298 (
        .din(new_Jinkela_wire_2689),
        .dout(new_Jinkela_wire_2690)
    );

    bfr new_Jinkela_buffer_7456 (
        .din(new_Jinkela_wire_9270),
        .dout(new_Jinkela_wire_9271)
    );

    bfr new_Jinkela_buffer_2259 (
        .din(new_Jinkela_wire_2645),
        .dout(new_Jinkela_wire_2646)
    );

    bfr new_Jinkela_buffer_7435 (
        .din(new_Jinkela_wire_9238),
        .dout(new_Jinkela_wire_9239)
    );

    bfr new_Jinkela_buffer_2352 (
        .din(new_Jinkela_wire_2748),
        .dout(new_Jinkela_wire_2749)
    );

    bfr new_Jinkela_buffer_7482 (
        .din(new_Jinkela_wire_9308),
        .dout(new_Jinkela_wire_9309)
    );

    bfr new_Jinkela_buffer_2260 (
        .din(new_Jinkela_wire_2646),
        .dout(new_Jinkela_wire_2647)
    );

    bfr new_Jinkela_buffer_7436 (
        .din(new_Jinkela_wire_9239),
        .dout(new_Jinkela_wire_9240)
    );

    bfr new_Jinkela_buffer_2299 (
        .din(new_Jinkela_wire_2690),
        .dout(new_Jinkela_wire_2691)
    );

    bfr new_Jinkela_buffer_7457 (
        .din(new_Jinkela_wire_9271),
        .dout(new_Jinkela_wire_9272)
    );

    bfr new_Jinkela_buffer_2261 (
        .din(new_Jinkela_wire_2647),
        .dout(new_Jinkela_wire_2648)
    );

    bfr new_Jinkela_buffer_7437 (
        .din(new_Jinkela_wire_9240),
        .dout(new_Jinkela_wire_9241)
    );

    bfr new_Jinkela_buffer_2484 (
        .din(N103),
        .dout(new_Jinkela_wire_2886)
    );

    spl2 new_Jinkela_splitter_735 (
        .a(new_Jinkela_wire_9338),
        .b(new_Jinkela_wire_9339),
        .c(new_Jinkela_wire_9340)
    );

    bfr new_Jinkela_buffer_2262 (
        .din(new_Jinkela_wire_2648),
        .dout(new_Jinkela_wire_2649)
    );

    bfr new_Jinkela_buffer_7438 (
        .din(new_Jinkela_wire_9241),
        .dout(new_Jinkela_wire_9242)
    );

    bfr new_Jinkela_buffer_2300 (
        .din(new_Jinkela_wire_2691),
        .dout(new_Jinkela_wire_2692)
    );

    bfr new_Jinkela_buffer_7458 (
        .din(new_Jinkela_wire_9272),
        .dout(new_Jinkela_wire_9273)
    );

    bfr new_Jinkela_buffer_2263 (
        .din(new_Jinkela_wire_2649),
        .dout(new_Jinkela_wire_2650)
    );

    bfr new_Jinkela_buffer_7439 (
        .din(new_Jinkela_wire_9242),
        .dout(new_Jinkela_wire_9243)
    );

    bfr new_Jinkela_buffer_2353 (
        .din(new_Jinkela_wire_2749),
        .dout(new_Jinkela_wire_2750)
    );

    bfr new_Jinkela_buffer_7483 (
        .din(new_Jinkela_wire_9309),
        .dout(new_Jinkela_wire_9310)
    );

    bfr new_Jinkela_buffer_2264 (
        .din(new_Jinkela_wire_2650),
        .dout(new_Jinkela_wire_2651)
    );

    spl2 new_Jinkela_splitter_724 (
        .a(new_Jinkela_wire_9243),
        .b(new_Jinkela_wire_9244),
        .c(new_Jinkela_wire_9245)
    );

    bfr new_Jinkela_buffer_4845 (
        .din(new_Jinkela_wire_5779),
        .dout(new_Jinkela_wire_5780)
    );

    spl2 new_Jinkela_splitter_163 (
        .a(n_1176_),
        .b(new_Jinkela_wire_3716),
        .c(new_Jinkela_wire_3717)
    );

    bfr new_Jinkela_buffer_1646 (
        .din(N213),
        .dout(new_Jinkela_wire_1990)
    );

    bfr new_Jinkela_buffer_3993 (
        .din(new_Jinkela_wire_4689),
        .dout(new_Jinkela_wire_4690)
    );

    bfr new_Jinkela_buffer_3224 (
        .din(new_Jinkela_wire_3682),
        .dout(new_Jinkela_wire_3683)
    );

    bfr new_Jinkela_buffer_3168 (
        .din(new_Jinkela_wire_3622),
        .dout(new_Jinkela_wire_3623)
    );

    bfr new_Jinkela_buffer_1522 (
        .din(new_Jinkela_wire_1859),
        .dout(new_Jinkela_wire_1860)
    );

    bfr new_Jinkela_buffer_4880 (
        .din(new_Jinkela_wire_5816),
        .dout(new_Jinkela_wire_5817)
    );

    bfr new_Jinkela_buffer_4846 (
        .din(new_Jinkela_wire_5780),
        .dout(new_Jinkela_wire_5781)
    );

    bfr new_Jinkela_buffer_4044 (
        .din(new_Jinkela_wire_4742),
        .dout(new_Jinkela_wire_4743)
    );

    bfr new_Jinkela_buffer_1575 (
        .din(new_Jinkela_wire_1918),
        .dout(new_Jinkela_wire_1919)
    );

    bfr new_Jinkela_buffer_3994 (
        .din(new_Jinkela_wire_4690),
        .dout(new_Jinkela_wire_4691)
    );

    bfr new_Jinkela_buffer_3237 (
        .din(new_Jinkela_wire_3705),
        .dout(new_Jinkela_wire_3706)
    );

    bfr new_Jinkela_buffer_3169 (
        .din(new_Jinkela_wire_3623),
        .dout(new_Jinkela_wire_3624)
    );

    bfr new_Jinkela_buffer_1523 (
        .din(new_Jinkela_wire_1860),
        .dout(new_Jinkela_wire_1861)
    );

    bfr new_Jinkela_buffer_4937 (
        .din(new_Jinkela_wire_5886),
        .dout(new_Jinkela_wire_5887)
    );

    bfr new_Jinkela_buffer_4847 (
        .din(new_Jinkela_wire_5781),
        .dout(new_Jinkela_wire_5782)
    );

    bfr new_Jinkela_buffer_4084 (
        .din(new_Jinkela_wire_4784),
        .dout(new_Jinkela_wire_4785)
    );

    bfr new_Jinkela_buffer_3235 (
        .din(new_Jinkela_wire_3701),
        .dout(new_Jinkela_wire_3702)
    );

    bfr new_Jinkela_buffer_1640 (
        .din(new_Jinkela_wire_1983),
        .dout(new_Jinkela_wire_1984)
    );

    bfr new_Jinkela_buffer_3995 (
        .din(new_Jinkela_wire_4691),
        .dout(new_Jinkela_wire_4692)
    );

    bfr new_Jinkela_buffer_3225 (
        .din(new_Jinkela_wire_3683),
        .dout(new_Jinkela_wire_3684)
    );

    bfr new_Jinkela_buffer_3170 (
        .din(new_Jinkela_wire_3624),
        .dout(new_Jinkela_wire_3625)
    );

    bfr new_Jinkela_buffer_1524 (
        .din(new_Jinkela_wire_1861),
        .dout(new_Jinkela_wire_1862)
    );

    bfr new_Jinkela_buffer_4881 (
        .din(new_Jinkela_wire_5817),
        .dout(new_Jinkela_wire_5818)
    );

    bfr new_Jinkela_buffer_4848 (
        .din(new_Jinkela_wire_5782),
        .dout(new_Jinkela_wire_5783)
    );

    bfr new_Jinkela_buffer_4045 (
        .din(new_Jinkela_wire_4743),
        .dout(new_Jinkela_wire_4744)
    );

    bfr new_Jinkela_buffer_1576 (
        .din(new_Jinkela_wire_1919),
        .dout(new_Jinkela_wire_1920)
    );

    bfr new_Jinkela_buffer_3996 (
        .din(new_Jinkela_wire_4692),
        .dout(new_Jinkela_wire_4693)
    );

    bfr new_Jinkela_buffer_3171 (
        .din(new_Jinkela_wire_3625),
        .dout(new_Jinkela_wire_3626)
    );

    bfr new_Jinkela_buffer_1525 (
        .din(new_Jinkela_wire_1862),
        .dout(new_Jinkela_wire_1863)
    );

    bfr new_Jinkela_buffer_4968 (
        .din(new_Jinkela_wire_5919),
        .dout(new_Jinkela_wire_5920)
    );

    bfr new_Jinkela_buffer_4849 (
        .din(new_Jinkela_wire_5783),
        .dout(new_Jinkela_wire_5784)
    );

    spl2 new_Jinkela_splitter_261 (
        .a(n_1248_),
        .b(new_Jinkela_wire_4856),
        .c(new_Jinkela_wire_4857)
    );

    bfr new_Jinkela_buffer_4118 (
        .din(new_Jinkela_wire_4818),
        .dout(new_Jinkela_wire_4819)
    );

    bfr new_Jinkela_buffer_1643 (
        .din(new_Jinkela_wire_1986),
        .dout(new_Jinkela_wire_1987)
    );

    bfr new_Jinkela_buffer_3997 (
        .din(new_Jinkela_wire_4693),
        .dout(new_Jinkela_wire_4694)
    );

    spl2 new_Jinkela_splitter_158 (
        .a(new_Jinkela_wire_3684),
        .b(new_Jinkela_wire_3685),
        .c(new_Jinkela_wire_3686)
    );

    bfr new_Jinkela_buffer_3172 (
        .din(new_Jinkela_wire_3626),
        .dout(new_Jinkela_wire_3627)
    );

    bfr new_Jinkela_buffer_1526 (
        .din(new_Jinkela_wire_1863),
        .dout(new_Jinkela_wire_1864)
    );

    bfr new_Jinkela_buffer_4882 (
        .din(new_Jinkela_wire_5818),
        .dout(new_Jinkela_wire_5819)
    );

    bfr new_Jinkela_buffer_4945 (
        .din(new_Jinkela_wire_5894),
        .dout(new_Jinkela_wire_5895)
    );

    bfr new_Jinkela_buffer_4850 (
        .din(new_Jinkela_wire_5784),
        .dout(new_Jinkela_wire_5785)
    );

    bfr new_Jinkela_buffer_4046 (
        .din(new_Jinkela_wire_4744),
        .dout(new_Jinkela_wire_4745)
    );

    bfr new_Jinkela_buffer_1577 (
        .din(new_Jinkela_wire_1920),
        .dout(new_Jinkela_wire_1921)
    );

    bfr new_Jinkela_buffer_3998 (
        .din(new_Jinkela_wire_4694),
        .dout(new_Jinkela_wire_4695)
    );

    bfr new_Jinkela_buffer_3226 (
        .din(new_Jinkela_wire_3686),
        .dout(new_Jinkela_wire_3687)
    );

    bfr new_Jinkela_buffer_3173 (
        .din(new_Jinkela_wire_3627),
        .dout(new_Jinkela_wire_3628)
    );

    bfr new_Jinkela_buffer_1527 (
        .din(new_Jinkela_wire_1864),
        .dout(new_Jinkela_wire_1865)
    );

    bfr new_Jinkela_buffer_4938 (
        .din(new_Jinkela_wire_5887),
        .dout(new_Jinkela_wire_5888)
    );

    bfr new_Jinkela_buffer_4851 (
        .din(new_Jinkela_wire_5785),
        .dout(new_Jinkela_wire_5786)
    );

    bfr new_Jinkela_buffer_4085 (
        .din(new_Jinkela_wire_4785),
        .dout(new_Jinkela_wire_4786)
    );

    bfr new_Jinkela_buffer_1641 (
        .din(new_Jinkela_wire_1984),
        .dout(new_Jinkela_wire_1985)
    );

    bfr new_Jinkela_buffer_3999 (
        .din(new_Jinkela_wire_4695),
        .dout(new_Jinkela_wire_4696)
    );

    bfr new_Jinkela_buffer_3174 (
        .din(new_Jinkela_wire_3628),
        .dout(new_Jinkela_wire_3629)
    );

    bfr new_Jinkela_buffer_1528 (
        .din(new_Jinkela_wire_1865),
        .dout(new_Jinkela_wire_1866)
    );

    bfr new_Jinkela_buffer_4883 (
        .din(new_Jinkela_wire_5819),
        .dout(new_Jinkela_wire_5820)
    );

    bfr new_Jinkela_buffer_4852 (
        .din(new_Jinkela_wire_5786),
        .dout(new_Jinkela_wire_5787)
    );

    bfr new_Jinkela_buffer_4047 (
        .din(new_Jinkela_wire_4745),
        .dout(new_Jinkela_wire_4746)
    );

    spl2 new_Jinkela_splitter_161 (
        .a(new_Jinkela_wire_3702),
        .b(new_Jinkela_wire_3703),
        .c(new_Jinkela_wire_3704)
    );

    bfr new_Jinkela_buffer_1578 (
        .din(new_Jinkela_wire_1921),
        .dout(new_Jinkela_wire_1922)
    );

    bfr new_Jinkela_buffer_4000 (
        .din(new_Jinkela_wire_4696),
        .dout(new_Jinkela_wire_4697)
    );

    bfr new_Jinkela_buffer_3175 (
        .din(new_Jinkela_wire_3629),
        .dout(new_Jinkela_wire_3630)
    );

    bfr new_Jinkela_buffer_1529 (
        .din(new_Jinkela_wire_1866),
        .dout(new_Jinkela_wire_1867)
    );

    bfr new_Jinkela_buffer_4853 (
        .din(new_Jinkela_wire_5787),
        .dout(new_Jinkela_wire_5788)
    );

    bfr new_Jinkela_buffer_1650 (
        .din(N135),
        .dout(new_Jinkela_wire_1994)
    );

    bfr new_Jinkela_buffer_4001 (
        .din(new_Jinkela_wire_4697),
        .dout(new_Jinkela_wire_4698)
    );

    bfr new_Jinkela_buffer_3227 (
        .din(new_Jinkela_wire_3687),
        .dout(new_Jinkela_wire_3688)
    );

    bfr new_Jinkela_buffer_3176 (
        .din(new_Jinkela_wire_3630),
        .dout(new_Jinkela_wire_3631)
    );

    bfr new_Jinkela_buffer_1530 (
        .din(new_Jinkela_wire_1867),
        .dout(new_Jinkela_wire_1868)
    );

    bfr new_Jinkela_buffer_4884 (
        .din(new_Jinkela_wire_5820),
        .dout(new_Jinkela_wire_5821)
    );

    bfr new_Jinkela_buffer_4854 (
        .din(new_Jinkela_wire_5788),
        .dout(new_Jinkela_wire_5789)
    );

    bfr new_Jinkela_buffer_4048 (
        .din(new_Jinkela_wire_4746),
        .dout(new_Jinkela_wire_4747)
    );

    bfr new_Jinkela_buffer_1579 (
        .din(new_Jinkela_wire_1922),
        .dout(new_Jinkela_wire_1923)
    );

    bfr new_Jinkela_buffer_4002 (
        .din(new_Jinkela_wire_4698),
        .dout(new_Jinkela_wire_4699)
    );

    spl3L new_Jinkela_splitter_164 (
        .a(n_0064_),
        .d(new_Jinkela_wire_3719),
        .b(new_Jinkela_wire_3720),
        .c(new_Jinkela_wire_3721)
    );

    bfr new_Jinkela_buffer_3177 (
        .din(new_Jinkela_wire_3631),
        .dout(new_Jinkela_wire_3632)
    );

    bfr new_Jinkela_buffer_1531 (
        .din(new_Jinkela_wire_1868),
        .dout(new_Jinkela_wire_1869)
    );

    bfr new_Jinkela_buffer_4855 (
        .din(new_Jinkela_wire_5789),
        .dout(new_Jinkela_wire_5790)
    );

    bfr new_Jinkela_buffer_4086 (
        .din(new_Jinkela_wire_4786),
        .dout(new_Jinkela_wire_4787)
    );

    bfr new_Jinkela_buffer_1644 (
        .din(new_Jinkela_wire_1987),
        .dout(new_Jinkela_wire_1988)
    );

    bfr new_Jinkela_buffer_4885 (
        .din(new_Jinkela_wire_5821),
        .dout(new_Jinkela_wire_5822)
    );

    bfr new_Jinkela_buffer_4003 (
        .din(new_Jinkela_wire_4699),
        .dout(new_Jinkela_wire_4700)
    );

    bfr new_Jinkela_buffer_3228 (
        .din(new_Jinkela_wire_3688),
        .dout(new_Jinkela_wire_3689)
    );

    bfr new_Jinkela_buffer_3178 (
        .din(new_Jinkela_wire_3632),
        .dout(new_Jinkela_wire_3633)
    );

    bfr new_Jinkela_buffer_1532 (
        .din(new_Jinkela_wire_1869),
        .dout(new_Jinkela_wire_1870)
    );

    bfr new_Jinkela_buffer_4974 (
        .din(n_0205_),
        .dout(new_Jinkela_wire_5928)
    );

    bfr new_Jinkela_buffer_4856 (
        .din(new_Jinkela_wire_5790),
        .dout(new_Jinkela_wire_5791)
    );

    bfr new_Jinkela_buffer_4049 (
        .din(new_Jinkela_wire_4747),
        .dout(new_Jinkela_wire_4748)
    );

    bfr new_Jinkela_buffer_1580 (
        .din(new_Jinkela_wire_1923),
        .dout(new_Jinkela_wire_1924)
    );

    bfr new_Jinkela_buffer_4004 (
        .din(new_Jinkela_wire_4700),
        .dout(new_Jinkela_wire_4701)
    );

    bfr new_Jinkela_buffer_3238 (
        .din(new_Jinkela_wire_3706),
        .dout(new_Jinkela_wire_3707)
    );

    bfr new_Jinkela_buffer_3179 (
        .din(new_Jinkela_wire_3633),
        .dout(new_Jinkela_wire_3634)
    );

    bfr new_Jinkela_buffer_1533 (
        .din(new_Jinkela_wire_1870),
        .dout(new_Jinkela_wire_1871)
    );

    bfr new_Jinkela_buffer_4939 (
        .din(new_Jinkela_wire_5888),
        .dout(new_Jinkela_wire_5889)
    );

    bfr new_Jinkela_buffer_4857 (
        .din(new_Jinkela_wire_5791),
        .dout(new_Jinkela_wire_5792)
    );

    spl2 new_Jinkela_splitter_262 (
        .a(n_0298_),
        .b(new_Jinkela_wire_4858),
        .c(new_Jinkela_wire_4859)
    );

    bfr new_Jinkela_buffer_4119 (
        .din(new_Jinkela_wire_4819),
        .dout(new_Jinkela_wire_4820)
    );

    bfr new_Jinkela_buffer_1647 (
        .din(new_Jinkela_wire_1990),
        .dout(new_Jinkela_wire_1991)
    );

    bfr new_Jinkela_buffer_4005 (
        .din(new_Jinkela_wire_4701),
        .dout(new_Jinkela_wire_4702)
    );

    bfr new_Jinkela_buffer_3229 (
        .din(new_Jinkela_wire_3689),
        .dout(new_Jinkela_wire_3690)
    );

    bfr new_Jinkela_buffer_3180 (
        .din(new_Jinkela_wire_3634),
        .dout(new_Jinkela_wire_3635)
    );

    bfr new_Jinkela_buffer_1534 (
        .din(new_Jinkela_wire_1871),
        .dout(new_Jinkela_wire_1872)
    );

    bfr new_Jinkela_buffer_4886 (
        .din(new_Jinkela_wire_5822),
        .dout(new_Jinkela_wire_5823)
    );

    bfr new_Jinkela_buffer_4946 (
        .din(new_Jinkela_wire_5895),
        .dout(new_Jinkela_wire_5896)
    );

    bfr new_Jinkela_buffer_4858 (
        .din(new_Jinkela_wire_5792),
        .dout(new_Jinkela_wire_5793)
    );

    bfr new_Jinkela_buffer_4050 (
        .din(new_Jinkela_wire_4748),
        .dout(new_Jinkela_wire_4749)
    );

    bfr new_Jinkela_buffer_1581 (
        .din(new_Jinkela_wire_1924),
        .dout(new_Jinkela_wire_1925)
    );

    bfr new_Jinkela_buffer_4006 (
        .din(new_Jinkela_wire_4702),
        .dout(new_Jinkela_wire_4703)
    );

    bfr new_Jinkela_buffer_3239 (
        .din(new_Jinkela_wire_3707),
        .dout(new_Jinkela_wire_3708)
    );

    bfr new_Jinkela_buffer_3181 (
        .din(new_Jinkela_wire_3635),
        .dout(new_Jinkela_wire_3636)
    );

    bfr new_Jinkela_buffer_1535 (
        .din(new_Jinkela_wire_1872),
        .dout(new_Jinkela_wire_1873)
    );

    bfr new_Jinkela_buffer_4940 (
        .din(new_Jinkela_wire_5889),
        .dout(new_Jinkela_wire_5890)
    );

    bfr new_Jinkela_buffer_4859 (
        .din(new_Jinkela_wire_5793),
        .dout(new_Jinkela_wire_5794)
    );

    bfr new_Jinkela_buffer_4087 (
        .din(new_Jinkela_wire_4787),
        .dout(new_Jinkela_wire_4788)
    );

    bfr new_Jinkela_buffer_1645 (
        .din(new_Jinkela_wire_1988),
        .dout(new_Jinkela_wire_1989)
    );

    bfr new_Jinkela_buffer_4007 (
        .din(new_Jinkela_wire_4703),
        .dout(new_Jinkela_wire_4704)
    );

    bfr new_Jinkela_buffer_3230 (
        .din(new_Jinkela_wire_3690),
        .dout(new_Jinkela_wire_3691)
    );

    bfr new_Jinkela_buffer_3182 (
        .din(new_Jinkela_wire_3636),
        .dout(new_Jinkela_wire_3637)
    );

    bfr new_Jinkela_buffer_1536 (
        .din(new_Jinkela_wire_1873),
        .dout(new_Jinkela_wire_1874)
    );

    bfr new_Jinkela_buffer_4887 (
        .din(new_Jinkela_wire_5823),
        .dout(new_Jinkela_wire_5824)
    );

    bfr new_Jinkela_buffer_4860 (
        .din(new_Jinkela_wire_5794),
        .dout(new_Jinkela_wire_5795)
    );

    bfr new_Jinkela_buffer_4051 (
        .din(new_Jinkela_wire_4749),
        .dout(new_Jinkela_wire_4750)
    );

    bfr new_Jinkela_buffer_1582 (
        .din(new_Jinkela_wire_1925),
        .dout(new_Jinkela_wire_1926)
    );

    bfr new_Jinkela_buffer_4008 (
        .din(new_Jinkela_wire_4704),
        .dout(new_Jinkela_wire_4705)
    );

    bfr new_Jinkela_buffer_3183 (
        .din(new_Jinkela_wire_3637),
        .dout(new_Jinkela_wire_3638)
    );

    bfr new_Jinkela_buffer_1537 (
        .din(new_Jinkela_wire_1874),
        .dout(new_Jinkela_wire_1875)
    );

    bfr new_Jinkela_buffer_1719 (
        .din(N32),
        .dout(new_Jinkela_wire_2065)
    );

    bfr new_Jinkela_buffer_1654 (
        .din(N248),
        .dout(new_Jinkela_wire_1998)
    );

    bfr new_Jinkela_buffer_3243 (
        .din(n_0573_),
        .dout(new_Jinkela_wire_3718)
    );

    bfr new_Jinkela_buffer_4861 (
        .din(new_Jinkela_wire_5795),
        .dout(new_Jinkela_wire_5796)
    );

    bfr new_Jinkela_buffer_4009 (
        .din(new_Jinkela_wire_4705),
        .dout(new_Jinkela_wire_4706)
    );

    bfr new_Jinkela_buffer_3231 (
        .din(new_Jinkela_wire_3691),
        .dout(new_Jinkela_wire_3692)
    );

    bfr new_Jinkela_buffer_3184 (
        .din(new_Jinkela_wire_3638),
        .dout(new_Jinkela_wire_3639)
    );

    bfr new_Jinkela_buffer_1538 (
        .din(new_Jinkela_wire_1875),
        .dout(new_Jinkela_wire_1876)
    );

    bfr new_Jinkela_buffer_4888 (
        .din(new_Jinkela_wire_5824),
        .dout(new_Jinkela_wire_5825)
    );

    bfr new_Jinkela_buffer_4862 (
        .din(new_Jinkela_wire_5796),
        .dout(new_Jinkela_wire_5797)
    );

    bfr new_Jinkela_buffer_4052 (
        .din(new_Jinkela_wire_4750),
        .dout(new_Jinkela_wire_4751)
    );

    bfr new_Jinkela_buffer_1583 (
        .din(new_Jinkela_wire_1926),
        .dout(new_Jinkela_wire_1927)
    );

    bfr new_Jinkela_buffer_4010 (
        .din(new_Jinkela_wire_4706),
        .dout(new_Jinkela_wire_4707)
    );

    bfr new_Jinkela_buffer_3240 (
        .din(new_Jinkela_wire_3708),
        .dout(new_Jinkela_wire_3709)
    );

    bfr new_Jinkela_buffer_3185 (
        .din(new_Jinkela_wire_3639),
        .dout(new_Jinkela_wire_3640)
    );

    bfr new_Jinkela_buffer_1539 (
        .din(new_Jinkela_wire_1876),
        .dout(new_Jinkela_wire_1877)
    );

    bfr new_Jinkela_buffer_4941 (
        .din(new_Jinkela_wire_5890),
        .dout(new_Jinkela_wire_5891)
    );

    bfr new_Jinkela_buffer_4863 (
        .din(new_Jinkela_wire_5797),
        .dout(new_Jinkela_wire_5798)
    );

    bfr new_Jinkela_buffer_4088 (
        .din(new_Jinkela_wire_4788),
        .dout(new_Jinkela_wire_4789)
    );

    bfr new_Jinkela_buffer_1648 (
        .din(new_Jinkela_wire_1991),
        .dout(new_Jinkela_wire_1992)
    );

    bfr new_Jinkela_buffer_4011 (
        .din(new_Jinkela_wire_4707),
        .dout(new_Jinkela_wire_4708)
    );

    bfr new_Jinkela_buffer_3232 (
        .din(new_Jinkela_wire_3692),
        .dout(new_Jinkela_wire_3693)
    );

    bfr new_Jinkela_buffer_3186 (
        .din(new_Jinkela_wire_3640),
        .dout(new_Jinkela_wire_3641)
    );

    bfr new_Jinkela_buffer_1540 (
        .din(new_Jinkela_wire_1877),
        .dout(new_Jinkela_wire_1878)
    );

    bfr new_Jinkela_buffer_4889 (
        .din(new_Jinkela_wire_5825),
        .dout(new_Jinkela_wire_5826)
    );

    bfr new_Jinkela_buffer_4864 (
        .din(new_Jinkela_wire_5798),
        .dout(new_Jinkela_wire_5799)
    );

    bfr new_Jinkela_buffer_4053 (
        .din(new_Jinkela_wire_4751),
        .dout(new_Jinkela_wire_4752)
    );

    bfr new_Jinkela_buffer_1584 (
        .din(new_Jinkela_wire_1927),
        .dout(new_Jinkela_wire_1928)
    );

    bfr new_Jinkela_buffer_4012 (
        .din(new_Jinkela_wire_4708),
        .dout(new_Jinkela_wire_4709)
    );

    spl4L new_Jinkela_splitter_165 (
        .a(n_1158_),
        .d(new_Jinkela_wire_3722),
        .b(new_Jinkela_wire_3723),
        .e(new_Jinkela_wire_3724),
        .c(new_Jinkela_wire_3725)
    );

    bfr new_Jinkela_buffer_3187 (
        .din(new_Jinkela_wire_3641),
        .dout(new_Jinkela_wire_3642)
    );

    bfr new_Jinkela_buffer_1541 (
        .din(new_Jinkela_wire_1878),
        .dout(new_Jinkela_wire_1879)
    );

    bfr new_Jinkela_buffer_4865 (
        .din(new_Jinkela_wire_5799),
        .dout(new_Jinkela_wire_5800)
    );

    spl2 new_Jinkela_splitter_263 (
        .a(n_0207_),
        .b(new_Jinkela_wire_4860),
        .c(new_Jinkela_wire_4861)
    );

    bfr new_Jinkela_buffer_4120 (
        .din(new_Jinkela_wire_4820),
        .dout(new_Jinkela_wire_4821)
    );

    bfr new_Jinkela_buffer_1651 (
        .din(new_Jinkela_wire_1994),
        .dout(new_Jinkela_wire_1995)
    );

    bfr new_Jinkela_buffer_4947 (
        .din(new_Jinkela_wire_5896),
        .dout(new_Jinkela_wire_5897)
    );

    bfr new_Jinkela_buffer_4013 (
        .din(new_Jinkela_wire_4709),
        .dout(new_Jinkela_wire_4710)
    );

    bfr new_Jinkela_buffer_3241 (
        .din(new_Jinkela_wire_3709),
        .dout(new_Jinkela_wire_3710)
    );

    bfr new_Jinkela_buffer_3188 (
        .din(new_Jinkela_wire_3642),
        .dout(new_Jinkela_wire_3643)
    );

    bfr new_Jinkela_buffer_1542 (
        .din(new_Jinkela_wire_1879),
        .dout(new_Jinkela_wire_1880)
    );

    bfr new_Jinkela_buffer_4890 (
        .din(new_Jinkela_wire_5826),
        .dout(new_Jinkela_wire_5827)
    );

    bfr new_Jinkela_buffer_5686 (
        .din(new_Jinkela_wire_6854),
        .dout(new_Jinkela_wire_6855)
    );

    bfr new_Jinkela_buffer_8436 (
        .din(new_Jinkela_wire_10601),
        .dout(new_Jinkela_wire_10602)
    );

    spl2 new_Jinkela_splitter_460 (
        .a(n_1051_),
        .b(new_Jinkela_wire_6927),
        .c(new_Jinkela_wire_6928)
    );

    bfr new_Jinkela_buffer_5731 (
        .din(new_Jinkela_wire_6907),
        .dout(new_Jinkela_wire_6908)
    );

    bfr new_Jinkela_buffer_5687 (
        .din(new_Jinkela_wire_6855),
        .dout(new_Jinkela_wire_6856)
    );

    bfr new_Jinkela_buffer_8437 (
        .din(new_Jinkela_wire_10602),
        .dout(new_Jinkela_wire_10603)
    );

    bfr new_Jinkela_buffer_5722 (
        .din(new_Jinkela_wire_6896),
        .dout(new_Jinkela_wire_6897)
    );

    bfr new_Jinkela_buffer_5688 (
        .din(new_Jinkela_wire_6856),
        .dout(new_Jinkela_wire_6857)
    );

    bfr new_Jinkela_buffer_8438 (
        .din(new_Jinkela_wire_10603),
        .dout(new_Jinkela_wire_10604)
    );

    bfr new_Jinkela_buffer_5689 (
        .din(new_Jinkela_wire_6857),
        .dout(new_Jinkela_wire_6858)
    );

    bfr new_Jinkela_buffer_8439 (
        .din(new_Jinkela_wire_10604),
        .dout(new_Jinkela_wire_10605)
    );

    bfr new_Jinkela_buffer_5723 (
        .din(new_Jinkela_wire_6897),
        .dout(new_Jinkela_wire_6898)
    );

    bfr new_Jinkela_buffer_5690 (
        .din(new_Jinkela_wire_6858),
        .dout(new_Jinkela_wire_6859)
    );

    bfr new_Jinkela_buffer_8440 (
        .din(new_Jinkela_wire_10605),
        .dout(new_Jinkela_wire_10606)
    );

    spl2 new_Jinkela_splitter_461 (
        .a(n_0046_),
        .b(new_Jinkela_wire_6929),
        .c(new_Jinkela_wire_6930)
    );

    bfr new_Jinkela_buffer_5727 (
        .din(new_Jinkela_wire_6903),
        .dout(new_Jinkela_wire_6904)
    );

    bfr new_Jinkela_buffer_5691 (
        .din(new_Jinkela_wire_6859),
        .dout(new_Jinkela_wire_6860)
    );

    bfr new_Jinkela_buffer_8441 (
        .din(new_Jinkela_wire_10606),
        .dout(new_Jinkela_wire_10607)
    );

    bfr new_Jinkela_buffer_5724 (
        .din(new_Jinkela_wire_6898),
        .dout(new_Jinkela_wire_6899)
    );

    bfr new_Jinkela_buffer_5692 (
        .din(new_Jinkela_wire_6860),
        .dout(new_Jinkela_wire_6861)
    );

    bfr new_Jinkela_buffer_8442 (
        .din(new_Jinkela_wire_10607),
        .dout(new_Jinkela_wire_10608)
    );

    spl3L new_Jinkela_splitter_462 (
        .a(n_0723_),
        .d(new_Jinkela_wire_6940),
        .b(new_Jinkela_wire_6941),
        .c(new_Jinkela_wire_6942)
    );

    bfr new_Jinkela_buffer_5693 (
        .din(new_Jinkela_wire_6861),
        .dout(new_Jinkela_wire_6862)
    );

    bfr new_Jinkela_buffer_8443 (
        .din(new_Jinkela_wire_10608),
        .dout(new_Jinkela_wire_10609)
    );

    spl2 new_Jinkela_splitter_457 (
        .a(new_Jinkela_wire_6899),
        .b(new_Jinkela_wire_6900),
        .c(new_Jinkela_wire_6901)
    );

    bfr new_Jinkela_buffer_5694 (
        .din(new_Jinkela_wire_6862),
        .dout(new_Jinkela_wire_6863)
    );

    bfr new_Jinkela_buffer_8444 (
        .din(new_Jinkela_wire_10609),
        .dout(new_Jinkela_wire_10610)
    );

    bfr new_Jinkela_buffer_5695 (
        .din(new_Jinkela_wire_6863),
        .dout(new_Jinkela_wire_6864)
    );

    bfr new_Jinkela_buffer_8445 (
        .din(new_Jinkela_wire_10610),
        .dout(new_Jinkela_wire_10611)
    );

    bfr new_Jinkela_buffer_5746 (
        .din(new_Jinkela_wire_6930),
        .dout(new_Jinkela_wire_6931)
    );

    bfr new_Jinkela_buffer_5728 (
        .din(new_Jinkela_wire_6904),
        .dout(new_Jinkela_wire_6905)
    );

    bfr new_Jinkela_buffer_5696 (
        .din(new_Jinkela_wire_6864),
        .dout(new_Jinkela_wire_6865)
    );

    bfr new_Jinkela_buffer_8446 (
        .din(new_Jinkela_wire_10611),
        .dout(new_Jinkela_wire_10612)
    );

    bfr new_Jinkela_buffer_5755 (
        .din(n_0590_),
        .dout(new_Jinkela_wire_6943)
    );

    bfr new_Jinkela_buffer_5729 (
        .din(new_Jinkela_wire_6905),
        .dout(new_Jinkela_wire_6906)
    );

    bfr new_Jinkela_buffer_5697 (
        .din(new_Jinkela_wire_6865),
        .dout(new_Jinkela_wire_6866)
    );

    bfr new_Jinkela_buffer_8447 (
        .din(new_Jinkela_wire_10612),
        .dout(new_Jinkela_wire_10613)
    );

    spl4L new_Jinkela_splitter_464 (
        .a(n_0162_),
        .d(new_Jinkela_wire_6947),
        .b(new_Jinkela_wire_6948),
        .e(new_Jinkela_wire_6949),
        .c(new_Jinkela_wire_6950)
    );

    bfr new_Jinkela_buffer_5698 (
        .din(new_Jinkela_wire_6866),
        .dout(new_Jinkela_wire_6867)
    );

    bfr new_Jinkela_buffer_8448 (
        .din(new_Jinkela_wire_10613),
        .dout(new_Jinkela_wire_10614)
    );

    bfr new_Jinkela_buffer_5756 (
        .din(new_Jinkela_wire_6943),
        .dout(new_Jinkela_wire_6944)
    );

    bfr new_Jinkela_buffer_5730 (
        .din(new_Jinkela_wire_6906),
        .dout(new_Jinkela_wire_6907)
    );

    bfr new_Jinkela_buffer_5699 (
        .din(new_Jinkela_wire_6867),
        .dout(new_Jinkela_wire_6868)
    );

    bfr new_Jinkela_buffer_8449 (
        .din(new_Jinkela_wire_10614),
        .dout(new_Jinkela_wire_10615)
    );

    bfr new_Jinkela_buffer_5817 (
        .din(n_0526_),
        .dout(new_Jinkela_wire_7011)
    );

    bfr new_Jinkela_buffer_5700 (
        .din(new_Jinkela_wire_6868),
        .dout(new_Jinkela_wire_6869)
    );

    bfr new_Jinkela_buffer_8450 (
        .din(new_Jinkela_wire_10615),
        .dout(new_Jinkela_wire_10616)
    );

    bfr new_Jinkela_buffer_5747 (
        .din(new_Jinkela_wire_6931),
        .dout(new_Jinkela_wire_6932)
    );

    bfr new_Jinkela_buffer_5732 (
        .din(new_Jinkela_wire_6908),
        .dout(new_Jinkela_wire_6909)
    );

    bfr new_Jinkela_buffer_5701 (
        .din(new_Jinkela_wire_6869),
        .dout(new_Jinkela_wire_6870)
    );

    bfr new_Jinkela_buffer_8451 (
        .din(new_Jinkela_wire_10616),
        .dout(new_Jinkela_wire_10617)
    );

    bfr new_Jinkela_buffer_5702 (
        .din(new_Jinkela_wire_6870),
        .dout(new_Jinkela_wire_6871)
    );

    bfr new_Jinkela_buffer_8452 (
        .din(new_Jinkela_wire_10617),
        .dout(new_Jinkela_wire_10618)
    );

    bfr new_Jinkela_buffer_5703 (
        .din(new_Jinkela_wire_6871),
        .dout(new_Jinkela_wire_6872)
    );

    bfr new_Jinkela_buffer_8453 (
        .din(new_Jinkela_wire_10618),
        .dout(new_Jinkela_wire_10619)
    );

    bfr new_Jinkela_buffer_5704 (
        .din(new_Jinkela_wire_6872),
        .dout(new_Jinkela_wire_6873)
    );

    bfr new_Jinkela_buffer_8454 (
        .din(new_Jinkela_wire_10619),
        .dout(new_Jinkela_wire_10620)
    );

    bfr new_Jinkela_buffer_5748 (
        .din(new_Jinkela_wire_6932),
        .dout(new_Jinkela_wire_6933)
    );

    bfr new_Jinkela_buffer_5733 (
        .din(new_Jinkela_wire_6909),
        .dout(new_Jinkela_wire_6910)
    );

    bfr new_Jinkela_buffer_5705 (
        .din(new_Jinkela_wire_6873),
        .dout(new_Jinkela_wire_6874)
    );

    bfr new_Jinkela_buffer_8455 (
        .din(new_Jinkela_wire_10620),
        .dout(new_Jinkela_wire_10621)
    );

    bfr new_Jinkela_buffer_5706 (
        .din(new_Jinkela_wire_6874),
        .dout(new_Jinkela_wire_6875)
    );

    bfr new_Jinkela_buffer_8456 (
        .din(new_Jinkela_wire_10621),
        .dout(new_Jinkela_wire_10622)
    );

    bfr new_Jinkela_buffer_989 (
        .din(new_Jinkela_wire_1063),
        .dout(new_Jinkela_wire_1064)
    );

    bfr new_Jinkela_buffer_1634 (
        .din(N203),
        .dout(new_Jinkela_wire_1978)
    );

    bfr new_Jinkela_buffer_1502 (
        .din(new_Jinkela_wire_1836),
        .dout(new_Jinkela_wire_1837)
    );

    spl2 new_Jinkela_splitter_94 (
        .a(new_Jinkela_wire_1405),
        .b(new_Jinkela_wire_1406),
        .c(new_Jinkela_wire_1407)
    );

    bfr new_Jinkela_buffer_7459 (
        .din(new_Jinkela_wire_9273),
        .dout(new_Jinkela_wire_9274)
    );

    bfr new_Jinkela_buffer_990 (
        .din(new_Jinkela_wire_1064),
        .dout(new_Jinkela_wire_1065)
    );

    bfr new_Jinkela_buffer_1565 (
        .din(new_Jinkela_wire_1902),
        .dout(new_Jinkela_wire_1903)
    );

    bfr new_Jinkela_buffer_7460 (
        .din(new_Jinkela_wire_9274),
        .dout(new_Jinkela_wire_9275)
    );

    bfr new_Jinkela_buffer_1503 (
        .din(new_Jinkela_wire_1837),
        .dout(new_Jinkela_wire_1838)
    );

    bfr new_Jinkela_buffer_1039 (
        .din(new_Jinkela_wire_1115),
        .dout(new_Jinkela_wire_1116)
    );

    bfr new_Jinkela_buffer_7484 (
        .din(new_Jinkela_wire_9310),
        .dout(new_Jinkela_wire_9311)
    );

    bfr new_Jinkela_buffer_991 (
        .din(new_Jinkela_wire_1065),
        .dout(new_Jinkela_wire_1066)
    );

    bfr new_Jinkela_buffer_1566 (
        .din(new_Jinkela_wire_1907),
        .dout(new_Jinkela_wire_1908)
    );

    bfr new_Jinkela_buffer_1631 (
        .din(new_Jinkela_wire_1974),
        .dout(new_Jinkela_wire_1975)
    );

    bfr new_Jinkela_buffer_7461 (
        .din(new_Jinkela_wire_9275),
        .dout(new_Jinkela_wire_9276)
    );

    spl3L new_Jinkela_splitter_106 (
        .a(new_Jinkela_wire_1838),
        .d(new_Jinkela_wire_1839),
        .b(new_Jinkela_wire_1840),
        .c(new_Jinkela_wire_1841)
    );

    spl2 new_Jinkela_splitter_738 (
        .a(new_Jinkela_wire_9346),
        .b(new_Jinkela_wire_9347),
        .c(new_Jinkela_wire_9348)
    );

    bfr new_Jinkela_buffer_992 (
        .din(new_Jinkela_wire_1066),
        .dout(new_Jinkela_wire_1067)
    );

    bfr new_Jinkela_buffer_7526 (
        .din(new_Jinkela_wire_9367),
        .dout(new_Jinkela_wire_9368)
    );

    bfr new_Jinkela_buffer_7462 (
        .din(new_Jinkela_wire_9276),
        .dout(new_Jinkela_wire_9277)
    );

    bfr new_Jinkela_buffer_1099 (
        .din(new_Jinkela_wire_1407),
        .dout(new_Jinkela_wire_1408)
    );

    bfr new_Jinkela_buffer_1504 (
        .din(new_Jinkela_wire_1841),
        .dout(new_Jinkela_wire_1842)
    );

    bfr new_Jinkela_buffer_1040 (
        .din(new_Jinkela_wire_1116),
        .dout(new_Jinkela_wire_1117)
    );

    bfr new_Jinkela_buffer_7485 (
        .din(new_Jinkela_wire_9311),
        .dout(new_Jinkela_wire_9312)
    );

    bfr new_Jinkela_buffer_993 (
        .din(new_Jinkela_wire_1067),
        .dout(new_Jinkela_wire_1068)
    );

    spl2 new_Jinkela_splitter_108 (
        .a(new_Jinkela_wire_1908),
        .b(new_Jinkela_wire_1909),
        .c(new_Jinkela_wire_1910)
    );

    bfr new_Jinkela_buffer_7463 (
        .din(new_Jinkela_wire_9277),
        .dout(new_Jinkela_wire_9278)
    );

    bfr new_Jinkela_buffer_1505 (
        .din(new_Jinkela_wire_1842),
        .dout(new_Jinkela_wire_1843)
    );

    bfr new_Jinkela_buffer_1289 (
        .din(N239),
        .dout(new_Jinkela_wire_1610)
    );

    bfr new_Jinkela_buffer_994 (
        .din(new_Jinkela_wire_1068),
        .dout(new_Jinkela_wire_1069)
    );

    bfr new_Jinkela_buffer_1567 (
        .din(new_Jinkela_wire_1910),
        .dout(new_Jinkela_wire_1911)
    );

    bfr new_Jinkela_buffer_7464 (
        .din(new_Jinkela_wire_9278),
        .dout(new_Jinkela_wire_9279)
    );

    spl2 new_Jinkela_splitter_96 (
        .a(new_Jinkela_wire_1474),
        .b(new_Jinkela_wire_1475),
        .c(new_Jinkela_wire_1476)
    );

    bfr new_Jinkela_buffer_1506 (
        .din(new_Jinkela_wire_1843),
        .dout(new_Jinkela_wire_1844)
    );

    bfr new_Jinkela_buffer_1041 (
        .din(new_Jinkela_wire_1117),
        .dout(new_Jinkela_wire_1118)
    );

    bfr new_Jinkela_buffer_7486 (
        .din(new_Jinkela_wire_9312),
        .dout(new_Jinkela_wire_9313)
    );

    bfr new_Jinkela_buffer_995 (
        .din(new_Jinkela_wire_1069),
        .dout(new_Jinkela_wire_1070)
    );

    bfr new_Jinkela_buffer_1638 (
        .din(N206),
        .dout(new_Jinkela_wire_1982)
    );

    bfr new_Jinkela_buffer_7465 (
        .din(new_Jinkela_wire_9279),
        .dout(new_Jinkela_wire_9280)
    );

    bfr new_Jinkela_buffer_1507 (
        .din(new_Jinkela_wire_1844),
        .dout(new_Jinkela_wire_1845)
    );

    bfr new_Jinkela_buffer_7511 (
        .din(new_Jinkela_wire_9348),
        .dout(new_Jinkela_wire_9349)
    );

    bfr new_Jinkela_buffer_996 (
        .din(new_Jinkela_wire_1070),
        .dout(new_Jinkela_wire_1071)
    );

    bfr new_Jinkela_buffer_1632 (
        .din(new_Jinkela_wire_1975),
        .dout(new_Jinkela_wire_1976)
    );

    bfr new_Jinkela_buffer_7528 (
        .din(n_0181_),
        .dout(new_Jinkela_wire_9370)
    );

    bfr new_Jinkela_buffer_7466 (
        .din(new_Jinkela_wire_9280),
        .dout(new_Jinkela_wire_9281)
    );

    bfr new_Jinkela_buffer_1100 (
        .din(new_Jinkela_wire_1408),
        .dout(new_Jinkela_wire_1409)
    );

    bfr new_Jinkela_buffer_1508 (
        .din(new_Jinkela_wire_1845),
        .dout(new_Jinkela_wire_1846)
    );

    bfr new_Jinkela_buffer_1042 (
        .din(new_Jinkela_wire_1118),
        .dout(new_Jinkela_wire_1119)
    );

    bfr new_Jinkela_buffer_7487 (
        .din(new_Jinkela_wire_9313),
        .dout(new_Jinkela_wire_9314)
    );

    bfr new_Jinkela_buffer_997 (
        .din(new_Jinkela_wire_1071),
        .dout(new_Jinkela_wire_1072)
    );

    bfr new_Jinkela_buffer_1568 (
        .din(new_Jinkela_wire_1911),
        .dout(new_Jinkela_wire_1912)
    );

    bfr new_Jinkela_buffer_7467 (
        .din(new_Jinkela_wire_9281),
        .dout(new_Jinkela_wire_9282)
    );

    bfr new_Jinkela_buffer_1509 (
        .din(new_Jinkela_wire_1846),
        .dout(new_Jinkela_wire_1847)
    );

    bfr new_Jinkela_buffer_998 (
        .din(new_Jinkela_wire_1072),
        .dout(new_Jinkela_wire_1073)
    );

    bfr new_Jinkela_buffer_1635 (
        .din(new_Jinkela_wire_1978),
        .dout(new_Jinkela_wire_1979)
    );

    spl2 new_Jinkela_splitter_741 (
        .a(n_0351_),
        .b(new_Jinkela_wire_9375),
        .c(new_Jinkela_wire_9376)
    );

    bfr new_Jinkela_buffer_7468 (
        .din(new_Jinkela_wire_9282),
        .dout(new_Jinkela_wire_9283)
    );

    bfr new_Jinkela_buffer_1162 (
        .din(new_Jinkela_wire_1473),
        .dout(new_Jinkela_wire_1474)
    );

    bfr new_Jinkela_buffer_1510 (
        .din(new_Jinkela_wire_1847),
        .dout(new_Jinkela_wire_1848)
    );

    bfr new_Jinkela_buffer_1043 (
        .din(new_Jinkela_wire_1119),
        .dout(new_Jinkela_wire_1120)
    );

    bfr new_Jinkela_buffer_7488 (
        .din(new_Jinkela_wire_9314),
        .dout(new_Jinkela_wire_9315)
    );

    bfr new_Jinkela_buffer_999 (
        .din(new_Jinkela_wire_1073),
        .dout(new_Jinkela_wire_1074)
    );

    bfr new_Jinkela_buffer_1569 (
        .din(new_Jinkela_wire_1912),
        .dout(new_Jinkela_wire_1913)
    );

    bfr new_Jinkela_buffer_7469 (
        .din(new_Jinkela_wire_9283),
        .dout(new_Jinkela_wire_9284)
    );

    bfr new_Jinkela_buffer_1511 (
        .din(new_Jinkela_wire_1848),
        .dout(new_Jinkela_wire_1849)
    );

    bfr new_Jinkela_buffer_1000 (
        .din(new_Jinkela_wire_1074),
        .dout(new_Jinkela_wire_1075)
    );

    bfr new_Jinkela_buffer_1633 (
        .din(new_Jinkela_wire_1976),
        .dout(new_Jinkela_wire_1977)
    );

    bfr new_Jinkela_buffer_7533 (
        .din(n_0184_),
        .dout(new_Jinkela_wire_9377)
    );

    bfr new_Jinkela_buffer_7470 (
        .din(new_Jinkela_wire_9284),
        .dout(new_Jinkela_wire_9285)
    );

    bfr new_Jinkela_buffer_1512 (
        .din(new_Jinkela_wire_1849),
        .dout(new_Jinkela_wire_1850)
    );

    bfr new_Jinkela_buffer_1044 (
        .din(new_Jinkela_wire_1120),
        .dout(new_Jinkela_wire_1121)
    );

    bfr new_Jinkela_buffer_7489 (
        .din(new_Jinkela_wire_9315),
        .dout(new_Jinkela_wire_9316)
    );

    bfr new_Jinkela_buffer_1001 (
        .din(new_Jinkela_wire_1075),
        .dout(new_Jinkela_wire_1076)
    );

    bfr new_Jinkela_buffer_1570 (
        .din(new_Jinkela_wire_1913),
        .dout(new_Jinkela_wire_1914)
    );

    bfr new_Jinkela_buffer_7471 (
        .din(new_Jinkela_wire_9285),
        .dout(new_Jinkela_wire_9286)
    );

    bfr new_Jinkela_buffer_1513 (
        .din(new_Jinkela_wire_1850),
        .dout(new_Jinkela_wire_1851)
    );

    bfr new_Jinkela_buffer_7529 (
        .din(new_Jinkela_wire_9370),
        .dout(new_Jinkela_wire_9371)
    );

    bfr new_Jinkela_buffer_1002 (
        .din(new_Jinkela_wire_1076),
        .dout(new_Jinkela_wire_1077)
    );

    bfr new_Jinkela_buffer_1642 (
        .din(N76),
        .dout(new_Jinkela_wire_1986)
    );

    bfr new_Jinkela_buffer_7512 (
        .din(new_Jinkela_wire_9349),
        .dout(new_Jinkela_wire_9350)
    );

    bfr new_Jinkela_buffer_7472 (
        .din(new_Jinkela_wire_9286),
        .dout(new_Jinkela_wire_9287)
    );

    bfr new_Jinkela_buffer_1514 (
        .din(new_Jinkela_wire_1851),
        .dout(new_Jinkela_wire_1852)
    );

    bfr new_Jinkela_buffer_1045 (
        .din(new_Jinkela_wire_1121),
        .dout(new_Jinkela_wire_1122)
    );

    bfr new_Jinkela_buffer_7490 (
        .din(new_Jinkela_wire_9316),
        .dout(new_Jinkela_wire_9317)
    );

    bfr new_Jinkela_buffer_1003 (
        .din(new_Jinkela_wire_1077),
        .dout(new_Jinkela_wire_1078)
    );

    bfr new_Jinkela_buffer_1571 (
        .din(new_Jinkela_wire_1914),
        .dout(new_Jinkela_wire_1915)
    );

    bfr new_Jinkela_buffer_7473 (
        .din(new_Jinkela_wire_9287),
        .dout(new_Jinkela_wire_9288)
    );

    bfr new_Jinkela_buffer_1515 (
        .din(new_Jinkela_wire_1852),
        .dout(new_Jinkela_wire_1853)
    );

    bfr new_Jinkela_buffer_1101 (
        .din(new_Jinkela_wire_1409),
        .dout(new_Jinkela_wire_1410)
    );

    bfr new_Jinkela_buffer_1004 (
        .din(new_Jinkela_wire_1078),
        .dout(new_Jinkela_wire_1079)
    );

    bfr new_Jinkela_buffer_1636 (
        .din(new_Jinkela_wire_1979),
        .dout(new_Jinkela_wire_1980)
    );

    bfr new_Jinkela_buffer_7527 (
        .din(new_Jinkela_wire_9368),
        .dout(new_Jinkela_wire_9369)
    );

    spl2 new_Jinkela_splitter_728 (
        .a(new_Jinkela_wire_9288),
        .b(new_Jinkela_wire_9289),
        .c(new_Jinkela_wire_9290)
    );

    bfr new_Jinkela_buffer_1516 (
        .din(new_Jinkela_wire_1853),
        .dout(new_Jinkela_wire_1854)
    );

    bfr new_Jinkela_buffer_1046 (
        .din(new_Jinkela_wire_1122),
        .dout(new_Jinkela_wire_1123)
    );

    bfr new_Jinkela_buffer_1005 (
        .din(new_Jinkela_wire_1079),
        .dout(new_Jinkela_wire_1080)
    );

    bfr new_Jinkela_buffer_1572 (
        .din(new_Jinkela_wire_1915),
        .dout(new_Jinkela_wire_1916)
    );

    spl2 new_Jinkela_splitter_739 (
        .a(new_Jinkela_wire_9350),
        .b(new_Jinkela_wire_9351),
        .c(new_Jinkela_wire_9352)
    );

    bfr new_Jinkela_buffer_7491 (
        .din(new_Jinkela_wire_9317),
        .dout(new_Jinkela_wire_9318)
    );

    bfr new_Jinkela_buffer_1517 (
        .din(new_Jinkela_wire_1854),
        .dout(new_Jinkela_wire_1855)
    );

    spl3L new_Jinkela_splitter_95 (
        .a(new_Jinkela_wire_1410),
        .d(new_Jinkela_wire_1411),
        .b(new_Jinkela_wire_1412),
        .c(new_Jinkela_wire_1413)
    );

    bfr new_Jinkela_buffer_7492 (
        .din(new_Jinkela_wire_9318),
        .dout(new_Jinkela_wire_9319)
    );

    bfr new_Jinkela_buffer_1006 (
        .din(new_Jinkela_wire_1080),
        .dout(new_Jinkela_wire_1081)
    );

    bfr new_Jinkela_buffer_1639 (
        .din(new_Jinkela_wire_1982),
        .dout(new_Jinkela_wire_1983)
    );

    bfr new_Jinkela_buffer_1518 (
        .din(new_Jinkela_wire_1855),
        .dout(new_Jinkela_wire_1856)
    );

    bfr new_Jinkela_buffer_7513 (
        .din(new_Jinkela_wire_9352),
        .dout(new_Jinkela_wire_9353)
    );

    bfr new_Jinkela_buffer_1047 (
        .din(new_Jinkela_wire_1123),
        .dout(new_Jinkela_wire_1124)
    );

    bfr new_Jinkela_buffer_7493 (
        .din(new_Jinkela_wire_9319),
        .dout(new_Jinkela_wire_9320)
    );

    bfr new_Jinkela_buffer_1007 (
        .din(new_Jinkela_wire_1081),
        .dout(new_Jinkela_wire_1082)
    );

    bfr new_Jinkela_buffer_1573 (
        .din(new_Jinkela_wire_1916),
        .dout(new_Jinkela_wire_1917)
    );

    bfr new_Jinkela_buffer_1519 (
        .din(new_Jinkela_wire_1856),
        .dout(new_Jinkela_wire_1857)
    );

    bfr new_Jinkela_buffer_1163 (
        .din(new_Jinkela_wire_1476),
        .dout(new_Jinkela_wire_1477)
    );

    bfr new_Jinkela_buffer_7494 (
        .din(new_Jinkela_wire_9320),
        .dout(new_Jinkela_wire_9321)
    );

    bfr new_Jinkela_buffer_1008 (
        .din(new_Jinkela_wire_1082),
        .dout(new_Jinkela_wire_1083)
    );

    bfr new_Jinkela_buffer_1637 (
        .din(new_Jinkela_wire_1980),
        .dout(new_Jinkela_wire_1981)
    );

    bfr new_Jinkela_buffer_1520 (
        .din(new_Jinkela_wire_1857),
        .dout(new_Jinkela_wire_1858)
    );

    bfr new_Jinkela_buffer_1048 (
        .din(new_Jinkela_wire_1124),
        .dout(new_Jinkela_wire_1125)
    );

    bfr new_Jinkela_buffer_7495 (
        .din(new_Jinkela_wire_9321),
        .dout(new_Jinkela_wire_9322)
    );

    bfr new_Jinkela_buffer_1009 (
        .din(new_Jinkela_wire_1083),
        .dout(new_Jinkela_wire_1084)
    );

    bfr new_Jinkela_buffer_1574 (
        .din(new_Jinkela_wire_1917),
        .dout(new_Jinkela_wire_1918)
    );

    bfr new_Jinkela_buffer_7530 (
        .din(new_Jinkela_wire_9371),
        .dout(new_Jinkela_wire_9372)
    );

    bfr new_Jinkela_buffer_1521 (
        .din(new_Jinkela_wire_1858),
        .dout(new_Jinkela_wire_1859)
    );

    bfr new_Jinkela_buffer_7514 (
        .din(new_Jinkela_wire_9353),
        .dout(new_Jinkela_wire_9354)
    );

    bfr new_Jinkela_buffer_7496 (
        .din(new_Jinkela_wire_9322),
        .dout(new_Jinkela_wire_9323)
    );

    bfr new_Jinkela_buffer_4054 (
        .din(new_Jinkela_wire_4752),
        .dout(new_Jinkela_wire_4753)
    );

    bfr new_Jinkela_buffer_2301 (
        .din(new_Jinkela_wire_2692),
        .dout(new_Jinkela_wire_2693)
    );

    bfr new_Jinkela_buffer_4014 (
        .din(new_Jinkela_wire_4710),
        .dout(new_Jinkela_wire_4711)
    );

    bfr new_Jinkela_buffer_2265 (
        .din(new_Jinkela_wire_2651),
        .dout(new_Jinkela_wire_2652)
    );

    bfr new_Jinkela_buffer_4089 (
        .din(new_Jinkela_wire_4789),
        .dout(new_Jinkela_wire_4790)
    );

    bfr new_Jinkela_buffer_2418 (
        .din(new_Jinkela_wire_2814),
        .dout(new_Jinkela_wire_2815)
    );

    bfr new_Jinkela_buffer_4015 (
        .din(new_Jinkela_wire_4711),
        .dout(new_Jinkela_wire_4712)
    );

    bfr new_Jinkela_buffer_2266 (
        .din(new_Jinkela_wire_2652),
        .dout(new_Jinkela_wire_2653)
    );

    bfr new_Jinkela_buffer_4055 (
        .din(new_Jinkela_wire_4753),
        .dout(new_Jinkela_wire_4754)
    );

    bfr new_Jinkela_buffer_2302 (
        .din(new_Jinkela_wire_2693),
        .dout(new_Jinkela_wire_2694)
    );

    bfr new_Jinkela_buffer_4016 (
        .din(new_Jinkela_wire_4712),
        .dout(new_Jinkela_wire_4713)
    );

    bfr new_Jinkela_buffer_2267 (
        .din(new_Jinkela_wire_2653),
        .dout(new_Jinkela_wire_2654)
    );

    bfr new_Jinkela_buffer_2354 (
        .din(new_Jinkela_wire_2750),
        .dout(new_Jinkela_wire_2751)
    );

    bfr new_Jinkela_buffer_4017 (
        .din(new_Jinkela_wire_4713),
        .dout(new_Jinkela_wire_4714)
    );

    bfr new_Jinkela_buffer_2268 (
        .din(new_Jinkela_wire_2654),
        .dout(new_Jinkela_wire_2655)
    );

    bfr new_Jinkela_buffer_4056 (
        .din(new_Jinkela_wire_4754),
        .dout(new_Jinkela_wire_4755)
    );

    bfr new_Jinkela_buffer_2303 (
        .din(new_Jinkela_wire_2694),
        .dout(new_Jinkela_wire_2695)
    );

    bfr new_Jinkela_buffer_4018 (
        .din(new_Jinkela_wire_4714),
        .dout(new_Jinkela_wire_4715)
    );

    bfr new_Jinkela_buffer_2269 (
        .din(new_Jinkela_wire_2655),
        .dout(new_Jinkela_wire_2656)
    );

    bfr new_Jinkela_buffer_4090 (
        .din(new_Jinkela_wire_4790),
        .dout(new_Jinkela_wire_4791)
    );

    bfr new_Jinkela_buffer_2488 (
        .din(N58),
        .dout(new_Jinkela_wire_2890)
    );

    bfr new_Jinkela_buffer_4019 (
        .din(new_Jinkela_wire_4715),
        .dout(new_Jinkela_wire_4716)
    );

    bfr new_Jinkela_buffer_2270 (
        .din(new_Jinkela_wire_2656),
        .dout(new_Jinkela_wire_2657)
    );

    bfr new_Jinkela_buffer_4057 (
        .din(new_Jinkela_wire_4755),
        .dout(new_Jinkela_wire_4756)
    );

    bfr new_Jinkela_buffer_2304 (
        .din(new_Jinkela_wire_2695),
        .dout(new_Jinkela_wire_2696)
    );

    bfr new_Jinkela_buffer_4020 (
        .din(new_Jinkela_wire_4716),
        .dout(new_Jinkela_wire_4717)
    );

    bfr new_Jinkela_buffer_2271 (
        .din(new_Jinkela_wire_2657),
        .dout(new_Jinkela_wire_2658)
    );

    bfr new_Jinkela_buffer_2355 (
        .din(new_Jinkela_wire_2751),
        .dout(new_Jinkela_wire_2752)
    );

    bfr new_Jinkela_buffer_4121 (
        .din(new_Jinkela_wire_4821),
        .dout(new_Jinkela_wire_4822)
    );

    bfr new_Jinkela_buffer_4021 (
        .din(new_Jinkela_wire_4717),
        .dout(new_Jinkela_wire_4718)
    );

    bfr new_Jinkela_buffer_2305 (
        .din(new_Jinkela_wire_2696),
        .dout(new_Jinkela_wire_2697)
    );

    bfr new_Jinkela_buffer_4058 (
        .din(new_Jinkela_wire_4756),
        .dout(new_Jinkela_wire_4757)
    );

    bfr new_Jinkela_buffer_2419 (
        .din(new_Jinkela_wire_2815),
        .dout(new_Jinkela_wire_2816)
    );

    bfr new_Jinkela_buffer_4022 (
        .din(new_Jinkela_wire_4718),
        .dout(new_Jinkela_wire_4719)
    );

    bfr new_Jinkela_buffer_2306 (
        .din(new_Jinkela_wire_2697),
        .dout(new_Jinkela_wire_2698)
    );

    bfr new_Jinkela_buffer_4091 (
        .din(new_Jinkela_wire_4791),
        .dout(new_Jinkela_wire_4792)
    );

    bfr new_Jinkela_buffer_2356 (
        .din(new_Jinkela_wire_2752),
        .dout(new_Jinkela_wire_2753)
    );

    bfr new_Jinkela_buffer_4023 (
        .din(new_Jinkela_wire_4719),
        .dout(new_Jinkela_wire_4720)
    );

    bfr new_Jinkela_buffer_2307 (
        .din(new_Jinkela_wire_2698),
        .dout(new_Jinkela_wire_2699)
    );

    bfr new_Jinkela_buffer_4059 (
        .din(new_Jinkela_wire_4757),
        .dout(new_Jinkela_wire_4758)
    );

    bfr new_Jinkela_buffer_2492 (
        .din(N216),
        .dout(new_Jinkela_wire_2894)
    );

    bfr new_Jinkela_buffer_4024 (
        .din(new_Jinkela_wire_4720),
        .dout(new_Jinkela_wire_4721)
    );

    bfr new_Jinkela_buffer_2308 (
        .din(new_Jinkela_wire_2699),
        .dout(new_Jinkela_wire_2700)
    );

    bfr new_Jinkela_buffer_2357 (
        .din(new_Jinkela_wire_2753),
        .dout(new_Jinkela_wire_2754)
    );

    bfr new_Jinkela_buffer_4025 (
        .din(new_Jinkela_wire_4721),
        .dout(new_Jinkela_wire_4722)
    );

    bfr new_Jinkela_buffer_2309 (
        .din(new_Jinkela_wire_2700),
        .dout(new_Jinkela_wire_2701)
    );

    bfr new_Jinkela_buffer_4060 (
        .din(new_Jinkela_wire_4758),
        .dout(new_Jinkela_wire_4759)
    );

    bfr new_Jinkela_buffer_2422 (
        .din(new_Jinkela_wire_2818),
        .dout(new_Jinkela_wire_2819)
    );

    bfr new_Jinkela_buffer_2485 (
        .din(new_Jinkela_wire_2886),
        .dout(new_Jinkela_wire_2887)
    );

    bfr new_Jinkela_buffer_4026 (
        .din(new_Jinkela_wire_4722),
        .dout(new_Jinkela_wire_4723)
    );

    bfr new_Jinkela_buffer_2310 (
        .din(new_Jinkela_wire_2701),
        .dout(new_Jinkela_wire_2702)
    );

    bfr new_Jinkela_buffer_4092 (
        .din(new_Jinkela_wire_4792),
        .dout(new_Jinkela_wire_4793)
    );

    bfr new_Jinkela_buffer_2358 (
        .din(new_Jinkela_wire_2754),
        .dout(new_Jinkela_wire_2755)
    );

    bfr new_Jinkela_buffer_4027 (
        .din(new_Jinkela_wire_4723),
        .dout(new_Jinkela_wire_4724)
    );

    bfr new_Jinkela_buffer_2311 (
        .din(new_Jinkela_wire_2702),
        .dout(new_Jinkela_wire_2703)
    );

    bfr new_Jinkela_buffer_4061 (
        .din(new_Jinkela_wire_4759),
        .dout(new_Jinkela_wire_4760)
    );

    bfr new_Jinkela_buffer_2421 (
        .din(new_Jinkela_wire_2817),
        .dout(new_Jinkela_wire_2818)
    );

    bfr new_Jinkela_buffer_4028 (
        .din(new_Jinkela_wire_4724),
        .dout(new_Jinkela_wire_4725)
    );

    bfr new_Jinkela_buffer_2312 (
        .din(new_Jinkela_wire_2703),
        .dout(new_Jinkela_wire_2704)
    );

    spl2 new_Jinkela_splitter_264 (
        .a(n_0321_),
        .b(new_Jinkela_wire_4862),
        .c(new_Jinkela_wire_4863)
    );

    bfr new_Jinkela_buffer_2359 (
        .din(new_Jinkela_wire_2755),
        .dout(new_Jinkela_wire_2756)
    );

    bfr new_Jinkela_buffer_4122 (
        .din(new_Jinkela_wire_4822),
        .dout(new_Jinkela_wire_4823)
    );

    bfr new_Jinkela_buffer_4029 (
        .din(new_Jinkela_wire_4725),
        .dout(new_Jinkela_wire_4726)
    );

    bfr new_Jinkela_buffer_2313 (
        .din(new_Jinkela_wire_2704),
        .dout(new_Jinkela_wire_2705)
    );

    bfr new_Jinkela_buffer_4062 (
        .din(new_Jinkela_wire_4760),
        .dout(new_Jinkela_wire_4761)
    );

    spl2 new_Jinkela_splitter_133 (
        .a(new_Jinkela_wire_2819),
        .b(new_Jinkela_wire_2820),
        .c(new_Jinkela_wire_2821)
    );

    bfr new_Jinkela_buffer_4030 (
        .din(new_Jinkela_wire_4726),
        .dout(new_Jinkela_wire_4727)
    );

    bfr new_Jinkela_buffer_2314 (
        .din(new_Jinkela_wire_2705),
        .dout(new_Jinkela_wire_2706)
    );

    bfr new_Jinkela_buffer_4093 (
        .din(new_Jinkela_wire_4793),
        .dout(new_Jinkela_wire_4794)
    );

    bfr new_Jinkela_buffer_2360 (
        .din(new_Jinkela_wire_2756),
        .dout(new_Jinkela_wire_2757)
    );

    bfr new_Jinkela_buffer_4031 (
        .din(new_Jinkela_wire_4727),
        .dout(new_Jinkela_wire_4728)
    );

    bfr new_Jinkela_buffer_2315 (
        .din(new_Jinkela_wire_2706),
        .dout(new_Jinkela_wire_2707)
    );

    bfr new_Jinkela_buffer_4063 (
        .din(new_Jinkela_wire_4761),
        .dout(new_Jinkela_wire_4762)
    );

    bfr new_Jinkela_buffer_2423 (
        .din(new_Jinkela_wire_2821),
        .dout(new_Jinkela_wire_2822)
    );

    bfr new_Jinkela_buffer_4032 (
        .din(new_Jinkela_wire_4728),
        .dout(new_Jinkela_wire_4729)
    );

    bfr new_Jinkela_buffer_2316 (
        .din(new_Jinkela_wire_2707),
        .dout(new_Jinkela_wire_2708)
    );

    bfr new_Jinkela_buffer_2361 (
        .din(new_Jinkela_wire_2757),
        .dout(new_Jinkela_wire_2758)
    );

    bfr new_Jinkela_buffer_4151 (
        .din(n_0479_),
        .dout(new_Jinkela_wire_4864)
    );

    bfr new_Jinkela_buffer_4033 (
        .din(new_Jinkela_wire_4729),
        .dout(new_Jinkela_wire_4730)
    );

    bfr new_Jinkela_buffer_2317 (
        .din(new_Jinkela_wire_2708),
        .dout(new_Jinkela_wire_2709)
    );

    bfr new_Jinkela_buffer_4064 (
        .din(new_Jinkela_wire_4762),
        .dout(new_Jinkela_wire_4763)
    );

    bfr new_Jinkela_buffer_4034 (
        .din(new_Jinkela_wire_4730),
        .dout(new_Jinkela_wire_4731)
    );

    bfr new_Jinkela_buffer_2318 (
        .din(new_Jinkela_wire_2709),
        .dout(new_Jinkela_wire_2710)
    );

    bfr new_Jinkela_buffer_5734 (
        .din(new_Jinkela_wire_6910),
        .dout(new_Jinkela_wire_6911)
    );

    and_bi n_2493_ (
        .a(new_Jinkela_wire_6885),
        .b(new_Jinkela_wire_4432),
        .c(n_0362_)
    );

    bfr new_Jinkela_buffer_5707 (
        .din(new_Jinkela_wire_6875),
        .dout(new_Jinkela_wire_6876)
    );

    bfr new_Jinkela_buffer_6610 (
        .din(n_0424_),
        .dout(new_Jinkela_wire_8086)
    );

    bfr new_Jinkela_buffer_6525 (
        .din(new_Jinkela_wire_7972),
        .dout(new_Jinkela_wire_7973)
    );

    or_bb n_2494_ (
        .a(n_0362_),
        .b(n_0361_),
        .c(new_net_2491)
    );

    bfr new_Jinkela_buffer_3189 (
        .din(new_Jinkela_wire_3643),
        .dout(new_Jinkela_wire_3644)
    );

    bfr new_Jinkela_buffer_6604 (
        .din(n_0954_),
        .dout(new_Jinkela_wire_8076)
    );

    and_bb n_2495_ (
        .a(new_Jinkela_wire_9578),
        .b(new_Jinkela_wire_6639),
        .c(n_0363_)
    );

    spl2 new_Jinkela_splitter_166 (
        .a(n_0317_),
        .b(new_Jinkela_wire_3726),
        .c(new_Jinkela_wire_3727)
    );

    bfr new_Jinkela_buffer_5708 (
        .din(new_Jinkela_wire_6876),
        .dout(new_Jinkela_wire_6877)
    );

    bfr new_Jinkela_buffer_3242 (
        .din(new_Jinkela_wire_3710),
        .dout(new_Jinkela_wire_3711)
    );

    bfr new_Jinkela_buffer_6526 (
        .din(new_Jinkela_wire_7973),
        .dout(new_Jinkela_wire_7974)
    );

    bfr new_Jinkela_buffer_6545 (
        .din(new_Jinkela_wire_8006),
        .dout(new_Jinkela_wire_8007)
    );

    and_ii n_2496_ (
        .a(n_0363_),
        .b(new_Jinkela_wire_5142),
        .c(n_0364_)
    );

    bfr new_Jinkela_buffer_3190 (
        .din(new_Jinkela_wire_3644),
        .dout(new_Jinkela_wire_3645)
    );

    bfr new_Jinkela_buffer_5749 (
        .din(new_Jinkela_wire_6933),
        .dout(new_Jinkela_wire_6934)
    );

    bfr new_Jinkela_buffer_5735 (
        .din(new_Jinkela_wire_6911),
        .dout(new_Jinkela_wire_6912)
    );

    and_bi n_2497_ (
        .a(new_Jinkela_wire_5227),
        .b(new_Jinkela_wire_9884),
        .c(n_0365_)
    );

    bfr new_Jinkela_buffer_5709 (
        .din(new_Jinkela_wire_6877),
        .dout(new_Jinkela_wire_6878)
    );

    bfr new_Jinkela_buffer_6548 (
        .din(new_Jinkela_wire_8011),
        .dout(new_Jinkela_wire_8012)
    );

    bfr new_Jinkela_buffer_6527 (
        .din(new_Jinkela_wire_7974),
        .dout(new_Jinkela_wire_7975)
    );

    and_bi n_2498_ (
        .a(new_Jinkela_wire_9885),
        .b(new_Jinkela_wire_5226),
        .c(n_0366_)
    );

    bfr new_Jinkela_buffer_3191 (
        .din(new_Jinkela_wire_3645),
        .dout(new_Jinkela_wire_3646)
    );

    or_bb n_2499_ (
        .a(n_0366_),
        .b(n_0365_),
        .c(new_net_2521)
    );

    bfr new_Jinkela_buffer_5710 (
        .din(new_Jinkela_wire_6878),
        .dout(new_Jinkela_wire_6879)
    );

    spl2 new_Jinkela_splitter_579 (
        .a(new_Jinkela_wire_8007),
        .b(new_Jinkela_wire_8008),
        .c(new_Jinkela_wire_8009)
    );

    spl3L new_Jinkela_splitter_167 (
        .a(n_1371_),
        .d(new_Jinkela_wire_3728),
        .b(new_Jinkela_wire_3729),
        .c(new_Jinkela_wire_3730)
    );

    bfr new_Jinkela_buffer_6528 (
        .din(new_Jinkela_wire_7975),
        .dout(new_Jinkela_wire_7976)
    );

    and_ii n_2500_ (
        .a(new_Jinkela_wire_4438),
        .b(new_Jinkela_wire_6799),
        .c(n_0367_)
    );

    bfr new_Jinkela_buffer_3192 (
        .din(new_Jinkela_wire_3646),
        .dout(new_Jinkela_wire_3647)
    );

    bfr new_Jinkela_buffer_5757 (
        .din(new_Jinkela_wire_6950),
        .dout(new_Jinkela_wire_6951)
    );

    bfr new_Jinkela_buffer_5736 (
        .din(new_Jinkela_wire_6912),
        .dout(new_Jinkela_wire_6913)
    );

    and_bi n_2501_ (
        .a(new_Jinkela_wire_9577),
        .b(new_Jinkela_wire_9199),
        .c(n_0368_)
    );

    bfr new_Jinkela_buffer_5711 (
        .din(new_Jinkela_wire_6879),
        .dout(new_Jinkela_wire_6880)
    );

    bfr new_Jinkela_buffer_6549 (
        .din(new_Jinkela_wire_8012),
        .dout(new_Jinkela_wire_8013)
    );

    bfr new_Jinkela_buffer_6529 (
        .din(new_Jinkela_wire_7976),
        .dout(new_Jinkela_wire_7977)
    );

    or_bb n_2502_ (
        .a(n_0368_),
        .b(new_Jinkela_wire_5053),
        .c(n_0369_)
    );

    bfr new_Jinkela_buffer_3193 (
        .din(new_Jinkela_wire_3647),
        .dout(new_Jinkela_wire_3648)
    );

    spl2 new_Jinkela_splitter_466 (
        .a(n_0176_),
        .b(new_Jinkela_wire_7014),
        .c(new_Jinkela_wire_7016)
    );

    or_ii n_2503_ (
        .a(new_Jinkela_wire_10555),
        .b(new_Jinkela_wire_5634),
        .c(n_0370_)
    );

    spl2 new_Jinkela_splitter_168 (
        .a(n_1285_),
        .b(new_Jinkela_wire_3731),
        .c(new_Jinkela_wire_3732)
    );

    bfr new_Jinkela_buffer_5712 (
        .din(new_Jinkela_wire_6880),
        .dout(new_Jinkela_wire_6881)
    );

    bfr new_Jinkela_buffer_6530 (
        .din(new_Jinkela_wire_7977),
        .dout(new_Jinkela_wire_7978)
    );

    spl2 new_Jinkela_splitter_583 (
        .a(new_Jinkela_wire_8076),
        .b(new_Jinkela_wire_8077),
        .c(new_Jinkela_wire_8078)
    );

    and_ii n_2504_ (
        .a(new_Jinkela_wire_10554),
        .b(new_Jinkela_wire_5633),
        .c(n_0371_)
    );

    bfr new_Jinkela_buffer_3194 (
        .din(new_Jinkela_wire_3648),
        .dout(new_Jinkela_wire_3649)
    );

    bfr new_Jinkela_buffer_5750 (
        .din(new_Jinkela_wire_6934),
        .dout(new_Jinkela_wire_6935)
    );

    bfr new_Jinkela_buffer_5737 (
        .din(new_Jinkela_wire_6913),
        .dout(new_Jinkela_wire_6914)
    );

    and_bi n_2505_ (
        .a(n_0370_),
        .b(n_0371_),
        .c(new_net_2566)
    );

    spl2 new_Jinkela_splitter_171 (
        .a(n_0942_),
        .b(new_Jinkela_wire_3769),
        .c(new_Jinkela_wire_3770)
    );

    bfr new_Jinkela_buffer_5713 (
        .din(new_Jinkela_wire_6881),
        .dout(new_Jinkela_wire_6882)
    );

    bfr new_Jinkela_buffer_3244 (
        .din(n_0080_),
        .dout(new_Jinkela_wire_3733)
    );

    bfr new_Jinkela_buffer_6531 (
        .din(new_Jinkela_wire_7978),
        .dout(new_Jinkela_wire_7979)
    );

    bfr new_Jinkela_buffer_6605 (
        .din(n_1344_),
        .dout(new_Jinkela_wire_8079)
    );

    and_ii n_2506_ (
        .a(new_Jinkela_wire_5013),
        .b(new_Jinkela_wire_9159),
        .c(n_0372_)
    );

    bfr new_Jinkela_buffer_3195 (
        .din(new_Jinkela_wire_3649),
        .dout(new_Jinkela_wire_3650)
    );

    or_ii n_2507_ (
        .a(new_Jinkela_wire_9573),
        .b(new_Jinkela_wire_7540),
        .c(n_0373_)
    );

    spl2 new_Jinkela_splitter_172 (
        .a(n_0912_),
        .b(new_Jinkela_wire_3771),
        .c(new_Jinkela_wire_3772)
    );

    bfr new_Jinkela_buffer_5714 (
        .din(new_Jinkela_wire_6882),
        .dout(new_Jinkela_wire_6883)
    );

    bfr new_Jinkela_buffer_3245 (
        .din(new_Jinkela_wire_3733),
        .dout(new_Jinkela_wire_3734)
    );

    bfr new_Jinkela_buffer_6532 (
        .din(new_Jinkela_wire_7979),
        .dout(new_Jinkela_wire_7980)
    );

    bfr new_Jinkela_buffer_6550 (
        .din(new_Jinkela_wire_8013),
        .dout(new_Jinkela_wire_8014)
    );

    and_ii n_2508_ (
        .a(new_Jinkela_wire_9575),
        .b(new_Jinkela_wire_7539),
        .c(n_0374_)
    );

    bfr new_Jinkela_buffer_3196 (
        .din(new_Jinkela_wire_3650),
        .dout(new_Jinkela_wire_3651)
    );

    spl2 new_Jinkela_splitter_463 (
        .a(new_Jinkela_wire_6944),
        .b(new_Jinkela_wire_6945),
        .c(new_Jinkela_wire_6946)
    );

    bfr new_Jinkela_buffer_5738 (
        .din(new_Jinkela_wire_6914),
        .dout(new_Jinkela_wire_6915)
    );

    and_bi n_2509_ (
        .a(n_0373_),
        .b(n_0374_),
        .c(new_net_2549)
    );

    bfr new_Jinkela_buffer_5715 (
        .din(new_Jinkela_wire_6883),
        .dout(new_Jinkela_wire_6884)
    );

    bfr new_Jinkela_buffer_6533 (
        .din(new_Jinkela_wire_7980),
        .dout(new_Jinkela_wire_7981)
    );

    or_ii n_2510_ (
        .a(new_Jinkela_wire_7019),
        .b(new_Jinkela_wire_8160),
        .c(n_0375_)
    );

    bfr new_Jinkela_buffer_3197 (
        .din(new_Jinkela_wire_3651),
        .dout(new_Jinkela_wire_3652)
    );

    and_bi n_2511_ (
        .a(new_Jinkela_wire_4736),
        .b(new_Jinkela_wire_7017),
        .c(n_0376_)
    );

    bfr new_Jinkela_buffer_3276 (
        .din(n_0866_),
        .dout(new_Jinkela_wire_3773)
    );

    spl2 new_Jinkela_splitter_454 (
        .a(new_Jinkela_wire_6884),
        .b(new_Jinkela_wire_6885),
        .c(new_Jinkela_wire_6886)
    );

    bfr new_Jinkela_buffer_3246 (
        .din(new_Jinkela_wire_3734),
        .dout(new_Jinkela_wire_3735)
    );

    bfr new_Jinkela_buffer_6534 (
        .din(new_Jinkela_wire_7981),
        .dout(new_Jinkela_wire_7982)
    );

    bfr new_Jinkela_buffer_6551 (
        .din(new_Jinkela_wire_8014),
        .dout(new_Jinkela_wire_8015)
    );

    and_bi n_2512_ (
        .a(n_0375_),
        .b(n_0376_),
        .c(n_0377_)
    );

    bfr new_Jinkela_buffer_3198 (
        .din(new_Jinkela_wire_3652),
        .dout(new_Jinkela_wire_3653)
    );

    or_ii n_2513_ (
        .a(new_Jinkela_wire_7263),
        .b(new_Jinkela_wire_7010),
        .c(n_0378_)
    );

    bfr new_Jinkela_buffer_5751 (
        .din(new_Jinkela_wire_6935),
        .dout(new_Jinkela_wire_6936)
    );

    bfr new_Jinkela_buffer_6606 (
        .din(new_Jinkela_wire_8079),
        .dout(new_Jinkela_wire_8080)
    );

    bfr new_Jinkela_buffer_5739 (
        .din(new_Jinkela_wire_6915),
        .dout(new_Jinkela_wire_6916)
    );

    bfr new_Jinkela_buffer_6535 (
        .din(new_Jinkela_wire_7982),
        .dout(new_Jinkela_wire_7983)
    );

    inv n_2514_ (
        .din(new_Jinkela_wire_6948),
        .dout(n_0379_)
    );

    bfr new_Jinkela_buffer_3199 (
        .din(new_Jinkela_wire_3653),
        .dout(new_Jinkela_wire_3654)
    );

    bfr new_Jinkela_buffer_5740 (
        .din(new_Jinkela_wire_6916),
        .dout(new_Jinkela_wire_6917)
    );

    and_bi n_2515_ (
        .a(new_Jinkela_wire_8070),
        .b(new_Jinkela_wire_7262),
        .c(n_0380_)
    );

    spl2 new_Jinkela_splitter_175 (
        .a(n_1207_),
        .b(new_Jinkela_wire_3783),
        .c(new_Jinkela_wire_3784)
    );

    bfr new_Jinkela_buffer_6552 (
        .din(new_Jinkela_wire_8015),
        .dout(new_Jinkela_wire_8016)
    );

    bfr new_Jinkela_buffer_3247 (
        .din(new_Jinkela_wire_3735),
        .dout(new_Jinkela_wire_3736)
    );

    bfr new_Jinkela_buffer_6536 (
        .din(new_Jinkela_wire_7983),
        .dout(new_Jinkela_wire_7984)
    );

    and_bi n_2516_ (
        .a(n_0378_),
        .b(n_0380_),
        .c(new_net_8)
    );

    bfr new_Jinkela_buffer_3200 (
        .din(new_Jinkela_wire_3654),
        .dout(new_Jinkela_wire_3655)
    );

    bfr new_Jinkela_buffer_5752 (
        .din(new_Jinkela_wire_6936),
        .dout(new_Jinkela_wire_6937)
    );

    bfr new_Jinkela_buffer_5741 (
        .din(new_Jinkela_wire_6917),
        .dout(new_Jinkela_wire_6918)
    );

    and_bb n_2517_ (
        .a(new_Jinkela_wire_7015),
        .b(new_Jinkela_wire_4392),
        .c(n_0381_)
    );

    bfr new_Jinkela_buffer_6607 (
        .din(new_Jinkela_wire_8080),
        .dout(new_Jinkela_wire_8081)
    );

    bfr new_Jinkela_buffer_3279 (
        .din(n_0450_),
        .dout(new_Jinkela_wire_3778)
    );

    and_bi n_2518_ (
        .a(new_Jinkela_wire_9136),
        .b(new_Jinkela_wire_10432),
        .c(new_net_9)
    );

    bfr new_Jinkela_buffer_3201 (
        .din(new_Jinkela_wire_3655),
        .dout(new_Jinkela_wire_3656)
    );

    bfr new_Jinkela_buffer_5819 (
        .din(n_1363_),
        .dout(new_Jinkela_wire_7021)
    );

    bfr new_Jinkela_buffer_5742 (
        .din(new_Jinkela_wire_6918),
        .dout(new_Jinkela_wire_6919)
    );

    bfr new_Jinkela_buffer_6553 (
        .din(new_Jinkela_wire_8016),
        .dout(new_Jinkela_wire_8017)
    );

    and_ii n_2519_ (
        .a(new_Jinkela_wire_6674),
        .b(new_Jinkela_wire_7651),
        .c(n_0382_)
    );

    bfr new_Jinkela_buffer_3277 (
        .din(new_Jinkela_wire_3773),
        .dout(new_Jinkela_wire_3774)
    );

    spl2 new_Jinkela_splitter_587 (
        .a(n_0783_),
        .b(new_Jinkela_wire_8093),
        .c(new_Jinkela_wire_8094)
    );

    bfr new_Jinkela_buffer_3248 (
        .din(new_Jinkela_wire_3736),
        .dout(new_Jinkela_wire_3737)
    );

    spl2 new_Jinkela_splitter_465 (
        .a(new_Jinkela_wire_7011),
        .b(new_Jinkela_wire_7012),
        .c(new_Jinkela_wire_7013)
    );

    or_bi n_2520_ (
        .a(new_Jinkela_wire_4120),
        .b(new_Jinkela_wire_8071),
        .c(n_0383_)
    );

    bfr new_Jinkela_buffer_3202 (
        .din(new_Jinkela_wire_3656),
        .dout(new_Jinkela_wire_3657)
    );

    bfr new_Jinkela_buffer_5753 (
        .din(new_Jinkela_wire_6937),
        .dout(new_Jinkela_wire_6938)
    );

    bfr new_Jinkela_buffer_5743 (
        .din(new_Jinkela_wire_6919),
        .dout(new_Jinkela_wire_6920)
    );

    bfr new_Jinkela_buffer_6554 (
        .din(new_Jinkela_wire_8017),
        .dout(new_Jinkela_wire_8018)
    );

    and_bi n_2521_ (
        .a(new_Jinkela_wire_4119),
        .b(new_Jinkela_wire_8072),
        .c(n_0384_)
    );

    spl2 new_Jinkela_splitter_586 (
        .a(n_1278_),
        .b(new_Jinkela_wire_8091),
        .c(new_Jinkela_wire_8092)
    );

    and_bi n_2522_ (
        .a(n_0383_),
        .b(n_0384_),
        .c(new_net_2509)
    );

    bfr new_Jinkela_buffer_3203 (
        .din(new_Jinkela_wire_3657),
        .dout(new_Jinkela_wire_3658)
    );

    bfr new_Jinkela_buffer_5758 (
        .din(new_Jinkela_wire_6951),
        .dout(new_Jinkela_wire_6952)
    );

    bfr new_Jinkela_buffer_5744 (
        .din(new_Jinkela_wire_6920),
        .dout(new_Jinkela_wire_6921)
    );

    bfr new_Jinkela_buffer_6555 (
        .din(new_Jinkela_wire_8018),
        .dout(new_Jinkela_wire_8019)
    );

    and_ii n_2523_ (
        .a(new_Jinkela_wire_6807),
        .b(new_Jinkela_wire_6534),
        .c(n_0385_)
    );

    bfr new_Jinkela_buffer_3282 (
        .din(n_1346_),
        .dout(new_Jinkela_wire_3787)
    );

    bfr new_Jinkela_buffer_6611 (
        .din(new_Jinkela_wire_8086),
        .dout(new_Jinkela_wire_8087)
    );

    bfr new_Jinkela_buffer_3249 (
        .din(new_Jinkela_wire_3737),
        .dout(new_Jinkela_wire_3738)
    );

    bfr new_Jinkela_buffer_6615 (
        .din(n_0219_),
        .dout(new_Jinkela_wire_8097)
    );

    and_bb n_2524_ (
        .a(new_Jinkela_wire_9422),
        .b(new_Jinkela_wire_5754),
        .c(n_0386_)
    );

    bfr new_Jinkela_buffer_3204 (
        .din(new_Jinkela_wire_3658),
        .dout(new_Jinkela_wire_3659)
    );

    bfr new_Jinkela_buffer_5754 (
        .din(new_Jinkela_wire_6938),
        .dout(new_Jinkela_wire_6939)
    );

    spl2 new_Jinkela_splitter_458 (
        .a(new_Jinkela_wire_6921),
        .b(new_Jinkela_wire_6922),
        .c(new_Jinkela_wire_6923)
    );

    spl3L new_Jinkela_splitter_580 (
        .a(new_Jinkela_wire_8019),
        .d(new_Jinkela_wire_8020),
        .b(new_Jinkela_wire_8021),
        .c(new_Jinkela_wire_8022)
    );

    and_ii n_2525_ (
        .a(n_0386_),
        .b(new_Jinkela_wire_10553),
        .c(n_0387_)
    );

    bfr new_Jinkela_buffer_6608 (
        .din(new_Jinkela_wire_8081),
        .dout(new_Jinkela_wire_8082)
    );

    bfr new_Jinkela_buffer_5745 (
        .din(new_Jinkela_wire_6923),
        .dout(new_Jinkela_wire_6924)
    );

    or_ii n_2526_ (
        .a(new_Jinkela_wire_8282),
        .b(new_Jinkela_wire_5196),
        .c(n_0388_)
    );

    bfr new_Jinkela_buffer_3205 (
        .din(new_Jinkela_wire_3659),
        .dout(new_Jinkela_wire_3660)
    );

    bfr new_Jinkela_buffer_6556 (
        .din(new_Jinkela_wire_8022),
        .dout(new_Jinkela_wire_8023)
    );

    or_bb n_2527_ (
        .a(new_Jinkela_wire_8281),
        .b(new_Jinkela_wire_5195),
        .c(n_0389_)
    );

    bfr new_Jinkela_buffer_3278 (
        .din(new_Jinkela_wire_3774),
        .dout(new_Jinkela_wire_3775)
    );

    bfr new_Jinkela_buffer_3250 (
        .din(new_Jinkela_wire_3738),
        .dout(new_Jinkela_wire_3739)
    );

    or_ii n_2528_ (
        .a(n_0389_),
        .b(n_0388_),
        .c(new_net_2503)
    );

    bfr new_Jinkela_buffer_3206 (
        .din(new_Jinkela_wire_3660),
        .dout(new_Jinkela_wire_3661)
    );

    bfr new_Jinkela_buffer_5759 (
        .din(new_Jinkela_wire_6952),
        .dout(new_Jinkela_wire_6953)
    );

    spl2 new_Jinkela_splitter_459 (
        .a(new_Jinkela_wire_6924),
        .b(new_Jinkela_wire_6925),
        .c(new_Jinkela_wire_6926)
    );

    bfr new_Jinkela_buffer_6557 (
        .din(new_Jinkela_wire_8023),
        .dout(new_Jinkela_wire_8024)
    );

    inv n_2529_ (
        .din(new_Jinkela_wire_3791),
        .dout(n_0390_)
    );

    bfr new_Jinkela_buffer_6609 (
        .din(new_Jinkela_wire_8082),
        .dout(new_Jinkela_wire_8083)
    );

    spl4L new_Jinkela_splitter_467 (
        .a(new_Jinkela_wire_7016),
        .d(new_Jinkela_wire_7017),
        .b(new_Jinkela_wire_7018),
        .e(new_Jinkela_wire_7019),
        .c(new_Jinkela_wire_7020)
    );

    and_ii n_2530_ (
        .a(new_Jinkela_wire_9423),
        .b(new_Jinkela_wire_4336),
        .c(n_0391_)
    );

    bfr new_Jinkela_buffer_3207 (
        .din(new_Jinkela_wire_3661),
        .dout(new_Jinkela_wire_3662)
    );

    bfr new_Jinkela_buffer_5760 (
        .din(new_Jinkela_wire_6953),
        .dout(new_Jinkela_wire_6954)
    );

    bfr new_Jinkela_buffer_6558 (
        .din(new_Jinkela_wire_8024),
        .dout(new_Jinkela_wire_8025)
    );

    or_bb n_2531_ (
        .a(n_0391_),
        .b(new_Jinkela_wire_9803),
        .c(n_0392_)
    );

    bfr new_Jinkela_buffer_6612 (
        .din(new_Jinkela_wire_8087),
        .dout(new_Jinkela_wire_8088)
    );

    bfr new_Jinkela_buffer_3251 (
        .din(new_Jinkela_wire_3739),
        .dout(new_Jinkela_wire_3740)
    );

    or_ii n_2532_ (
        .a(new_Jinkela_wire_6098),
        .b(new_Jinkela_wire_8356),
        .c(n_0393_)
    );

    bfr new_Jinkela_buffer_3208 (
        .din(new_Jinkela_wire_3662),
        .dout(new_Jinkela_wire_3663)
    );

    bfr new_Jinkela_buffer_6559 (
        .din(new_Jinkela_wire_8025),
        .dout(new_Jinkela_wire_8026)
    );

    and_bi n_2533_ (
        .a(new_Jinkela_wire_3821),
        .b(new_Jinkela_wire_6097),
        .c(n_0394_)
    );

    spl4L new_Jinkela_splitter_174 (
        .a(n_1306_),
        .d(new_Jinkela_wire_3779),
        .b(new_Jinkela_wire_3780),
        .e(new_Jinkela_wire_3781),
        .c(new_Jinkela_wire_3782)
    );

    bfr new_Jinkela_buffer_5761 (
        .din(new_Jinkela_wire_6954),
        .dout(new_Jinkela_wire_6955)
    );

    spl2 new_Jinkela_splitter_584 (
        .a(new_Jinkela_wire_8083),
        .b(new_Jinkela_wire_8084),
        .c(new_Jinkela_wire_8085)
    );

    and_bi n_2534_ (
        .a(n_0393_),
        .b(n_0394_),
        .c(new_net_2574)
    );

    bfr new_Jinkela_buffer_3209 (
        .din(new_Jinkela_wire_3663),
        .dout(new_Jinkela_wire_3664)
    );

    bfr new_Jinkela_buffer_5818 (
        .din(new_Jinkela_wire_7014),
        .dout(new_Jinkela_wire_7015)
    );

    bfr new_Jinkela_buffer_6560 (
        .din(new_Jinkela_wire_8026),
        .dout(new_Jinkela_wire_8027)
    );

    bfr new_Jinkela_buffer_4866 (
        .din(new_Jinkela_wire_5800),
        .dout(new_Jinkela_wire_5801)
    );

    and_ii n_1779_ (
        .a(new_Jinkela_wire_7077),
        .b(new_Jinkela_wire_8166),
        .c(n_1046_)
    );

    bfr new_Jinkela_buffer_8457 (
        .din(new_Jinkela_wire_10622),
        .dout(new_Jinkela_wire_10623)
    );

    and_bb n_1780_ (
        .a(new_Jinkela_wire_7076),
        .b(new_Jinkela_wire_8165),
        .c(n_1047_)
    );

    bfr new_Jinkela_buffer_4942 (
        .din(new_Jinkela_wire_5891),
        .dout(new_Jinkela_wire_5892)
    );

    bfr new_Jinkela_buffer_4867 (
        .din(new_Jinkela_wire_5801),
        .dout(new_Jinkela_wire_5802)
    );

    and_ii n_1781_ (
        .a(n_1047_),
        .b(n_1046_),
        .c(n_1048_)
    );

    bfr new_Jinkela_buffer_8458 (
        .din(new_Jinkela_wire_10623),
        .dout(new_Jinkela_wire_10624)
    );

    and_bi n_1782_ (
        .a(new_Jinkela_wire_2893),
        .b(new_Jinkela_wire_1353),
        .c(n_1049_)
    );

    bfr new_Jinkela_buffer_4891 (
        .din(new_Jinkela_wire_5827),
        .dout(new_Jinkela_wire_5828)
    );

    spl2 new_Jinkela_splitter_356 (
        .a(new_Jinkela_wire_5802),
        .b(new_Jinkela_wire_5803),
        .c(new_Jinkela_wire_5804)
    );

    and_bi n_1783_ (
        .a(new_Jinkela_wire_1273),
        .b(new_Jinkela_wire_363),
        .c(n_1050_)
    );

    spl2 new_Jinkela_splitter_364 (
        .a(n_0471_),
        .b(new_Jinkela_wire_5933),
        .c(new_Jinkela_wire_5934)
    );

    spl4L new_Jinkela_splitter_870 (
        .a(new_Jinkela_wire_10624),
        .d(new_Jinkela_wire_10625),
        .b(new_Jinkela_wire_10626),
        .e(new_Jinkela_wire_10627),
        .c(new_Jinkela_wire_10628)
    );

    and_ii n_1784_ (
        .a(n_1050_),
        .b(n_1049_),
        .c(n_1051_)
    );

    bfr new_Jinkela_buffer_4892 (
        .din(new_Jinkela_wire_5828),
        .dout(new_Jinkela_wire_5829)
    );

    and_bi n_1785_ (
        .a(new_Jinkela_wire_2076),
        .b(new_Jinkela_wire_1348),
        .c(n_1052_)
    );

    and_bi n_1786_ (
        .a(new_Jinkela_wire_1241),
        .b(new_Jinkela_wire_3205),
        .c(n_1053_)
    );

    spl2 new_Jinkela_splitter_365 (
        .a(n_0081_),
        .b(new_Jinkela_wire_5935),
        .c(new_Jinkela_wire_5936)
    );

    bfr new_Jinkela_buffer_4948 (
        .din(new_Jinkela_wire_5897),
        .dout(new_Jinkela_wire_5898)
    );

    and_ii n_1787_ (
        .a(n_1053_),
        .b(n_1052_),
        .c(n_1054_)
    );

    bfr new_Jinkela_buffer_4893 (
        .din(new_Jinkela_wire_5829),
        .dout(new_Jinkela_wire_5830)
    );

    and_ii n_1788_ (
        .a(new_Jinkela_wire_4234),
        .b(new_Jinkela_wire_6928),
        .c(n_1055_)
    );

    bfr new_Jinkela_buffer_4969 (
        .din(new_Jinkela_wire_5920),
        .dout(new_Jinkela_wire_5921)
    );

    and_bb n_1789_ (
        .a(new_Jinkela_wire_4233),
        .b(new_Jinkela_wire_6927),
        .c(n_1056_)
    );

    bfr new_Jinkela_buffer_4894 (
        .din(new_Jinkela_wire_5830),
        .dout(new_Jinkela_wire_5831)
    );

    and_ii n_1790_ (
        .a(n_1056_),
        .b(n_1055_),
        .c(n_1057_)
    );

    bfr new_Jinkela_buffer_4949 (
        .din(new_Jinkela_wire_5898),
        .dout(new_Jinkela_wire_5899)
    );

    and_ii n_1791_ (
        .a(new_Jinkela_wire_8822),
        .b(new_Jinkela_wire_6246),
        .c(n_1058_)
    );

    bfr new_Jinkela_buffer_4895 (
        .din(new_Jinkela_wire_5831),
        .dout(new_Jinkela_wire_5832)
    );

    and_bb n_1792_ (
        .a(new_Jinkela_wire_8821),
        .b(new_Jinkela_wire_6245),
        .c(n_1059_)
    );

    bfr new_Jinkela_buffer_4975 (
        .din(new_Jinkela_wire_5928),
        .dout(new_Jinkela_wire_5929)
    );

    and_ii n_1793_ (
        .a(n_1059_),
        .b(n_1058_),
        .c(n_1060_)
    );

    bfr new_Jinkela_buffer_4896 (
        .din(new_Jinkela_wire_5832),
        .dout(new_Jinkela_wire_5833)
    );

    or_bb n_1794_ (
        .a(new_Jinkela_wire_7346),
        .b(new_Jinkela_wire_8075),
        .c(n_1061_)
    );

    bfr new_Jinkela_buffer_4950 (
        .din(new_Jinkela_wire_5899),
        .dout(new_Jinkela_wire_5900)
    );

    and_bb n_1795_ (
        .a(new_Jinkela_wire_7345),
        .b(new_Jinkela_wire_8074),
        .c(n_1062_)
    );

    bfr new_Jinkela_buffer_4897 (
        .din(new_Jinkela_wire_5833),
        .dout(new_Jinkela_wire_5834)
    );

    and_bi n_1796_ (
        .a(n_1061_),
        .b(n_1062_),
        .c(n_1063_)
    );

    bfr new_Jinkela_buffer_4970 (
        .din(new_Jinkela_wire_5921),
        .dout(new_Jinkela_wire_5922)
    );

    and_bi n_1797_ (
        .a(new_Jinkela_wire_176),
        .b(new_Jinkela_wire_1367),
        .c(n_1064_)
    );

    bfr new_Jinkela_buffer_4898 (
        .din(new_Jinkela_wire_5834),
        .dout(new_Jinkela_wire_5835)
    );

    and_bi n_1798_ (
        .a(new_Jinkela_wire_1175),
        .b(new_Jinkela_wire_2084),
        .c(n_1065_)
    );

    bfr new_Jinkela_buffer_4951 (
        .din(new_Jinkela_wire_5900),
        .dout(new_Jinkela_wire_5901)
    );

    and_ii n_1799_ (
        .a(n_1065_),
        .b(n_1064_),
        .c(n_1066_)
    );

    bfr new_Jinkela_buffer_4899 (
        .din(new_Jinkela_wire_5835),
        .dout(new_Jinkela_wire_5836)
    );

    and_bi n_1800_ (
        .a(new_Jinkela_wire_787),
        .b(new_Jinkela_wire_1332),
        .c(n_1067_)
    );

    bfr new_Jinkela_buffer_5010 (
        .din(n_0171_),
        .dout(new_Jinkela_wire_5970)
    );

    and_bi n_1801_ (
        .a(new_Jinkela_wire_1380),
        .b(new_Jinkela_wire_442),
        .c(n_1068_)
    );

    bfr new_Jinkela_buffer_4900 (
        .din(new_Jinkela_wire_5836),
        .dout(new_Jinkela_wire_5837)
    );

    and_ii n_1802_ (
        .a(n_1068_),
        .b(n_1067_),
        .c(n_1069_)
    );

    bfr new_Jinkela_buffer_4952 (
        .din(new_Jinkela_wire_5901),
        .dout(new_Jinkela_wire_5902)
    );

    or_bb n_1803_ (
        .a(new_Jinkela_wire_8751),
        .b(new_Jinkela_wire_3584),
        .c(n_1070_)
    );

    bfr new_Jinkela_buffer_4901 (
        .din(new_Jinkela_wire_5837),
        .dout(new_Jinkela_wire_5838)
    );

    and_bb n_1804_ (
        .a(new_Jinkela_wire_8752),
        .b(new_Jinkela_wire_3583),
        .c(n_1071_)
    );

    spl2 new_Jinkela_splitter_363 (
        .a(new_Jinkela_wire_5922),
        .b(new_Jinkela_wire_5923),
        .c(new_Jinkela_wire_5924)
    );

    and_bi n_1805_ (
        .a(n_1070_),
        .b(n_1071_),
        .c(n_1072_)
    );

    bfr new_Jinkela_buffer_4902 (
        .din(new_Jinkela_wire_5838),
        .dout(new_Jinkela_wire_5839)
    );

    and_bi n_1806_ (
        .a(new_Jinkela_wire_594),
        .b(new_Jinkela_wire_1364),
        .c(n_1073_)
    );

    bfr new_Jinkela_buffer_4953 (
        .din(new_Jinkela_wire_5902),
        .dout(new_Jinkela_wire_5903)
    );

    and_bi n_1807_ (
        .a(new_Jinkela_wire_1173),
        .b(new_Jinkela_wire_2666),
        .c(n_1074_)
    );

    bfr new_Jinkela_buffer_4903 (
        .din(new_Jinkela_wire_5839),
        .dout(new_Jinkela_wire_5840)
    );

    and_ii n_1808_ (
        .a(n_1074_),
        .b(n_1073_),
        .c(n_1075_)
    );

    bfr new_Jinkela_buffer_4971 (
        .din(new_Jinkela_wire_5924),
        .dout(new_Jinkela_wire_5925)
    );

    and_bi n_1809_ (
        .a(new_Jinkela_wire_3442),
        .b(new_Jinkela_wire_1191),
        .c(n_1076_)
    );

    bfr new_Jinkela_buffer_4904 (
        .din(new_Jinkela_wire_5840),
        .dout(new_Jinkela_wire_5841)
    );

    and_bi n_1810_ (
        .a(new_Jinkela_wire_1229),
        .b(new_Jinkela_wire_3124),
        .c(n_1077_)
    );

    bfr new_Jinkela_buffer_4954 (
        .din(new_Jinkela_wire_5903),
        .dout(new_Jinkela_wire_5904)
    );

    and_ii n_1811_ (
        .a(n_1077_),
        .b(n_1076_),
        .c(n_1078_)
    );

    bfr new_Jinkela_buffer_4905 (
        .din(new_Jinkela_wire_5841),
        .dout(new_Jinkela_wire_5842)
    );

    or_bi n_1812_ (
        .a(new_Jinkela_wire_9544),
        .b(new_Jinkela_wire_7093),
        .c(n_1079_)
    );

    bfr new_Jinkela_buffer_4976 (
        .din(new_Jinkela_wire_5929),
        .dout(new_Jinkela_wire_5930)
    );

    and_bi n_1813_ (
        .a(new_Jinkela_wire_9543),
        .b(new_Jinkela_wire_7092),
        .c(n_1080_)
    );

    bfr new_Jinkela_buffer_4906 (
        .din(new_Jinkela_wire_5842),
        .dout(new_Jinkela_wire_5843)
    );

    and_bi n_1814_ (
        .a(n_1079_),
        .b(n_1080_),
        .c(n_1081_)
    );

    bfr new_Jinkela_buffer_4955 (
        .din(new_Jinkela_wire_5904),
        .dout(new_Jinkela_wire_5905)
    );

    and_ii n_1815_ (
        .a(new_Jinkela_wire_7296),
        .b(new_Jinkela_wire_8716),
        .c(n_1082_)
    );

    bfr new_Jinkela_buffer_4907 (
        .din(new_Jinkela_wire_5843),
        .dout(new_Jinkela_wire_5844)
    );

    and_bb n_1816_ (
        .a(new_Jinkela_wire_7295),
        .b(new_Jinkela_wire_8715),
        .c(n_1083_)
    );

    and_ii n_1817_ (
        .a(n_1083_),
        .b(n_1082_),
        .c(n_1084_)
    );

    bfr new_Jinkela_buffer_4908 (
        .din(new_Jinkela_wire_5844),
        .dout(new_Jinkela_wire_5845)
    );

    and_bi n_1818_ (
        .a(new_Jinkela_wire_79),
        .b(new_Jinkela_wire_1197),
        .c(n_1085_)
    );

    bfr new_Jinkela_buffer_4956 (
        .din(new_Jinkela_wire_5905),
        .dout(new_Jinkela_wire_5906)
    );

    and_bi n_1819_ (
        .a(new_Jinkela_wire_1356),
        .b(new_Jinkela_wire_3446),
        .c(n_1086_)
    );

    bfr new_Jinkela_buffer_4909 (
        .din(new_Jinkela_wire_5845),
        .dout(new_Jinkela_wire_5846)
    );

    and_ii n_1820_ (
        .a(n_1086_),
        .b(n_1085_),
        .c(n_1087_)
    );

    bfr new_Jinkela_buffer_4094 (
        .din(new_Jinkela_wire_4794),
        .dout(new_Jinkela_wire_4795)
    );

    bfr new_Jinkela_buffer_4035 (
        .din(new_Jinkela_wire_4731),
        .dout(new_Jinkela_wire_4732)
    );

    bfr new_Jinkela_buffer_4065 (
        .din(new_Jinkela_wire_4763),
        .dout(new_Jinkela_wire_4764)
    );

    bfr new_Jinkela_buffer_4036 (
        .din(new_Jinkela_wire_4732),
        .dout(new_Jinkela_wire_4733)
    );

    spl3L new_Jinkela_splitter_269 (
        .a(n_0401_),
        .d(new_Jinkela_wire_4914),
        .b(new_Jinkela_wire_4915),
        .c(new_Jinkela_wire_4916)
    );

    bfr new_Jinkela_buffer_4123 (
        .din(new_Jinkela_wire_4823),
        .dout(new_Jinkela_wire_4824)
    );

    bfr new_Jinkela_buffer_4037 (
        .din(new_Jinkela_wire_4733),
        .dout(new_Jinkela_wire_4734)
    );

    bfr new_Jinkela_buffer_4066 (
        .din(new_Jinkela_wire_4764),
        .dout(new_Jinkela_wire_4765)
    );

    bfr new_Jinkela_buffer_4038 (
        .din(new_Jinkela_wire_4734),
        .dout(new_Jinkela_wire_4735)
    );

    bfr new_Jinkela_buffer_4095 (
        .din(new_Jinkela_wire_4795),
        .dout(new_Jinkela_wire_4796)
    );

    spl2 new_Jinkela_splitter_257 (
        .a(new_Jinkela_wire_4735),
        .b(new_Jinkela_wire_4736),
        .c(new_Jinkela_wire_4737)
    );

    spl4L new_Jinkela_splitter_266 (
        .a(n_1160_),
        .d(new_Jinkela_wire_4871),
        .b(new_Jinkela_wire_4872),
        .e(new_Jinkela_wire_4873),
        .c(new_Jinkela_wire_4874)
    );

    bfr new_Jinkela_buffer_4067 (
        .din(new_Jinkela_wire_4765),
        .dout(new_Jinkela_wire_4766)
    );

    bfr new_Jinkela_buffer_4068 (
        .din(new_Jinkela_wire_4766),
        .dout(new_Jinkela_wire_4767)
    );

    bfr new_Jinkela_buffer_4096 (
        .din(new_Jinkela_wire_4796),
        .dout(new_Jinkela_wire_4797)
    );

    bfr new_Jinkela_buffer_4069 (
        .din(new_Jinkela_wire_4767),
        .dout(new_Jinkela_wire_4768)
    );

    bfr new_Jinkela_buffer_4153 (
        .din(new_Jinkela_wire_4865),
        .dout(new_Jinkela_wire_4866)
    );

    bfr new_Jinkela_buffer_4124 (
        .din(new_Jinkela_wire_4824),
        .dout(new_Jinkela_wire_4825)
    );

    bfr new_Jinkela_buffer_4070 (
        .din(new_Jinkela_wire_4768),
        .dout(new_Jinkela_wire_4769)
    );

    bfr new_Jinkela_buffer_4097 (
        .din(new_Jinkela_wire_4797),
        .dout(new_Jinkela_wire_4798)
    );

    bfr new_Jinkela_buffer_4071 (
        .din(new_Jinkela_wire_4769),
        .dout(new_Jinkela_wire_4770)
    );

    bfr new_Jinkela_buffer_4152 (
        .din(new_Jinkela_wire_4864),
        .dout(new_Jinkela_wire_4865)
    );

    bfr new_Jinkela_buffer_4072 (
        .din(new_Jinkela_wire_4770),
        .dout(new_Jinkela_wire_4771)
    );

    bfr new_Jinkela_buffer_4098 (
        .din(new_Jinkela_wire_4798),
        .dout(new_Jinkela_wire_4799)
    );

    bfr new_Jinkela_buffer_4073 (
        .din(new_Jinkela_wire_4771),
        .dout(new_Jinkela_wire_4772)
    );

    bfr new_Jinkela_buffer_4125 (
        .din(new_Jinkela_wire_4825),
        .dout(new_Jinkela_wire_4826)
    );

    bfr new_Jinkela_buffer_4074 (
        .din(new_Jinkela_wire_4772),
        .dout(new_Jinkela_wire_4773)
    );

    bfr new_Jinkela_buffer_4099 (
        .din(new_Jinkela_wire_4799),
        .dout(new_Jinkela_wire_4800)
    );

    bfr new_Jinkela_buffer_4075 (
        .din(new_Jinkela_wire_4773),
        .dout(new_Jinkela_wire_4774)
    );

    bfr new_Jinkela_buffer_4076 (
        .din(new_Jinkela_wire_4774),
        .dout(new_Jinkela_wire_4775)
    );

    bfr new_Jinkela_buffer_4100 (
        .din(new_Jinkela_wire_4800),
        .dout(new_Jinkela_wire_4801)
    );

    bfr new_Jinkela_buffer_4077 (
        .din(new_Jinkela_wire_4775),
        .dout(new_Jinkela_wire_4776)
    );

    bfr new_Jinkela_buffer_4126 (
        .din(new_Jinkela_wire_4826),
        .dout(new_Jinkela_wire_4827)
    );

    bfr new_Jinkela_buffer_4078 (
        .din(new_Jinkela_wire_4776),
        .dout(new_Jinkela_wire_4777)
    );

    bfr new_Jinkela_buffer_4101 (
        .din(new_Jinkela_wire_4801),
        .dout(new_Jinkela_wire_4802)
    );

    bfr new_Jinkela_buffer_4079 (
        .din(new_Jinkela_wire_4777),
        .dout(new_Jinkela_wire_4778)
    );

    bfr new_Jinkela_buffer_4080 (
        .din(new_Jinkela_wire_4778),
        .dout(new_Jinkela_wire_4779)
    );

    bfr new_Jinkela_buffer_4102 (
        .din(new_Jinkela_wire_4802),
        .dout(new_Jinkela_wire_4803)
    );

    bfr new_Jinkela_buffer_4081 (
        .din(new_Jinkela_wire_4779),
        .dout(new_Jinkela_wire_4780)
    );

    bfr new_Jinkela_buffer_4156 (
        .din(n_0079_),
        .dout(new_Jinkela_wire_4875)
    );

    bfr new_Jinkela_buffer_4127 (
        .din(new_Jinkela_wire_4827),
        .dout(new_Jinkela_wire_4828)
    );

    bfr new_Jinkela_buffer_4103 (
        .din(new_Jinkela_wire_4803),
        .dout(new_Jinkela_wire_4804)
    );

    bfr new_Jinkela_buffer_1010 (
        .din(new_Jinkela_wire_1084),
        .dout(new_Jinkela_wire_1085)
    );

    bfr new_Jinkela_buffer_1102 (
        .din(new_Jinkela_wire_1413),
        .dout(new_Jinkela_wire_1414)
    );

    bfr new_Jinkela_buffer_1049 (
        .din(new_Jinkela_wire_1125),
        .dout(new_Jinkela_wire_1126)
    );

    bfr new_Jinkela_buffer_7497 (
        .din(new_Jinkela_wire_9323),
        .dout(new_Jinkela_wire_9324)
    );

    bfr new_Jinkela_buffer_7534 (
        .din(new_Jinkela_wire_9377),
        .dout(new_Jinkela_wire_9378)
    );

    bfr new_Jinkela_buffer_7515 (
        .din(new_Jinkela_wire_9354),
        .dout(new_Jinkela_wire_9355)
    );

    bfr new_Jinkela_buffer_1050 (
        .din(new_Jinkela_wire_1126),
        .dout(new_Jinkela_wire_1127)
    );

    bfr new_Jinkela_buffer_7498 (
        .din(new_Jinkela_wire_9324),
        .dout(new_Jinkela_wire_9325)
    );

    bfr new_Jinkela_buffer_1103 (
        .din(new_Jinkela_wire_1414),
        .dout(new_Jinkela_wire_1415)
    );

    spl4L new_Jinkela_splitter_742 (
        .a(n_1235_),
        .d(new_Jinkela_wire_9381),
        .b(new_Jinkela_wire_9382),
        .e(new_Jinkela_wire_9383),
        .c(new_Jinkela_wire_9384)
    );

    bfr new_Jinkela_buffer_1293 (
        .din(N296),
        .dout(new_Jinkela_wire_1614)
    );

    bfr new_Jinkela_buffer_1051 (
        .din(new_Jinkela_wire_1127),
        .dout(new_Jinkela_wire_1128)
    );

    bfr new_Jinkela_buffer_7499 (
        .din(new_Jinkela_wire_9325),
        .dout(new_Jinkela_wire_9326)
    );

    bfr new_Jinkela_buffer_7531 (
        .din(new_Jinkela_wire_9372),
        .dout(new_Jinkela_wire_9373)
    );

    bfr new_Jinkela_buffer_7516 (
        .din(new_Jinkela_wire_9355),
        .dout(new_Jinkela_wire_9356)
    );

    bfr new_Jinkela_buffer_1052 (
        .din(new_Jinkela_wire_1128),
        .dout(new_Jinkela_wire_1129)
    );

    bfr new_Jinkela_buffer_7500 (
        .din(new_Jinkela_wire_9326),
        .dout(new_Jinkela_wire_9327)
    );

    bfr new_Jinkela_buffer_1104 (
        .din(new_Jinkela_wire_1415),
        .dout(new_Jinkela_wire_1416)
    );

    bfr new_Jinkela_buffer_1225 (
        .din(new_Jinkela_wire_1543),
        .dout(new_Jinkela_wire_1544)
    );

    bfr new_Jinkela_buffer_1053 (
        .din(new_Jinkela_wire_1129),
        .dout(new_Jinkela_wire_1130)
    );

    bfr new_Jinkela_buffer_7501 (
        .din(new_Jinkela_wire_9327),
        .dout(new_Jinkela_wire_9328)
    );

    spl4L new_Jinkela_splitter_50 (
        .a(new_Jinkela_wire_1221),
        .d(new_Jinkela_wire_1222),
        .b(new_Jinkela_wire_1243),
        .e(new_Jinkela_wire_1264),
        .c(new_Jinkela_wire_1285)
    );

    bfr new_Jinkela_buffer_7537 (
        .din(n_1184_),
        .dout(new_Jinkela_wire_9385)
    );

    bfr new_Jinkela_buffer_7517 (
        .din(new_Jinkela_wire_9356),
        .dout(new_Jinkela_wire_9357)
    );

    bfr new_Jinkela_buffer_1054 (
        .din(new_Jinkela_wire_1130),
        .dout(new_Jinkela_wire_1131)
    );

    bfr new_Jinkela_buffer_7502 (
        .din(new_Jinkela_wire_9328),
        .dout(new_Jinkela_wire_9329)
    );

    spl3L new_Jinkela_splitter_36 (
        .a(new_Jinkela_wire_1167),
        .d(new_Jinkela_wire_1168),
        .b(new_Jinkela_wire_1179),
        .c(new_Jinkela_wire_1200)
    );

    bfr new_Jinkela_buffer_1055 (
        .din(new_Jinkela_wire_1131),
        .dout(new_Jinkela_wire_1132)
    );

    bfr new_Jinkela_buffer_7503 (
        .din(new_Jinkela_wire_9329),
        .dout(new_Jinkela_wire_9330)
    );

    spl4L new_Jinkela_splitter_40 (
        .a(new_Jinkela_wire_1179),
        .d(new_Jinkela_wire_1180),
        .b(new_Jinkela_wire_1185),
        .e(new_Jinkela_wire_1190),
        .c(new_Jinkela_wire_1195)
    );

    bfr new_Jinkela_buffer_7532 (
        .din(new_Jinkela_wire_9373),
        .dout(new_Jinkela_wire_9374)
    );

    bfr new_Jinkela_buffer_7518 (
        .din(new_Jinkela_wire_9357),
        .dout(new_Jinkela_wire_9358)
    );

    bfr new_Jinkela_buffer_1056 (
        .din(new_Jinkela_wire_1132),
        .dout(new_Jinkela_wire_1133)
    );

    bfr new_Jinkela_buffer_7504 (
        .din(new_Jinkela_wire_9330),
        .dout(new_Jinkela_wire_9331)
    );

    spl2 new_Jinkela_splitter_37 (
        .a(new_Jinkela_wire_1168),
        .b(new_Jinkela_wire_1169),
        .c(new_Jinkela_wire_1174)
    );

    bfr new_Jinkela_buffer_1057 (
        .din(new_Jinkela_wire_1133),
        .dout(new_Jinkela_wire_1134)
    );

    bfr new_Jinkela_buffer_7505 (
        .din(new_Jinkela_wire_9331),
        .dout(new_Jinkela_wire_9332)
    );

    spl4L new_Jinkela_splitter_39 (
        .a(new_Jinkela_wire_1174),
        .d(new_Jinkela_wire_1175),
        .b(new_Jinkela_wire_1176),
        .e(new_Jinkela_wire_1177),
        .c(new_Jinkela_wire_1178)
    );

    bfr new_Jinkela_buffer_7540 (
        .din(n_0628_),
        .dout(new_Jinkela_wire_9390)
    );

    bfr new_Jinkela_buffer_7519 (
        .din(new_Jinkela_wire_9358),
        .dout(new_Jinkela_wire_9359)
    );

    bfr new_Jinkela_buffer_1058 (
        .din(new_Jinkela_wire_1134),
        .dout(new_Jinkela_wire_1135)
    );

    bfr new_Jinkela_buffer_7506 (
        .din(new_Jinkela_wire_9332),
        .dout(new_Jinkela_wire_9333)
    );

    spl4L new_Jinkela_splitter_38 (
        .a(new_Jinkela_wire_1169),
        .d(new_Jinkela_wire_1170),
        .b(new_Jinkela_wire_1171),
        .e(new_Jinkela_wire_1172),
        .c(new_Jinkela_wire_1173)
    );

    bfr new_Jinkela_buffer_1059 (
        .din(new_Jinkela_wire_1135),
        .dout(new_Jinkela_wire_1136)
    );

    bfr new_Jinkela_buffer_7507 (
        .din(new_Jinkela_wire_9333),
        .dout(new_Jinkela_wire_9334)
    );

    spl4L new_Jinkela_splitter_41 (
        .a(new_Jinkela_wire_1180),
        .d(new_Jinkela_wire_1181),
        .b(new_Jinkela_wire_1182),
        .e(new_Jinkela_wire_1183),
        .c(new_Jinkela_wire_1184)
    );

    bfr new_Jinkela_buffer_7535 (
        .din(new_Jinkela_wire_9378),
        .dout(new_Jinkela_wire_9379)
    );

    bfr new_Jinkela_buffer_7520 (
        .din(new_Jinkela_wire_9359),
        .dout(new_Jinkela_wire_9360)
    );

    bfr new_Jinkela_buffer_1060 (
        .din(new_Jinkela_wire_1136),
        .dout(new_Jinkela_wire_1137)
    );

    bfr new_Jinkela_buffer_7508 (
        .din(new_Jinkela_wire_9334),
        .dout(new_Jinkela_wire_9335)
    );

    spl4L new_Jinkela_splitter_45 (
        .a(new_Jinkela_wire_1200),
        .d(new_Jinkela_wire_1201),
        .b(new_Jinkela_wire_1206),
        .e(new_Jinkela_wire_1211),
        .c(new_Jinkela_wire_1216)
    );

    bfr new_Jinkela_buffer_1061 (
        .din(new_Jinkela_wire_1137),
        .dout(new_Jinkela_wire_1138)
    );

    spl2 new_Jinkela_splitter_744 (
        .a(n_0826_),
        .b(new_Jinkela_wire_9392),
        .c(new_Jinkela_wire_9393)
    );

    bfr new_Jinkela_buffer_7521 (
        .din(new_Jinkela_wire_9360),
        .dout(new_Jinkela_wire_9361)
    );

    spl4L new_Jinkela_splitter_42 (
        .a(new_Jinkela_wire_1185),
        .d(new_Jinkela_wire_1186),
        .b(new_Jinkela_wire_1187),
        .e(new_Jinkela_wire_1188),
        .c(new_Jinkela_wire_1189)
    );

    bfr new_Jinkela_buffer_7539 (
        .din(new_Jinkela_wire_9386),
        .dout(new_Jinkela_wire_9387)
    );

    bfr new_Jinkela_buffer_1062 (
        .din(new_Jinkela_wire_1138),
        .dout(new_Jinkela_wire_1139)
    );

    bfr new_Jinkela_buffer_7536 (
        .din(new_Jinkela_wire_9379),
        .dout(new_Jinkela_wire_9380)
    );

    bfr new_Jinkela_buffer_7522 (
        .din(new_Jinkela_wire_9361),
        .dout(new_Jinkela_wire_9362)
    );

    spl4L new_Jinkela_splitter_46 (
        .a(new_Jinkela_wire_1201),
        .d(new_Jinkela_wire_1202),
        .b(new_Jinkela_wire_1203),
        .e(new_Jinkela_wire_1204),
        .c(new_Jinkela_wire_1205)
    );

    bfr new_Jinkela_buffer_1063 (
        .din(new_Jinkela_wire_1139),
        .dout(new_Jinkela_wire_1140)
    );

    bfr new_Jinkela_buffer_7523 (
        .din(new_Jinkela_wire_9362),
        .dout(new_Jinkela_wire_9363)
    );

    spl4L new_Jinkela_splitter_43 (
        .a(new_Jinkela_wire_1190),
        .d(new_Jinkela_wire_1191),
        .b(new_Jinkela_wire_1192),
        .e(new_Jinkela_wire_1193),
        .c(new_Jinkela_wire_1194)
    );

    bfr new_Jinkela_buffer_7538 (
        .din(n_0792_),
        .dout(new_Jinkela_wire_9386)
    );

    bfr new_Jinkela_buffer_1064 (
        .din(new_Jinkela_wire_1140),
        .dout(new_Jinkela_wire_1141)
    );

    bfr new_Jinkela_buffer_7524 (
        .din(new_Jinkela_wire_9363),
        .dout(new_Jinkela_wire_9364)
    );

    spl4L new_Jinkela_splitter_44 (
        .a(new_Jinkela_wire_1195),
        .d(new_Jinkela_wire_1196),
        .b(new_Jinkela_wire_1197),
        .e(new_Jinkela_wire_1198),
        .c(new_Jinkela_wire_1199)
    );

    bfr new_Jinkela_buffer_1065 (
        .din(new_Jinkela_wire_1141),
        .dout(new_Jinkela_wire_1142)
    );

    bfr new_Jinkela_buffer_7525 (
        .din(new_Jinkela_wire_9364),
        .dout(new_Jinkela_wire_9365)
    );

    spl4L new_Jinkela_splitter_71 (
        .a(new_Jinkela_wire_1306),
        .d(new_Jinkela_wire_1307),
        .b(new_Jinkela_wire_1328),
        .e(new_Jinkela_wire_1349),
        .c(new_Jinkela_wire_1370)
    );

    bfr new_Jinkela_buffer_7542 (
        .din(n_1179_),
        .dout(new_Jinkela_wire_9394)
    );

    bfr new_Jinkela_buffer_1066 (
        .din(new_Jinkela_wire_1142),
        .dout(new_Jinkela_wire_1143)
    );

    bfr new_Jinkela_buffer_7541 (
        .din(new_Jinkela_wire_9390),
        .dout(new_Jinkela_wire_9391)
    );

    spl2 new_Jinkela_splitter_743 (
        .a(new_Jinkela_wire_9387),
        .b(new_Jinkela_wire_9388),
        .c(new_Jinkela_wire_9389)
    );

    spl4L new_Jinkela_splitter_47 (
        .a(new_Jinkela_wire_1206),
        .d(new_Jinkela_wire_1207),
        .b(new_Jinkela_wire_1208),
        .e(new_Jinkela_wire_1209),
        .c(new_Jinkela_wire_1210)
    );

    bfr new_Jinkela_buffer_1067 (
        .din(new_Jinkela_wire_1143),
        .dout(new_Jinkela_wire_1144)
    );

    spl4L new_Jinkela_splitter_49 (
        .a(new_Jinkela_wire_1216),
        .d(new_Jinkela_wire_1217),
        .b(new_Jinkela_wire_1218),
        .e(new_Jinkela_wire_1219),
        .c(new_Jinkela_wire_1220)
    );

    bfr new_Jinkela_buffer_1068 (
        .din(new_Jinkela_wire_1144),
        .dout(new_Jinkela_wire_1145)
    );

    spl2 new_Jinkela_splitter_745 (
        .a(n_1324_),
        .b(new_Jinkela_wire_9395),
        .c(new_Jinkela_wire_9396)
    );

    bfr new_Jinkela_buffer_7543 (
        .din(n_0066_),
        .dout(new_Jinkela_wire_9401)
    );

    spl4L new_Jinkela_splitter_48 (
        .a(new_Jinkela_wire_1211),
        .d(new_Jinkela_wire_1212),
        .b(new_Jinkela_wire_1213),
        .e(new_Jinkela_wire_1214),
        .c(new_Jinkela_wire_1215)
    );

    spl2 new_Jinkela_splitter_746 (
        .a(new_Jinkela_wire_9396),
        .b(new_Jinkela_wire_9397),
        .c(new_Jinkela_wire_9398)
    );

    bfr new_Jinkela_buffer_1069 (
        .din(new_Jinkela_wire_1145),
        .dout(new_Jinkela_wire_1146)
    );

    bfr new_Jinkela_buffer_7551 (
        .din(new_net_2497),
        .dout(new_Jinkela_wire_9411)
    );

    spl2 new_Jinkela_splitter_173 (
        .a(new_Jinkela_wire_3775),
        .b(new_Jinkela_wire_3776),
        .c(new_Jinkela_wire_3777)
    );

    bfr new_Jinkela_buffer_3210 (
        .din(new_Jinkela_wire_3664),
        .dout(new_Jinkela_wire_3665)
    );

    bfr new_Jinkela_buffer_3253 (
        .din(new_Jinkela_wire_3741),
        .dout(new_Jinkela_wire_3742)
    );

    bfr new_Jinkela_buffer_3211 (
        .din(new_Jinkela_wire_3665),
        .dout(new_Jinkela_wire_3666)
    );

    bfr new_Jinkela_buffer_3252 (
        .din(new_Jinkela_wire_3740),
        .dout(new_Jinkela_wire_3741)
    );

    bfr new_Jinkela_buffer_3212 (
        .din(new_Jinkela_wire_3666),
        .dout(new_Jinkela_wire_3667)
    );

    bfr new_Jinkela_buffer_3280 (
        .din(new_Jinkela_wire_3784),
        .dout(new_Jinkela_wire_3785)
    );

    bfr new_Jinkela_buffer_3213 (
        .din(new_Jinkela_wire_3667),
        .dout(new_Jinkela_wire_3668)
    );

    spl4L new_Jinkela_splitter_176 (
        .a(n_1314_),
        .d(new_Jinkela_wire_3791),
        .b(new_Jinkela_wire_3792),
        .e(new_Jinkela_wire_3793),
        .c(new_Jinkela_wire_3794)
    );

    bfr new_Jinkela_buffer_3254 (
        .din(new_Jinkela_wire_3742),
        .dout(new_Jinkela_wire_3743)
    );

    bfr new_Jinkela_buffer_3214 (
        .din(new_Jinkela_wire_3668),
        .dout(new_Jinkela_wire_3669)
    );

    bfr new_Jinkela_buffer_3215 (
        .din(new_Jinkela_wire_3669),
        .dout(new_Jinkela_wire_3670)
    );

    bfr new_Jinkela_buffer_3313 (
        .din(n_0600_),
        .dout(new_Jinkela_wire_3822)
    );

    bfr new_Jinkela_buffer_3255 (
        .din(new_Jinkela_wire_3743),
        .dout(new_Jinkela_wire_3744)
    );

    bfr new_Jinkela_buffer_3216 (
        .din(new_Jinkela_wire_3670),
        .dout(new_Jinkela_wire_3671)
    );

    bfr new_Jinkela_buffer_3283 (
        .din(new_Jinkela_wire_3787),
        .dout(new_Jinkela_wire_3788)
    );

    bfr new_Jinkela_buffer_3217 (
        .din(new_Jinkela_wire_3671),
        .dout(new_Jinkela_wire_3672)
    );

    bfr new_Jinkela_buffer_3281 (
        .din(new_Jinkela_wire_3785),
        .dout(new_Jinkela_wire_3786)
    );

    bfr new_Jinkela_buffer_3256 (
        .din(new_Jinkela_wire_3744),
        .dout(new_Jinkela_wire_3745)
    );

    bfr new_Jinkela_buffer_3218 (
        .din(new_Jinkela_wire_3672),
        .dout(new_Jinkela_wire_3673)
    );

    bfr new_Jinkela_buffer_3219 (
        .din(new_Jinkela_wire_3673),
        .dout(new_Jinkela_wire_3674)
    );

    bfr new_Jinkela_buffer_3257 (
        .din(new_Jinkela_wire_3745),
        .dout(new_Jinkela_wire_3746)
    );

    bfr new_Jinkela_buffer_3286 (
        .din(new_Jinkela_wire_3794),
        .dout(new_Jinkela_wire_3795)
    );

    bfr new_Jinkela_buffer_3258 (
        .din(new_Jinkela_wire_3746),
        .dout(new_Jinkela_wire_3747)
    );

    bfr new_Jinkela_buffer_3284 (
        .din(new_Jinkela_wire_3788),
        .dout(new_Jinkela_wire_3789)
    );

    bfr new_Jinkela_buffer_3259 (
        .din(new_Jinkela_wire_3747),
        .dout(new_Jinkela_wire_3748)
    );

    bfr new_Jinkela_buffer_3326 (
        .din(n_0478_),
        .dout(new_Jinkela_wire_3835)
    );

    bfr new_Jinkela_buffer_3260 (
        .din(new_Jinkela_wire_3748),
        .dout(new_Jinkela_wire_3749)
    );

    bfr new_Jinkela_buffer_3285 (
        .din(new_Jinkela_wire_3789),
        .dout(new_Jinkela_wire_3790)
    );

    bfr new_Jinkela_buffer_3261 (
        .din(new_Jinkela_wire_3749),
        .dout(new_Jinkela_wire_3750)
    );

    bfr new_Jinkela_buffer_3314 (
        .din(n_0331_),
        .dout(new_Jinkela_wire_3823)
    );

    bfr new_Jinkela_buffer_3262 (
        .din(new_Jinkela_wire_3750),
        .dout(new_Jinkela_wire_3751)
    );

    bfr new_Jinkela_buffer_3287 (
        .din(new_Jinkela_wire_3795),
        .dout(new_Jinkela_wire_3796)
    );

    bfr new_Jinkela_buffer_3263 (
        .din(new_Jinkela_wire_3751),
        .dout(new_Jinkela_wire_3752)
    );

    bfr new_Jinkela_buffer_3264 (
        .din(new_Jinkela_wire_3752),
        .dout(new_Jinkela_wire_3753)
    );

    bfr new_Jinkela_buffer_3315 (
        .din(new_Jinkela_wire_3823),
        .dout(new_Jinkela_wire_3824)
    );

    bfr new_Jinkela_buffer_3288 (
        .din(new_Jinkela_wire_3796),
        .dout(new_Jinkela_wire_3797)
    );

    bfr new_Jinkela_buffer_3265 (
        .din(new_Jinkela_wire_3753),
        .dout(new_Jinkela_wire_3754)
    );

    bfr new_Jinkela_buffer_3266 (
        .din(new_Jinkela_wire_3754),
        .dout(new_Jinkela_wire_3755)
    );

    spl2 new_Jinkela_splitter_177 (
        .a(n_0877_),
        .b(new_Jinkela_wire_3836),
        .c(new_Jinkela_wire_3837)
    );

    bfr new_Jinkela_buffer_3289 (
        .din(new_Jinkela_wire_3797),
        .dout(new_Jinkela_wire_3798)
    );

    bfr new_Jinkela_buffer_3267 (
        .din(new_Jinkela_wire_3755),
        .dout(new_Jinkela_wire_3756)
    );

    bfr new_Jinkela_buffer_2362 (
        .din(new_Jinkela_wire_2758),
        .dout(new_Jinkela_wire_2759)
    );

    spl2 new_Jinkela_splitter_585 (
        .a(new_Jinkela_wire_8088),
        .b(new_Jinkela_wire_8089),
        .c(new_Jinkela_wire_8090)
    );

    bfr new_Jinkela_buffer_2319 (
        .din(new_Jinkela_wire_2710),
        .dout(new_Jinkela_wire_2711)
    );

    bfr new_Jinkela_buffer_6561 (
        .din(new_Jinkela_wire_8027),
        .dout(new_Jinkela_wire_8028)
    );

    bfr new_Jinkela_buffer_2486 (
        .din(new_Jinkela_wire_2887),
        .dout(new_Jinkela_wire_2888)
    );

    bfr new_Jinkela_buffer_6613 (
        .din(new_Jinkela_wire_8094),
        .dout(new_Jinkela_wire_8095)
    );

    bfr new_Jinkela_buffer_2320 (
        .din(new_Jinkela_wire_2711),
        .dout(new_Jinkela_wire_2712)
    );

    bfr new_Jinkela_buffer_6562 (
        .din(new_Jinkela_wire_8028),
        .dout(new_Jinkela_wire_8029)
    );

    bfr new_Jinkela_buffer_2363 (
        .din(new_Jinkela_wire_2759),
        .dout(new_Jinkela_wire_2760)
    );

    spl2 new_Jinkela_splitter_589 (
        .a(n_0167_),
        .b(new_Jinkela_wire_8104),
        .c(new_Jinkela_wire_8105)
    );

    bfr new_Jinkela_buffer_2321 (
        .din(new_Jinkela_wire_2712),
        .dout(new_Jinkela_wire_2713)
    );

    bfr new_Jinkela_buffer_6616 (
        .din(new_Jinkela_wire_8097),
        .dout(new_Jinkela_wire_8098)
    );

    bfr new_Jinkela_buffer_6563 (
        .din(new_Jinkela_wire_8029),
        .dout(new_Jinkela_wire_8030)
    );

    bfr new_Jinkela_buffer_2489 (
        .din(new_Jinkela_wire_2890),
        .dout(new_Jinkela_wire_2891)
    );

    bfr new_Jinkela_buffer_2322 (
        .din(new_Jinkela_wire_2713),
        .dout(new_Jinkela_wire_2714)
    );

    spl2 new_Jinkela_splitter_588 (
        .a(n_1218_),
        .b(new_Jinkela_wire_8102),
        .c(new_Jinkela_wire_8103)
    );

    bfr new_Jinkela_buffer_6564 (
        .din(new_Jinkela_wire_8030),
        .dout(new_Jinkela_wire_8031)
    );

    bfr new_Jinkela_buffer_2364 (
        .din(new_Jinkela_wire_2760),
        .dout(new_Jinkela_wire_2761)
    );

    bfr new_Jinkela_buffer_6614 (
        .din(new_Jinkela_wire_8095),
        .dout(new_Jinkela_wire_8096)
    );

    bfr new_Jinkela_buffer_2323 (
        .din(new_Jinkela_wire_2714),
        .dout(new_Jinkela_wire_2715)
    );

    bfr new_Jinkela_buffer_6565 (
        .din(new_Jinkela_wire_8031),
        .dout(new_Jinkela_wire_8032)
    );

    bfr new_Jinkela_buffer_2424 (
        .din(new_Jinkela_wire_2822),
        .dout(new_Jinkela_wire_2823)
    );

    bfr new_Jinkela_buffer_2324 (
        .din(new_Jinkela_wire_2715),
        .dout(new_Jinkela_wire_2716)
    );

    bfr new_Jinkela_buffer_6566 (
        .din(new_Jinkela_wire_8032),
        .dout(new_Jinkela_wire_8033)
    );

    bfr new_Jinkela_buffer_2365 (
        .din(new_Jinkela_wire_2761),
        .dout(new_Jinkela_wire_2762)
    );

    bfr new_Jinkela_buffer_2325 (
        .din(new_Jinkela_wire_2716),
        .dout(new_Jinkela_wire_2717)
    );

    bfr new_Jinkela_buffer_6617 (
        .din(new_Jinkela_wire_8098),
        .dout(new_Jinkela_wire_8099)
    );

    bfr new_Jinkela_buffer_6567 (
        .din(new_Jinkela_wire_8033),
        .dout(new_Jinkela_wire_8034)
    );

    bfr new_Jinkela_buffer_2487 (
        .din(new_Jinkela_wire_2888),
        .dout(new_Jinkela_wire_2889)
    );

    bfr new_Jinkela_buffer_2326 (
        .din(new_Jinkela_wire_2717),
        .dout(new_Jinkela_wire_2718)
    );

    bfr new_Jinkela_buffer_6568 (
        .din(new_Jinkela_wire_8034),
        .dout(new_Jinkela_wire_8035)
    );

    bfr new_Jinkela_buffer_2366 (
        .din(new_Jinkela_wire_2762),
        .dout(new_Jinkela_wire_2763)
    );

    spl3L new_Jinkela_splitter_592 (
        .a(n_1042_),
        .d(new_Jinkela_wire_8165),
        .b(new_Jinkela_wire_8166),
        .c(new_Jinkela_wire_8167)
    );

    bfr new_Jinkela_buffer_2327 (
        .din(new_Jinkela_wire_2718),
        .dout(new_Jinkela_wire_2719)
    );

    bfr new_Jinkela_buffer_6618 (
        .din(new_Jinkela_wire_8099),
        .dout(new_Jinkela_wire_8100)
    );

    bfr new_Jinkela_buffer_6569 (
        .din(new_Jinkela_wire_8035),
        .dout(new_Jinkela_wire_8036)
    );

    bfr new_Jinkela_buffer_2425 (
        .din(new_Jinkela_wire_2823),
        .dout(new_Jinkela_wire_2824)
    );

    bfr new_Jinkela_buffer_2328 (
        .din(new_Jinkela_wire_2719),
        .dout(new_Jinkela_wire_2720)
    );

    spl2 new_Jinkela_splitter_591 (
        .a(n_0538_),
        .b(new_Jinkela_wire_8163),
        .c(new_Jinkela_wire_8164)
    );

    bfr new_Jinkela_buffer_6570 (
        .din(new_Jinkela_wire_8036),
        .dout(new_Jinkela_wire_8037)
    );

    bfr new_Jinkela_buffer_2367 (
        .din(new_Jinkela_wire_2763),
        .dout(new_Jinkela_wire_2764)
    );

    spl2 new_Jinkela_splitter_595 (
        .a(n_0787_),
        .b(new_Jinkela_wire_8173),
        .c(new_Jinkela_wire_8174)
    );

    bfr new_Jinkela_buffer_2329 (
        .din(new_Jinkela_wire_2720),
        .dout(new_Jinkela_wire_2721)
    );

    bfr new_Jinkela_buffer_6619 (
        .din(new_Jinkela_wire_8100),
        .dout(new_Jinkela_wire_8101)
    );

    bfr new_Jinkela_buffer_6571 (
        .din(new_Jinkela_wire_8037),
        .dout(new_Jinkela_wire_8038)
    );

    bfr new_Jinkela_buffer_2496 (
        .din(N220),
        .dout(new_Jinkela_wire_2898)
    );

    bfr new_Jinkela_buffer_2330 (
        .din(new_Jinkela_wire_2721),
        .dout(new_Jinkela_wire_2722)
    );

    bfr new_Jinkela_buffer_6620 (
        .din(new_Jinkela_wire_8105),
        .dout(new_Jinkela_wire_8106)
    );

    bfr new_Jinkela_buffer_6572 (
        .din(new_Jinkela_wire_8038),
        .dout(new_Jinkela_wire_8039)
    );

    bfr new_Jinkela_buffer_2368 (
        .din(new_Jinkela_wire_2764),
        .dout(new_Jinkela_wire_2765)
    );

    bfr new_Jinkela_buffer_2331 (
        .din(new_Jinkela_wire_2722),
        .dout(new_Jinkela_wire_2723)
    );

    bfr new_Jinkela_buffer_6573 (
        .din(new_Jinkela_wire_8039),
        .dout(new_Jinkela_wire_8040)
    );

    spl3L new_Jinkela_splitter_134 (
        .a(new_Jinkela_wire_2824),
        .d(new_Jinkela_wire_2825),
        .b(new_Jinkela_wire_2826),
        .c(new_Jinkela_wire_2827)
    );

    spl3L new_Jinkela_splitter_594 (
        .a(n_0697_),
        .d(new_Jinkela_wire_8170),
        .b(new_Jinkela_wire_8171),
        .c(new_Jinkela_wire_8172)
    );

    bfr new_Jinkela_buffer_2332 (
        .din(new_Jinkela_wire_2723),
        .dout(new_Jinkela_wire_2724)
    );

    bfr new_Jinkela_buffer_6621 (
        .din(new_Jinkela_wire_8106),
        .dout(new_Jinkela_wire_8107)
    );

    bfr new_Jinkela_buffer_6574 (
        .din(new_Jinkela_wire_8040),
        .dout(new_Jinkela_wire_8041)
    );

    bfr new_Jinkela_buffer_2369 (
        .din(new_Jinkela_wire_2765),
        .dout(new_Jinkela_wire_2766)
    );

    bfr new_Jinkela_buffer_2333 (
        .din(new_Jinkela_wire_2724),
        .dout(new_Jinkela_wire_2725)
    );

    bfr new_Jinkela_buffer_6575 (
        .din(new_Jinkela_wire_8041),
        .dout(new_Jinkela_wire_8042)
    );

    bfr new_Jinkela_buffer_2490 (
        .din(new_Jinkela_wire_2891),
        .dout(new_Jinkela_wire_2892)
    );

    bfr new_Jinkela_buffer_2334 (
        .din(new_Jinkela_wire_2725),
        .dout(new_Jinkela_wire_2726)
    );

    bfr new_Jinkela_buffer_6622 (
        .din(new_Jinkela_wire_8107),
        .dout(new_Jinkela_wire_8108)
    );

    bfr new_Jinkela_buffer_6576 (
        .din(new_Jinkela_wire_8042),
        .dout(new_Jinkela_wire_8043)
    );

    bfr new_Jinkela_buffer_2370 (
        .din(new_Jinkela_wire_2766),
        .dout(new_Jinkela_wire_2767)
    );

    bfr new_Jinkela_buffer_2335 (
        .din(new_Jinkela_wire_2726),
        .dout(new_Jinkela_wire_2727)
    );

    spl2 new_Jinkela_splitter_593 (
        .a(new_Jinkela_wire_8167),
        .b(new_Jinkela_wire_8168),
        .c(new_Jinkela_wire_8169)
    );

    bfr new_Jinkela_buffer_6577 (
        .din(new_Jinkela_wire_8043),
        .dout(new_Jinkela_wire_8044)
    );

    bfr new_Jinkela_buffer_2426 (
        .din(new_Jinkela_wire_2827),
        .dout(new_Jinkela_wire_2828)
    );

    spl2 new_Jinkela_splitter_596 (
        .a(n_0602_),
        .b(new_Jinkela_wire_8175),
        .c(new_Jinkela_wire_8176)
    );

    bfr new_Jinkela_buffer_2336 (
        .din(new_Jinkela_wire_2727),
        .dout(new_Jinkela_wire_2728)
    );

    bfr new_Jinkela_buffer_6623 (
        .din(new_Jinkela_wire_8108),
        .dout(new_Jinkela_wire_8109)
    );

    bfr new_Jinkela_buffer_6578 (
        .din(new_Jinkela_wire_8044),
        .dout(new_Jinkela_wire_8045)
    );

    bfr new_Jinkela_buffer_2371 (
        .din(new_Jinkela_wire_2767),
        .dout(new_Jinkela_wire_2768)
    );

    bfr new_Jinkela_buffer_2337 (
        .din(new_Jinkela_wire_2728),
        .dout(new_Jinkela_wire_2729)
    );

    bfr new_Jinkela_buffer_6579 (
        .din(new_Jinkela_wire_8045),
        .dout(new_Jinkela_wire_8046)
    );

    bfr new_Jinkela_buffer_2493 (
        .din(new_Jinkela_wire_2894),
        .dout(new_Jinkela_wire_2895)
    );

    bfr new_Jinkela_buffer_2338 (
        .din(new_Jinkela_wire_2729),
        .dout(new_Jinkela_wire_2730)
    );

    bfr new_Jinkela_buffer_6624 (
        .din(new_Jinkela_wire_8109),
        .dout(new_Jinkela_wire_8110)
    );

    bfr new_Jinkela_buffer_6580 (
        .din(new_Jinkela_wire_8046),
        .dout(new_Jinkela_wire_8047)
    );

    bfr new_Jinkela_buffer_2372 (
        .din(new_Jinkela_wire_2768),
        .dout(new_Jinkela_wire_2769)
    );

    bfr new_Jinkela_buffer_2339 (
        .din(new_Jinkela_wire_2730),
        .dout(new_Jinkela_wire_2731)
    );

    spl2 new_Jinkela_splitter_597 (
        .a(n_0100_),
        .b(new_Jinkela_wire_8177),
        .c(new_Jinkela_wire_8178)
    );

    bfr new_Jinkela_buffer_6581 (
        .din(new_Jinkela_wire_8047),
        .dout(new_Jinkela_wire_8048)
    );

    bfr new_Jinkela_buffer_7 (
        .din(new_Jinkela_wire_8),
        .dout(new_Jinkela_wire_9)
    );

    spl2 new_Jinkela_splitter_749 (
        .a(n_0015_),
        .b(new_Jinkela_wire_9417),
        .c(new_Jinkela_wire_9421)
    );

    bfr new_Jinkela_buffer_70 (
        .din(new_Jinkela_wire_77),
        .dout(new_Jinkela_wire_78)
    );

    spl2 new_Jinkela_splitter_747 (
        .a(new_Jinkela_wire_9398),
        .b(new_Jinkela_wire_9399),
        .c(new_Jinkela_wire_9400)
    );

    bfr new_Jinkela_buffer_8 (
        .din(new_Jinkela_wire_9),
        .dout(new_Jinkela_wire_10)
    );

    bfr new_Jinkela_buffer_7544 (
        .din(new_Jinkela_wire_9401),
        .dout(new_Jinkela_wire_9402)
    );

    bfr new_Jinkela_buffer_73 (
        .din(new_Jinkela_wire_80),
        .dout(new_Jinkela_wire_81)
    );

    bfr new_Jinkela_buffer_7545 (
        .din(new_Jinkela_wire_9402),
        .dout(new_Jinkela_wire_9403)
    );

    bfr new_Jinkela_buffer_9 (
        .din(new_Jinkela_wire_10),
        .dout(new_Jinkela_wire_11)
    );

    bfr new_Jinkela_buffer_7552 (
        .din(new_Jinkela_wire_9411),
        .dout(new_Jinkela_wire_9412)
    );

    bfr new_Jinkela_buffer_71 (
        .din(new_Jinkela_wire_78),
        .dout(new_Jinkela_wire_79)
    );

    spl4L new_Jinkela_splitter_751 (
        .a(new_Jinkela_wire_9421),
        .d(new_Jinkela_wire_9422),
        .b(new_Jinkela_wire_9423),
        .e(new_Jinkela_wire_9424),
        .c(new_Jinkela_wire_9425)
    );

    bfr new_Jinkela_buffer_10 (
        .din(new_Jinkela_wire_11),
        .dout(new_Jinkela_wire_12)
    );

    bfr new_Jinkela_buffer_7546 (
        .din(new_Jinkela_wire_9403),
        .dout(new_Jinkela_wire_9404)
    );

    bfr new_Jinkela_buffer_80 (
        .din(N180),
        .dout(new_Jinkela_wire_88)
    );

    bfr new_Jinkela_buffer_7553 (
        .din(new_Jinkela_wire_9412),
        .dout(new_Jinkela_wire_9413)
    );

    bfr new_Jinkela_buffer_11 (
        .din(new_Jinkela_wire_12),
        .dout(new_Jinkela_wire_13)
    );

    bfr new_Jinkela_buffer_7547 (
        .din(new_Jinkela_wire_9404),
        .dout(new_Jinkela_wire_9405)
    );

    bfr new_Jinkela_buffer_74 (
        .din(new_Jinkela_wire_81),
        .dout(new_Jinkela_wire_82)
    );

    spl4L new_Jinkela_splitter_754 (
        .a(new_Jinkela_wire_9430),
        .d(new_Jinkela_wire_9431),
        .b(new_Jinkela_wire_9432),
        .e(new_Jinkela_wire_9433),
        .c(new_Jinkela_wire_9434)
    );

    bfr new_Jinkela_buffer_12 (
        .din(new_Jinkela_wire_13),
        .dout(new_Jinkela_wire_14)
    );

    bfr new_Jinkela_buffer_7548 (
        .din(new_Jinkela_wire_9405),
        .dout(new_Jinkela_wire_9406)
    );

    bfr new_Jinkela_buffer_77 (
        .din(new_Jinkela_wire_84),
        .dout(new_Jinkela_wire_85)
    );

    bfr new_Jinkela_buffer_7554 (
        .din(new_Jinkela_wire_9413),
        .dout(new_Jinkela_wire_9414)
    );

    bfr new_Jinkela_buffer_13 (
        .din(new_Jinkela_wire_14),
        .dout(new_Jinkela_wire_15)
    );

    bfr new_Jinkela_buffer_7549 (
        .din(new_Jinkela_wire_9406),
        .dout(new_Jinkela_wire_9407)
    );

    bfr new_Jinkela_buffer_75 (
        .din(new_Jinkela_wire_82),
        .dout(new_Jinkela_wire_83)
    );

    spl2 new_Jinkela_splitter_752 (
        .a(n_0005_),
        .b(new_Jinkela_wire_9426),
        .c(new_Jinkela_wire_9430)
    );

    bfr new_Jinkela_buffer_14 (
        .din(new_Jinkela_wire_15),
        .dout(new_Jinkela_wire_16)
    );

    spl2 new_Jinkela_splitter_748 (
        .a(new_Jinkela_wire_9407),
        .b(new_Jinkela_wire_9408),
        .c(new_Jinkela_wire_9409)
    );

    bfr new_Jinkela_buffer_84 (
        .din(N55),
        .dout(new_Jinkela_wire_92)
    );

    bfr new_Jinkela_buffer_7550 (
        .din(new_Jinkela_wire_9409),
        .dout(new_Jinkela_wire_9410)
    );

    bfr new_Jinkela_buffer_15 (
        .din(new_Jinkela_wire_16),
        .dout(new_Jinkela_wire_17)
    );

    bfr new_Jinkela_buffer_7555 (
        .din(new_Jinkela_wire_9414),
        .dout(new_Jinkela_wire_9415)
    );

    bfr new_Jinkela_buffer_78 (
        .din(new_Jinkela_wire_85),
        .dout(new_Jinkela_wire_86)
    );

    bfr new_Jinkela_buffer_7560 (
        .din(n_0537_),
        .dout(new_Jinkela_wire_9476)
    );

    bfr new_Jinkela_buffer_16 (
        .din(new_Jinkela_wire_17),
        .dout(new_Jinkela_wire_18)
    );

    bfr new_Jinkela_buffer_7556 (
        .din(new_Jinkela_wire_9415),
        .dout(new_Jinkela_wire_9416)
    );

    bfr new_Jinkela_buffer_81 (
        .din(new_Jinkela_wire_88),
        .dout(new_Jinkela_wire_89)
    );

    spl3L new_Jinkela_splitter_750 (
        .a(new_Jinkela_wire_9417),
        .d(new_Jinkela_wire_9418),
        .b(new_Jinkela_wire_9419),
        .c(new_Jinkela_wire_9420)
    );

    bfr new_Jinkela_buffer_17 (
        .din(new_Jinkela_wire_18),
        .dout(new_Jinkela_wire_19)
    );

    spl3L new_Jinkela_splitter_765 (
        .a(n_1209_),
        .d(new_Jinkela_wire_9473),
        .b(new_Jinkela_wire_9474),
        .c(new_Jinkela_wire_9475)
    );

    bfr new_Jinkela_buffer_79 (
        .din(new_Jinkela_wire_86),
        .dout(new_Jinkela_wire_87)
    );

    bfr new_Jinkela_buffer_18 (
        .din(new_Jinkela_wire_19),
        .dout(new_Jinkela_wire_20)
    );

    bfr new_Jinkela_buffer_7557 (
        .din(n_0718_),
        .dout(new_Jinkela_wire_9435)
    );

    spl3L new_Jinkela_splitter_753 (
        .a(new_Jinkela_wire_9426),
        .d(new_Jinkela_wire_9427),
        .b(new_Jinkela_wire_9428),
        .c(new_Jinkela_wire_9429)
    );

    bfr new_Jinkela_buffer_88 (
        .din(N57),
        .dout(new_Jinkela_wire_96)
    );

    spl2 new_Jinkela_splitter_766 (
        .a(n_0511_),
        .b(new_Jinkela_wire_9480),
        .c(new_Jinkela_wire_9481)
    );

    bfr new_Jinkela_buffer_7564 (
        .din(n_0582_),
        .dout(new_Jinkela_wire_9482)
    );

    bfr new_Jinkela_buffer_19 (
        .din(new_Jinkela_wire_20),
        .dout(new_Jinkela_wire_21)
    );

    bfr new_Jinkela_buffer_7561 (
        .din(new_Jinkela_wire_9476),
        .dout(new_Jinkela_wire_9477)
    );

    bfr new_Jinkela_buffer_82 (
        .din(new_Jinkela_wire_89),
        .dout(new_Jinkela_wire_90)
    );

    bfr new_Jinkela_buffer_7559 (
        .din(n_0235_),
        .dout(new_Jinkela_wire_9468)
    );

    bfr new_Jinkela_buffer_20 (
        .din(new_Jinkela_wire_21),
        .dout(new_Jinkela_wire_22)
    );

    spl4L new_Jinkela_splitter_764 (
        .a(n_0887_),
        .d(new_Jinkela_wire_9469),
        .b(new_Jinkela_wire_9470),
        .e(new_Jinkela_wire_9471),
        .c(new_Jinkela_wire_9472)
    );

    bfr new_Jinkela_buffer_85 (
        .din(new_Jinkela_wire_92),
        .dout(new_Jinkela_wire_93)
    );

    spl2 new_Jinkela_splitter_755 (
        .a(new_Jinkela_wire_9436),
        .b(new_Jinkela_wire_9437),
        .c(new_Jinkela_wire_9445)
    );

    bfr new_Jinkela_buffer_21 (
        .din(new_Jinkela_wire_22),
        .dout(new_Jinkela_wire_23)
    );

    spl4L new_Jinkela_splitter_758 (
        .a(new_Jinkela_wire_9445),
        .d(new_Jinkela_wire_9446),
        .b(new_Jinkela_wire_9451),
        .e(new_Jinkela_wire_9456),
        .c(new_Jinkela_wire_9461)
    );

    bfr new_Jinkela_buffer_83 (
        .din(new_Jinkela_wire_90),
        .dout(new_Jinkela_wire_91)
    );

    bfr new_Jinkela_buffer_22 (
        .din(new_Jinkela_wire_23),
        .dout(new_Jinkela_wire_24)
    );

    bfr new_Jinkela_buffer_7558 (
        .din(new_Jinkela_wire_9435),
        .dout(new_Jinkela_wire_9436)
    );

    bfr new_Jinkela_buffer_89 (
        .din(N65),
        .dout(new_Jinkela_wire_97)
    );

    spl4L new_Jinkela_splitter_756 (
        .a(new_Jinkela_wire_9437),
        .d(new_Jinkela_wire_9438),
        .b(new_Jinkela_wire_9439),
        .e(new_Jinkela_wire_9440),
        .c(new_Jinkela_wire_9441)
    );

    bfr new_Jinkela_buffer_23 (
        .din(new_Jinkela_wire_24),
        .dout(new_Jinkela_wire_25)
    );

    spl3L new_Jinkela_splitter_757 (
        .a(new_Jinkela_wire_9441),
        .d(new_Jinkela_wire_9442),
        .b(new_Jinkela_wire_9443),
        .c(new_Jinkela_wire_9444)
    );

    bfr new_Jinkela_buffer_86 (
        .din(new_Jinkela_wire_93),
        .dout(new_Jinkela_wire_94)
    );

    bfr new_Jinkela_buffer_7566 (
        .din(n_0014_),
        .dout(new_Jinkela_wire_9486)
    );

    bfr new_Jinkela_buffer_7562 (
        .din(new_Jinkela_wire_9477),
        .dout(new_Jinkela_wire_9478)
    );

    bfr new_Jinkela_buffer_24 (
        .din(new_Jinkela_wire_25),
        .dout(new_Jinkela_wire_26)
    );

    spl4L new_Jinkela_splitter_760 (
        .a(new_Jinkela_wire_9451),
        .d(new_Jinkela_wire_9452),
        .b(new_Jinkela_wire_9453),
        .e(new_Jinkela_wire_9454),
        .c(new_Jinkela_wire_9455)
    );

    bfr new_Jinkela_buffer_93 (
        .din(N144),
        .dout(new_Jinkela_wire_101)
    );

    spl4L new_Jinkela_splitter_759 (
        .a(new_Jinkela_wire_9446),
        .d(new_Jinkela_wire_9447),
        .b(new_Jinkela_wire_9448),
        .e(new_Jinkela_wire_9449),
        .c(new_Jinkela_wire_9450)
    );

    bfr new_Jinkela_buffer_25 (
        .din(new_Jinkela_wire_26),
        .dout(new_Jinkela_wire_27)
    );

    spl2 new_Jinkela_splitter_763 (
        .a(new_Jinkela_wire_9465),
        .b(new_Jinkela_wire_9466),
        .c(new_Jinkela_wire_9467)
    );

    bfr new_Jinkela_buffer_87 (
        .din(new_Jinkela_wire_94),
        .dout(new_Jinkela_wire_95)
    );

    spl4L new_Jinkela_splitter_761 (
        .a(new_Jinkela_wire_9456),
        .d(new_Jinkela_wire_9457),
        .b(new_Jinkela_wire_9458),
        .e(new_Jinkela_wire_9459),
        .c(new_Jinkela_wire_9460)
    );

    bfr new_Jinkela_buffer_26 (
        .din(new_Jinkela_wire_27),
        .dout(new_Jinkela_wire_28)
    );

    spl4L new_Jinkela_splitter_762 (
        .a(new_Jinkela_wire_9461),
        .d(new_Jinkela_wire_9462),
        .b(new_Jinkela_wire_9463),
        .e(new_Jinkela_wire_9464),
        .c(new_Jinkela_wire_9465)
    );

    bfr new_Jinkela_buffer_90 (
        .din(new_Jinkela_wire_97),
        .dout(new_Jinkela_wire_98)
    );

    bfr new_Jinkela_buffer_27 (
        .din(new_Jinkela_wire_28),
        .dout(new_Jinkela_wire_29)
    );

    bfr new_Jinkela_buffer_7563 (
        .din(new_Jinkela_wire_9478),
        .dout(new_Jinkela_wire_9479)
    );

    spl2 new_Jinkela_splitter_3 (
        .a(N343),
        .b(new_Jinkela_wire_105),
        .c(new_Jinkela_wire_106)
    );

    bfr new_Jinkela_buffer_161 (
        .din(N85),
        .dout(new_Jinkela_wire_173)
    );

    bfr new_Jinkela_buffer_7565 (
        .din(n_0295_),
        .dout(new_Jinkela_wire_9485)
    );

    bfr new_Jinkela_buffer_4972 (
        .din(new_Jinkela_wire_5925),
        .dout(new_Jinkela_wire_5926)
    );

    spl4L new_Jinkela_splitter_73 (
        .a(new_Jinkela_wire_1308),
        .d(new_Jinkela_wire_1309),
        .b(new_Jinkela_wire_1310),
        .e(new_Jinkela_wire_1311),
        .c(new_Jinkela_wire_1312)
    );

    bfr new_Jinkela_buffer_4910 (
        .din(new_Jinkela_wire_5846),
        .dout(new_Jinkela_wire_5847)
    );

    spl4L new_Jinkela_splitter_78 (
        .a(new_Jinkela_wire_1329),
        .d(new_Jinkela_wire_1330),
        .b(new_Jinkela_wire_1331),
        .e(new_Jinkela_wire_1332),
        .c(new_Jinkela_wire_1333)
    );

    bfr new_Jinkela_buffer_4957 (
        .din(new_Jinkela_wire_5906),
        .dout(new_Jinkela_wire_5907)
    );

    spl4L new_Jinkela_splitter_75 (
        .a(new_Jinkela_wire_1318),
        .d(new_Jinkela_wire_1319),
        .b(new_Jinkela_wire_1320),
        .e(new_Jinkela_wire_1321),
        .c(new_Jinkela_wire_1322)
    );

    bfr new_Jinkela_buffer_4911 (
        .din(new_Jinkela_wire_5847),
        .dout(new_Jinkela_wire_5848)
    );

    spl4L new_Jinkela_splitter_76 (
        .a(new_Jinkela_wire_1323),
        .d(new_Jinkela_wire_1324),
        .b(new_Jinkela_wire_1325),
        .e(new_Jinkela_wire_1326),
        .c(new_Jinkela_wire_1327)
    );

    bfr new_Jinkela_buffer_4977 (
        .din(new_Jinkela_wire_5930),
        .dout(new_Jinkela_wire_5931)
    );

    spl4L new_Jinkela_splitter_82 (
        .a(new_Jinkela_wire_1349),
        .d(new_Jinkela_wire_1350),
        .b(new_Jinkela_wire_1355),
        .e(new_Jinkela_wire_1360),
        .c(new_Jinkela_wire_1365)
    );

    bfr new_Jinkela_buffer_4912 (
        .din(new_Jinkela_wire_5848),
        .dout(new_Jinkela_wire_5849)
    );

    spl4L new_Jinkela_splitter_79 (
        .a(new_Jinkela_wire_1334),
        .d(new_Jinkela_wire_1335),
        .b(new_Jinkela_wire_1336),
        .e(new_Jinkela_wire_1337),
        .c(new_Jinkela_wire_1338)
    );

    bfr new_Jinkela_buffer_4958 (
        .din(new_Jinkela_wire_5907),
        .dout(new_Jinkela_wire_5908)
    );

    spl4L new_Jinkela_splitter_83 (
        .a(new_Jinkela_wire_1350),
        .d(new_Jinkela_wire_1351),
        .b(new_Jinkela_wire_1352),
        .e(new_Jinkela_wire_1353),
        .c(new_Jinkela_wire_1354)
    );

    bfr new_Jinkela_buffer_4913 (
        .din(new_Jinkela_wire_5849),
        .dout(new_Jinkela_wire_5850)
    );

    spl4L new_Jinkela_splitter_80 (
        .a(new_Jinkela_wire_1339),
        .d(new_Jinkela_wire_1340),
        .b(new_Jinkela_wire_1341),
        .e(new_Jinkela_wire_1342),
        .c(new_Jinkela_wire_1343)
    );

    spl4L new_Jinkela_splitter_81 (
        .a(new_Jinkela_wire_1344),
        .d(new_Jinkela_wire_1345),
        .b(new_Jinkela_wire_1346),
        .e(new_Jinkela_wire_1347),
        .c(new_Jinkela_wire_1348)
    );

    bfr new_Jinkela_buffer_4914 (
        .din(new_Jinkela_wire_5850),
        .dout(new_Jinkela_wire_5851)
    );

    spl4L new_Jinkela_splitter_87 (
        .a(new_Jinkela_wire_1370),
        .d(new_Jinkela_wire_1371),
        .b(new_Jinkela_wire_1376),
        .e(new_Jinkela_wire_1381),
        .c(new_Jinkela_wire_1386)
    );

    bfr new_Jinkela_buffer_5017 (
        .din(n_0547_),
        .dout(new_Jinkela_wire_5977)
    );

    bfr new_Jinkela_buffer_4959 (
        .din(new_Jinkela_wire_5908),
        .dout(new_Jinkela_wire_5909)
    );

    spl4L new_Jinkela_splitter_84 (
        .a(new_Jinkela_wire_1355),
        .d(new_Jinkela_wire_1356),
        .b(new_Jinkela_wire_1357),
        .e(new_Jinkela_wire_1358),
        .c(new_Jinkela_wire_1359)
    );

    bfr new_Jinkela_buffer_4915 (
        .din(new_Jinkela_wire_5851),
        .dout(new_Jinkela_wire_5852)
    );

    spl4L new_Jinkela_splitter_88 (
        .a(new_Jinkela_wire_1371),
        .d(new_Jinkela_wire_1372),
        .b(new_Jinkela_wire_1373),
        .e(new_Jinkela_wire_1374),
        .c(new_Jinkela_wire_1375)
    );

    bfr new_Jinkela_buffer_4978 (
        .din(new_Jinkela_wire_5931),
        .dout(new_Jinkela_wire_5932)
    );

    spl4L new_Jinkela_splitter_85 (
        .a(new_Jinkela_wire_1360),
        .d(new_Jinkela_wire_1361),
        .b(new_Jinkela_wire_1362),
        .e(new_Jinkela_wire_1363),
        .c(new_Jinkela_wire_1364)
    );

    bfr new_Jinkela_buffer_4916 (
        .din(new_Jinkela_wire_5852),
        .dout(new_Jinkela_wire_5853)
    );

    spl4L new_Jinkela_splitter_86 (
        .a(new_Jinkela_wire_1365),
        .d(new_Jinkela_wire_1366),
        .b(new_Jinkela_wire_1367),
        .e(new_Jinkela_wire_1368),
        .c(new_Jinkela_wire_1369)
    );

    bfr new_Jinkela_buffer_4960 (
        .din(new_Jinkela_wire_5909),
        .dout(new_Jinkela_wire_5910)
    );

    bfr new_Jinkela_buffer_4917 (
        .din(new_Jinkela_wire_5853),
        .dout(new_Jinkela_wire_5854)
    );

    bfr new_Jinkela_buffer_1105 (
        .din(new_Jinkela_wire_1416),
        .dout(new_Jinkela_wire_1417)
    );

    spl4L new_Jinkela_splitter_89 (
        .a(new_Jinkela_wire_1376),
        .d(new_Jinkela_wire_1377),
        .b(new_Jinkela_wire_1378),
        .e(new_Jinkela_wire_1379),
        .c(new_Jinkela_wire_1380)
    );

    spl2 new_Jinkela_splitter_92 (
        .a(new_Jinkela_wire_1390),
        .b(new_Jinkela_wire_1391),
        .c(new_Jinkela_wire_1392)
    );

    bfr new_Jinkela_buffer_4918 (
        .din(new_Jinkela_wire_5854),
        .dout(new_Jinkela_wire_5855)
    );

    spl4L new_Jinkela_splitter_90 (
        .a(new_Jinkela_wire_1381),
        .d(new_Jinkela_wire_1382),
        .b(new_Jinkela_wire_1383),
        .e(new_Jinkela_wire_1384),
        .c(new_Jinkela_wire_1385)
    );

    bfr new_Jinkela_buffer_4979 (
        .din(new_Jinkela_wire_5936),
        .dout(new_Jinkela_wire_5937)
    );

    bfr new_Jinkela_buffer_4961 (
        .din(new_Jinkela_wire_5910),
        .dout(new_Jinkela_wire_5911)
    );

    spl4L new_Jinkela_splitter_91 (
        .a(new_Jinkela_wire_1386),
        .d(new_Jinkela_wire_1387),
        .b(new_Jinkela_wire_1388),
        .e(new_Jinkela_wire_1389),
        .c(new_Jinkela_wire_1390)
    );

    bfr new_Jinkela_buffer_4919 (
        .din(new_Jinkela_wire_5855),
        .dout(new_Jinkela_wire_5856)
    );

    bfr new_Jinkela_buffer_5011 (
        .din(new_Jinkela_wire_5970),
        .dout(new_Jinkela_wire_5971)
    );

    bfr new_Jinkela_buffer_1290 (
        .din(new_Jinkela_wire_1610),
        .dout(new_Jinkela_wire_1611)
    );

    bfr new_Jinkela_buffer_4920 (
        .din(new_Jinkela_wire_5856),
        .dout(new_Jinkela_wire_5857)
    );

    bfr new_Jinkela_buffer_1106 (
        .din(new_Jinkela_wire_1417),
        .dout(new_Jinkela_wire_1418)
    );

    spl2 new_Jinkela_splitter_93 (
        .a(new_Jinkela_wire_1392),
        .b(new_Jinkela_wire_1393),
        .c(new_Jinkela_wire_1394)
    );

    bfr new_Jinkela_buffer_4962 (
        .din(new_Jinkela_wire_5911),
        .dout(new_Jinkela_wire_5912)
    );

    bfr new_Jinkela_buffer_4921 (
        .din(new_Jinkela_wire_5857),
        .dout(new_Jinkela_wire_5858)
    );

    bfr new_Jinkela_buffer_1165 (
        .din(new_Jinkela_wire_1478),
        .dout(new_Jinkela_wire_1479)
    );

    bfr new_Jinkela_buffer_4980 (
        .din(new_Jinkela_wire_5937),
        .dout(new_Jinkela_wire_5938)
    );

    spl2 new_Jinkela_splitter_99 (
        .a(new_Jinkela_wire_1544),
        .b(new_Jinkela_wire_1545),
        .c(new_Jinkela_wire_1546)
    );

    bfr new_Jinkela_buffer_4922 (
        .din(new_Jinkela_wire_5858),
        .dout(new_Jinkela_wire_5859)
    );

    bfr new_Jinkela_buffer_1107 (
        .din(new_Jinkela_wire_1418),
        .dout(new_Jinkela_wire_1419)
    );

    bfr new_Jinkela_buffer_4963 (
        .din(new_Jinkela_wire_5912),
        .dout(new_Jinkela_wire_5913)
    );

    bfr new_Jinkela_buffer_1108 (
        .din(new_Jinkela_wire_1419),
        .dout(new_Jinkela_wire_1420)
    );

    bfr new_Jinkela_buffer_4923 (
        .din(new_Jinkela_wire_5859),
        .dout(new_Jinkela_wire_5860)
    );

    spl3L new_Jinkela_splitter_97 (
        .a(new_Jinkela_wire_1479),
        .d(new_Jinkela_wire_1480),
        .b(new_Jinkela_wire_1481),
        .c(new_Jinkela_wire_1482)
    );

    bfr new_Jinkela_buffer_5018 (
        .din(n_1164_),
        .dout(new_Jinkela_wire_5978)
    );

    bfr new_Jinkela_buffer_1109 (
        .din(new_Jinkela_wire_1420),
        .dout(new_Jinkela_wire_1421)
    );

    bfr new_Jinkela_buffer_4924 (
        .din(new_Jinkela_wire_5860),
        .dout(new_Jinkela_wire_5861)
    );

    bfr new_Jinkela_buffer_1226 (
        .din(new_Jinkela_wire_1546),
        .dout(new_Jinkela_wire_1547)
    );

    bfr new_Jinkela_buffer_4964 (
        .din(new_Jinkela_wire_5913),
        .dout(new_Jinkela_wire_5914)
    );

    bfr new_Jinkela_buffer_1110 (
        .din(new_Jinkela_wire_1421),
        .dout(new_Jinkela_wire_1422)
    );

    bfr new_Jinkela_buffer_4925 (
        .din(new_Jinkela_wire_5861),
        .dout(new_Jinkela_wire_5862)
    );

    bfr new_Jinkela_buffer_1166 (
        .din(new_Jinkela_wire_1482),
        .dout(new_Jinkela_wire_1483)
    );

    bfr new_Jinkela_buffer_4981 (
        .din(new_Jinkela_wire_5938),
        .dout(new_Jinkela_wire_5939)
    );

    bfr new_Jinkela_buffer_1111 (
        .din(new_Jinkela_wire_1422),
        .dout(new_Jinkela_wire_1423)
    );

    bfr new_Jinkela_buffer_4926 (
        .din(new_Jinkela_wire_5862),
        .dout(new_Jinkela_wire_5863)
    );

    bfr new_Jinkela_buffer_1357 (
        .din(N81),
        .dout(new_Jinkela_wire_1683)
    );

    bfr new_Jinkela_buffer_4965 (
        .din(new_Jinkela_wire_5914),
        .dout(new_Jinkela_wire_5915)
    );

    bfr new_Jinkela_buffer_1112 (
        .din(new_Jinkela_wire_1423),
        .dout(new_Jinkela_wire_1424)
    );

    bfr new_Jinkela_buffer_4927 (
        .din(new_Jinkela_wire_5863),
        .dout(new_Jinkela_wire_5864)
    );

    bfr new_Jinkela_buffer_1167 (
        .din(new_Jinkela_wire_1483),
        .dout(new_Jinkela_wire_1484)
    );

    bfr new_Jinkela_buffer_5012 (
        .din(new_Jinkela_wire_5971),
        .dout(new_Jinkela_wire_5972)
    );

    bfr new_Jinkela_buffer_1113 (
        .din(new_Jinkela_wire_1424),
        .dout(new_Jinkela_wire_1425)
    );

    bfr new_Jinkela_buffer_4928 (
        .din(new_Jinkela_wire_5864),
        .dout(new_Jinkela_wire_5865)
    );

    bfr new_Jinkela_buffer_1291 (
        .din(new_Jinkela_wire_1611),
        .dout(new_Jinkela_wire_1612)
    );

    bfr new_Jinkela_buffer_4966 (
        .din(new_Jinkela_wire_5915),
        .dout(new_Jinkela_wire_5916)
    );

    bfr new_Jinkela_buffer_1114 (
        .din(new_Jinkela_wire_1425),
        .dout(new_Jinkela_wire_1426)
    );

    bfr new_Jinkela_buffer_4929 (
        .din(new_Jinkela_wire_5865),
        .dout(new_Jinkela_wire_5866)
    );

    bfr new_Jinkela_buffer_1168 (
        .din(new_Jinkela_wire_1484),
        .dout(new_Jinkela_wire_1485)
    );

    bfr new_Jinkela_buffer_4982 (
        .din(new_Jinkela_wire_5939),
        .dout(new_Jinkela_wire_5940)
    );

    bfr new_Jinkela_buffer_1115 (
        .din(new_Jinkela_wire_1426),
        .dout(new_Jinkela_wire_1427)
    );

    bfr new_Jinkela_buffer_4930 (
        .din(new_Jinkela_wire_5866),
        .dout(new_Jinkela_wire_5867)
    );

    bfr new_Jinkela_buffer_1227 (
        .din(new_Jinkela_wire_1547),
        .dout(new_Jinkela_wire_1548)
    );

    and_bi n_1821_ (
        .a(new_Jinkela_wire_100),
        .b(new_Jinkela_wire_1247),
        .c(n_1088_)
    );

    or_bi n_2535_ (
        .a(new_Jinkela_wire_10416),
        .b(new_Jinkela_wire_9419),
        .c(n_0395_)
    );

    bfr new_Jinkela_buffer_5762 (
        .din(new_Jinkela_wire_6955),
        .dout(new_Jinkela_wire_6956)
    );

    and_bi n_1822_ (
        .a(new_Jinkela_wire_1343),
        .b(new_Jinkela_wire_2595),
        .c(n_1089_)
    );

    and_bi n_2536_ (
        .a(new_Jinkela_wire_10415),
        .b(new_Jinkela_wire_9420),
        .c(n_0396_)
    );

    bfr new_Jinkela_buffer_5821 (
        .din(new_net_2489),
        .dout(new_Jinkela_wire_7023)
    );

    spl3L new_Jinkela_splitter_468 (
        .a(n_0113_),
        .d(new_Jinkela_wire_7024),
        .b(new_Jinkela_wire_7025),
        .c(new_Jinkela_wire_7026)
    );

    and_ii n_1823_ (
        .a(n_1089_),
        .b(n_1088_),
        .c(n_1090_)
    );

    and_bi n_2537_ (
        .a(n_0395_),
        .b(n_0396_),
        .c(new_net_2576)
    );

    bfr new_Jinkela_buffer_5763 (
        .din(new_Jinkela_wire_6956),
        .dout(new_Jinkela_wire_6957)
    );

    and_bi n_1824_ (
        .a(new_Jinkela_wire_4655),
        .b(new_Jinkela_wire_7117),
        .c(n_1091_)
    );

    and_ii n_2538_ (
        .a(new_Jinkela_wire_9252),
        .b(new_Jinkela_wire_8663),
        .c(n_0397_)
    );

    spl2 new_Jinkela_splitter_469 (
        .a(n_0349_),
        .b(new_Jinkela_wire_7067),
        .c(new_Jinkela_wire_7068)
    );

    bfr new_Jinkela_buffer_5820 (
        .din(new_Jinkela_wire_7021),
        .dout(new_Jinkela_wire_7022)
    );

    and_bi n_1825_ (
        .a(new_Jinkela_wire_7116),
        .b(new_Jinkela_wire_4654),
        .c(n_1092_)
    );

    or_bb n_2539_ (
        .a(new_Jinkela_wire_7385),
        .b(new_Jinkela_wire_7416),
        .c(n_0398_)
    );

    bfr new_Jinkela_buffer_5764 (
        .din(new_Jinkela_wire_6957),
        .dout(new_Jinkela_wire_6958)
    );

    and_ii n_1826_ (
        .a(n_1092_),
        .b(n_1091_),
        .c(n_1093_)
    );

    and_bi n_2540_ (
        .a(new_Jinkela_wire_8481),
        .b(new_Jinkela_wire_8409),
        .c(n_0399_)
    );

    spl3L new_Jinkela_splitter_470 (
        .a(n_0782_),
        .d(new_Jinkela_wire_7069),
        .b(new_Jinkela_wire_7070),
        .c(new_Jinkela_wire_7071)
    );

    and_bi n_1827_ (
        .a(new_Jinkela_wire_83),
        .b(new_Jinkela_wire_1236),
        .c(n_1094_)
    );

    and_bi n_2541_ (
        .a(new_Jinkela_wire_8408),
        .b(new_Jinkela_wire_8480),
        .c(n_0400_)
    );

    bfr new_Jinkela_buffer_5765 (
        .din(new_Jinkela_wire_6958),
        .dout(new_Jinkela_wire_6959)
    );

    and_bi n_1828_ (
        .a(new_Jinkela_wire_1171),
        .b(new_Jinkela_wire_3367),
        .c(n_1095_)
    );

    and_ii n_2542_ (
        .a(n_0400_),
        .b(n_0399_),
        .c(n_0401_)
    );

    bfr new_Jinkela_buffer_5862 (
        .din(n_0630_),
        .dout(new_Jinkela_wire_7083)
    );

    bfr new_Jinkela_buffer_5822 (
        .din(new_Jinkela_wire_7026),
        .dout(new_Jinkela_wire_7027)
    );

    and_ii n_1829_ (
        .a(n_1095_),
        .b(n_1094_),
        .c(n_1096_)
    );

    and_ii n_2543_ (
        .a(new_Jinkela_wire_4916),
        .b(new_Jinkela_wire_9410),
        .c(n_0402_)
    );

    bfr new_Jinkela_buffer_5766 (
        .din(new_Jinkela_wire_6959),
        .dout(new_Jinkela_wire_6960)
    );

    or_ii n_1830_ (
        .a(new_Jinkela_wire_8321),
        .b(new_Jinkela_wire_5236),
        .c(n_1097_)
    );

    and_bi n_2544_ (
        .a(new_Jinkela_wire_7956),
        .b(new_Jinkela_wire_4018),
        .c(n_0403_)
    );

    or_bb n_1831_ (
        .a(new_Jinkela_wire_8320),
        .b(new_Jinkela_wire_5235),
        .c(n_1098_)
    );

    and_bi n_2545_ (
        .a(new_Jinkela_wire_9342),
        .b(new_Jinkela_wire_7334),
        .c(n_0404_)
    );

    bfr new_Jinkela_buffer_5767 (
        .din(new_Jinkela_wire_6960),
        .dout(new_Jinkela_wire_6961)
    );

    or_ii n_1832_ (
        .a(n_1098_),
        .b(n_1097_),
        .c(n_1099_)
    );

    and_ii n_2546_ (
        .a(new_Jinkela_wire_4537),
        .b(new_Jinkela_wire_9341),
        .c(n_0405_)
    );

    and_bi n_1833_ (
        .a(new_Jinkela_wire_3562),
        .b(new_Jinkela_wire_1287),
        .c(n_1100_)
    );

    and_ii n_2547_ (
        .a(n_0405_),
        .b(n_0404_),
        .c(n_0406_)
    );

    bfr new_Jinkela_buffer_5768 (
        .din(new_Jinkela_wire_6961),
        .dout(new_Jinkela_wire_6962)
    );

    and_bi n_1834_ (
        .a(new_Jinkela_wire_1274),
        .b(new_Jinkela_wire_952),
        .c(n_1101_)
    );

    and_bi n_2548_ (
        .a(new_Jinkela_wire_9340),
        .b(new_Jinkela_wire_7922),
        .c(n_0407_)
    );

    bfr new_Jinkela_buffer_5823 (
        .din(new_Jinkela_wire_7027),
        .dout(new_Jinkela_wire_7028)
    );

    and_ii n_1835_ (
        .a(n_1101_),
        .b(n_1100_),
        .c(n_1102_)
    );

    and_bi n_2549_ (
        .a(new_Jinkela_wire_7921),
        .b(new_Jinkela_wire_9339),
        .c(n_0408_)
    );

    bfr new_Jinkela_buffer_5769 (
        .din(new_Jinkela_wire_6962),
        .dout(new_Jinkela_wire_6963)
    );

    and_bi n_1836_ (
        .a(new_Jinkela_wire_608),
        .b(new_Jinkela_wire_1342),
        .c(n_1103_)
    );

    and_ii n_2550_ (
        .a(n_0408_),
        .b(n_0407_),
        .c(n_0409_)
    );

    spl2 new_Jinkela_splitter_471 (
        .a(n_1163_),
        .b(new_Jinkela_wire_7072),
        .c(new_Jinkela_wire_7073)
    );

    spl2 new_Jinkela_splitter_472 (
        .a(n_0418_),
        .b(new_Jinkela_wire_7074),
        .c(new_Jinkela_wire_7075)
    );

    and_bi n_1837_ (
        .a(new_Jinkela_wire_1333),
        .b(new_Jinkela_wire_1617),
        .c(n_1104_)
    );

    and_bb n_2551_ (
        .a(new_Jinkela_wire_8449),
        .b(new_Jinkela_wire_7302),
        .c(n_0410_)
    );

    bfr new_Jinkela_buffer_5770 (
        .din(new_Jinkela_wire_6963),
        .dout(new_Jinkela_wire_6964)
    );

    and_ii n_1838_ (
        .a(n_1104_),
        .b(n_1103_),
        .c(n_1105_)
    );

    and_ii n_2552_ (
        .a(new_Jinkela_wire_8448),
        .b(new_Jinkela_wire_7301),
        .c(n_0411_)
    );

    bfr new_Jinkela_buffer_5824 (
        .din(new_Jinkela_wire_7028),
        .dout(new_Jinkela_wire_7029)
    );

    and_bi n_1839_ (
        .a(new_Jinkela_wire_7247),
        .b(new_Jinkela_wire_8397),
        .c(n_1106_)
    );

    or_bb n_2553_ (
        .a(n_0411_),
        .b(n_0410_),
        .c(n_0412_)
    );

    bfr new_Jinkela_buffer_5771 (
        .din(new_Jinkela_wire_6964),
        .dout(new_Jinkela_wire_6965)
    );

    and_bi n_1840_ (
        .a(new_Jinkela_wire_8396),
        .b(new_Jinkela_wire_7246),
        .c(n_1107_)
    );

    or_bb n_2554_ (
        .a(new_Jinkela_wire_10447),
        .b(new_Jinkela_wire_7269),
        .c(n_0413_)
    );

    and_ii n_1841_ (
        .a(n_1107_),
        .b(n_1106_),
        .c(n_1108_)
    );

    and_bb n_2555_ (
        .a(new_Jinkela_wire_10446),
        .b(new_Jinkela_wire_7268),
        .c(n_0414_)
    );

    bfr new_Jinkela_buffer_5772 (
        .din(new_Jinkela_wire_6965),
        .dout(new_Jinkela_wire_6966)
    );

    and_bi n_1842_ (
        .a(new_Jinkela_wire_2808),
        .b(new_Jinkela_wire_1234),
        .c(n_1109_)
    );

    and_bi n_2556_ (
        .a(n_0413_),
        .b(n_0414_),
        .c(n_0415_)
    );

    bfr new_Jinkela_buffer_5825 (
        .din(new_Jinkela_wire_7029),
        .dout(new_Jinkela_wire_7030)
    );

    and_bi n_1843_ (
        .a(new_Jinkela_wire_1288),
        .b(new_Jinkela_wire_1406),
        .c(n_1110_)
    );

    or_bb n_2557_ (
        .a(new_Jinkela_wire_7294),
        .b(new_Jinkela_wire_8375),
        .c(n_0416_)
    );

    bfr new_Jinkela_buffer_5773 (
        .din(new_Jinkela_wire_6966),
        .dout(new_Jinkela_wire_6967)
    );

    and_ii n_1844_ (
        .a(n_1110_),
        .b(n_1109_),
        .c(n_1111_)
    );

    and_ii n_2558_ (
        .a(new_Jinkela_wire_7336),
        .b(new_Jinkela_wire_7462),
        .c(n_0417_)
    );

    spl3L new_Jinkela_splitter_473 (
        .a(n_1045_),
        .d(new_Jinkela_wire_7076),
        .b(new_Jinkela_wire_7077),
        .c(new_Jinkela_wire_7078)
    );

    or_bb n_1845_ (
        .a(new_Jinkela_wire_10228),
        .b(new_Jinkela_wire_4504),
        .c(n_1112_)
    );

    and_ii n_2559_ (
        .a(new_Jinkela_wire_6791),
        .b(new_Jinkela_wire_7234),
        .c(n_0418_)
    );

    bfr new_Jinkela_buffer_5774 (
        .din(new_Jinkela_wire_6967),
        .dout(new_Jinkela_wire_6968)
    );

    or_ii n_1846_ (
        .a(new_Jinkela_wire_10227),
        .b(new_Jinkela_wire_4503),
        .c(n_1113_)
    );

    and_bi n_2560_ (
        .a(new_Jinkela_wire_7075),
        .b(new_Jinkela_wire_4877),
        .c(n_0419_)
    );

    bfr new_Jinkela_buffer_5826 (
        .din(new_Jinkela_wire_7030),
        .dout(new_Jinkela_wire_7031)
    );

    or_ii n_1847_ (
        .a(n_1113_),
        .b(n_1112_),
        .c(n_1114_)
    );

    and_bi n_2561_ (
        .a(new_Jinkela_wire_4876),
        .b(new_Jinkela_wire_7074),
        .c(n_0420_)
    );

    bfr new_Jinkela_buffer_5775 (
        .din(new_Jinkela_wire_6968),
        .dout(new_Jinkela_wire_6969)
    );

    and_ii n_1848_ (
        .a(new_Jinkela_wire_9090),
        .b(new_Jinkela_wire_4628),
        .c(n_1115_)
    );

    and_ii n_2562_ (
        .a(n_0420_),
        .b(n_0419_),
        .c(n_0421_)
    );

    spl2 new_Jinkela_splitter_474 (
        .a(new_Jinkela_wire_7078),
        .b(new_Jinkela_wire_7079),
        .c(new_Jinkela_wire_7080)
    );

    spl2 new_Jinkela_splitter_475 (
        .a(n_0811_),
        .b(new_Jinkela_wire_7081),
        .c(new_Jinkela_wire_7082)
    );

    and_bb n_1849_ (
        .a(new_Jinkela_wire_9089),
        .b(new_Jinkela_wire_4627),
        .c(n_1116_)
    );

    and_bi n_2563_ (
        .a(new_Jinkela_wire_7952),
        .b(new_Jinkela_wire_8373),
        .c(n_0422_)
    );

    bfr new_Jinkela_buffer_5776 (
        .din(new_Jinkela_wire_6969),
        .dout(new_Jinkela_wire_6970)
    );

    and_ii n_1850_ (
        .a(n_1116_),
        .b(n_1115_),
        .c(n_1117_)
    );

    and_bi n_2564_ (
        .a(new_Jinkela_wire_8372),
        .b(new_Jinkela_wire_7954),
        .c(n_0423_)
    );

    bfr new_Jinkela_buffer_5827 (
        .din(new_Jinkela_wire_7031),
        .dout(new_Jinkela_wire_7032)
    );

    and_bi n_1851_ (
        .a(new_Jinkela_wire_6334),
        .b(new_Jinkela_wire_7989),
        .c(n_1118_)
    );

    and_ii n_2565_ (
        .a(n_0423_),
        .b(n_0422_),
        .c(n_0424_)
    );

    bfr new_Jinkela_buffer_5777 (
        .din(new_Jinkela_wire_6970),
        .dout(new_Jinkela_wire_6971)
    );

    and_bi n_1852_ (
        .a(new_Jinkela_wire_7988),
        .b(new_Jinkela_wire_6333),
        .c(n_1119_)
    );

    and_bb n_2566_ (
        .a(new_Jinkela_wire_8090),
        .b(new_Jinkela_wire_4914),
        .c(n_0425_)
    );

    spl2 new_Jinkela_splitter_476 (
        .a(n_0253_),
        .b(new_Jinkela_wire_7086),
        .c(new_Jinkela_wire_7087)
    );

    or_bb n_1853_ (
        .a(n_1119_),
        .b(n_1118_),
        .c(n_1120_)
    );

    and_ii n_2567_ (
        .a(new_Jinkela_wire_8089),
        .b(new_Jinkela_wire_4915),
        .c(n_0426_)
    );

    bfr new_Jinkela_buffer_5778 (
        .din(new_Jinkela_wire_6971),
        .dout(new_Jinkela_wire_6972)
    );

    or_bb n_1854_ (
        .a(n_1120_),
        .b(n_1063_),
        .c(n_1121_)
    );

    or_bb n_2568_ (
        .a(n_0426_),
        .b(n_0425_),
        .c(n_0427_)
    );

    bfr new_Jinkela_buffer_5828 (
        .din(new_Jinkela_wire_7032),
        .dout(new_Jinkela_wire_7033)
    );

    or_bb n_1855_ (
        .a(n_1121_),
        .b(n_1006_),
        .c(new_net_6)
    );

    and_bi n_2569_ (
        .a(new_Jinkela_wire_8376),
        .b(new_Jinkela_wire_8994),
        .c(n_0428_)
    );

    bfr new_Jinkela_buffer_5779 (
        .din(new_Jinkela_wire_6972),
        .dout(new_Jinkela_wire_6973)
    );

    and_ii n_1856_ (
        .a(new_Jinkela_wire_6261),
        .b(new_Jinkela_wire_2156),
        .c(n_1122_)
    );

    and_bi n_2570_ (
        .a(n_0416_),
        .b(n_0428_),
        .c(n_0429_)
    );

    bfr new_Jinkela_buffer_5863 (
        .din(new_Jinkela_wire_7083),
        .dout(new_Jinkela_wire_7084)
    );

    and_bi n_1857_ (
        .a(new_Jinkela_wire_1193),
        .b(new_Jinkela_wire_1814),
        .c(n_1123_)
    );

    and_ii n_2571_ (
        .a(new_Jinkela_wire_3719),
        .b(new_Jinkela_wire_9111),
        .c(n_0430_)
    );

    bfr new_Jinkela_buffer_5780 (
        .din(new_Jinkela_wire_6973),
        .dout(new_Jinkela_wire_6974)
    );

    and_ii n_1858_ (
        .a(new_Jinkela_wire_6891),
        .b(new_Jinkela_wire_9455),
        .c(n_1124_)
    );

    or_bb n_2572_ (
        .a(new_Jinkela_wire_4502),
        .b(new_Jinkela_wire_7453),
        .c(n_0431_)
    );

    bfr new_Jinkela_buffer_5829 (
        .din(new_Jinkela_wire_7033),
        .dout(new_Jinkela_wire_7034)
    );

    and_bi n_1859_ (
        .a(new_Jinkela_wire_1176),
        .b(new_Jinkela_wire_271),
        .c(n_1125_)
    );

    or_bi n_2573_ (
        .a(new_Jinkela_wire_8370),
        .b(new_Jinkela_wire_6671),
        .c(n_0432_)
    );

    bfr new_Jinkela_buffer_5781 (
        .din(new_Jinkela_wire_6974),
        .dout(new_Jinkela_wire_6975)
    );

    and_bb n_1860_ (
        .a(new_Jinkela_wire_5400),
        .b(new_Jinkela_wire_7309),
        .c(n_1126_)
    );

    and_bi n_2574_ (
        .a(new_Jinkela_wire_8369),
        .b(new_Jinkela_wire_6670),
        .c(n_0433_)
    );

    spl3L new_Jinkela_splitter_477 (
        .a(n_0785_),
        .d(new_Jinkela_wire_7089),
        .b(new_Jinkela_wire_7090),
        .c(new_Jinkela_wire_7091)
    );

    or_bb n_1861_ (
        .a(new_Jinkela_wire_5397),
        .b(new_Jinkela_wire_9450),
        .c(n_1127_)
    );

    and_bi n_2575_ (
        .a(n_0432_),
        .b(n_0433_),
        .c(n_0434_)
    );

    bfr new_Jinkela_buffer_5782 (
        .din(new_Jinkela_wire_6975),
        .dout(new_Jinkela_wire_6976)
    );

    and_bi n_1862_ (
        .a(new_Jinkela_wire_6894),
        .b(new_Jinkela_wire_9603),
        .c(n_1128_)
    );

    and_bi n_2576_ (
        .a(new_Jinkela_wire_5106),
        .b(new_Jinkela_wire_10428),
        .c(n_0435_)
    );

    bfr new_Jinkela_buffer_5830 (
        .din(new_Jinkela_wire_7034),
        .dout(new_Jinkela_wire_7035)
    );

    spl3L new_Jinkela_splitter_598 (
        .a(n_1364_),
        .d(new_Jinkela_wire_8181),
        .b(new_Jinkela_wire_8182),
        .c(new_Jinkela_wire_8183)
    );

    bfr new_Jinkela_buffer_6625 (
        .din(new_Jinkela_wire_8110),
        .dout(new_Jinkela_wire_8111)
    );

    bfr new_Jinkela_buffer_6582 (
        .din(new_Jinkela_wire_8048),
        .dout(new_Jinkela_wire_8049)
    );

    bfr new_Jinkela_buffer_6583 (
        .din(new_Jinkela_wire_8049),
        .dout(new_Jinkela_wire_8050)
    );

    bfr new_Jinkela_buffer_6626 (
        .din(new_Jinkela_wire_8111),
        .dout(new_Jinkela_wire_8112)
    );

    bfr new_Jinkela_buffer_6584 (
        .din(new_Jinkela_wire_8050),
        .dout(new_Jinkela_wire_8051)
    );

    bfr new_Jinkela_buffer_6675 (
        .din(n_1152_),
        .dout(new_Jinkela_wire_8179)
    );

    bfr new_Jinkela_buffer_6585 (
        .din(new_Jinkela_wire_8051),
        .dout(new_Jinkela_wire_8052)
    );

    bfr new_Jinkela_buffer_6627 (
        .din(new_Jinkela_wire_8112),
        .dout(new_Jinkela_wire_8113)
    );

    bfr new_Jinkela_buffer_6586 (
        .din(new_Jinkela_wire_8052),
        .dout(new_Jinkela_wire_8053)
    );

    bfr new_Jinkela_buffer_6676 (
        .din(n_1272_),
        .dout(new_Jinkela_wire_8180)
    );

    bfr new_Jinkela_buffer_6587 (
        .din(new_Jinkela_wire_8053),
        .dout(new_Jinkela_wire_8054)
    );

    spl4L new_Jinkela_splitter_599 (
        .a(n_1180_),
        .d(new_Jinkela_wire_8184),
        .b(new_Jinkela_wire_8185),
        .e(new_Jinkela_wire_8186),
        .c(new_Jinkela_wire_8187)
    );

    bfr new_Jinkela_buffer_6628 (
        .din(new_Jinkela_wire_8113),
        .dout(new_Jinkela_wire_8114)
    );

    bfr new_Jinkela_buffer_6588 (
        .din(new_Jinkela_wire_8054),
        .dout(new_Jinkela_wire_8055)
    );

    spl2 new_Jinkela_splitter_600 (
        .a(n_0541_),
        .b(new_Jinkela_wire_8188),
        .c(new_Jinkela_wire_8189)
    );

    bfr new_Jinkela_buffer_6589 (
        .din(new_Jinkela_wire_8055),
        .dout(new_Jinkela_wire_8056)
    );

    bfr new_Jinkela_buffer_6629 (
        .din(new_Jinkela_wire_8114),
        .dout(new_Jinkela_wire_8115)
    );

    bfr new_Jinkela_buffer_6590 (
        .din(new_Jinkela_wire_8056),
        .dout(new_Jinkela_wire_8057)
    );

    spl2 new_Jinkela_splitter_601 (
        .a(n_0839_),
        .b(new_Jinkela_wire_8190),
        .c(new_Jinkela_wire_8191)
    );

    bfr new_Jinkela_buffer_6591 (
        .din(new_Jinkela_wire_8057),
        .dout(new_Jinkela_wire_8058)
    );

    bfr new_Jinkela_buffer_6630 (
        .din(new_Jinkela_wire_8115),
        .dout(new_Jinkela_wire_8116)
    );

    bfr new_Jinkela_buffer_6592 (
        .din(new_Jinkela_wire_8058),
        .dout(new_Jinkela_wire_8059)
    );

    bfr new_Jinkela_buffer_6677 (
        .din(n_0987_),
        .dout(new_Jinkela_wire_8192)
    );

    bfr new_Jinkela_buffer_6593 (
        .din(new_Jinkela_wire_8059),
        .dout(new_Jinkela_wire_8060)
    );

    bfr new_Jinkela_buffer_6631 (
        .din(new_Jinkela_wire_8116),
        .dout(new_Jinkela_wire_8117)
    );

    bfr new_Jinkela_buffer_6594 (
        .din(new_Jinkela_wire_8060),
        .dout(new_Jinkela_wire_8061)
    );

    bfr new_Jinkela_buffer_6595 (
        .din(new_Jinkela_wire_8061),
        .dout(new_Jinkela_wire_8062)
    );

    bfr new_Jinkela_buffer_6632 (
        .din(new_Jinkela_wire_8117),
        .dout(new_Jinkela_wire_8118)
    );

    bfr new_Jinkela_buffer_6596 (
        .din(new_Jinkela_wire_8062),
        .dout(new_Jinkela_wire_8063)
    );

    bfr new_Jinkela_buffer_6597 (
        .din(new_Jinkela_wire_8063),
        .dout(new_Jinkela_wire_8064)
    );

    bfr new_Jinkela_buffer_6633 (
        .din(new_Jinkela_wire_8118),
        .dout(new_Jinkela_wire_8119)
    );

    bfr new_Jinkela_buffer_6598 (
        .din(new_Jinkela_wire_8064),
        .dout(new_Jinkela_wire_8065)
    );

    spl2 new_Jinkela_splitter_604 (
        .a(new_net_1),
        .b(new_Jinkela_wire_8199),
        .c(new_Jinkela_wire_8200)
    );

    bfr new_Jinkela_buffer_6599 (
        .din(new_Jinkela_wire_8065),
        .dout(new_Jinkela_wire_8066)
    );

    spl4L new_Jinkela_splitter_605 (
        .a(n_0103_),
        .d(new_Jinkela_wire_8264),
        .b(new_Jinkela_wire_8265),
        .e(new_Jinkela_wire_8266),
        .c(new_Jinkela_wire_8267)
    );

    bfr new_Jinkela_buffer_6634 (
        .din(new_Jinkela_wire_8119),
        .dout(new_Jinkela_wire_8120)
    );

    bfr new_Jinkela_buffer_6600 (
        .din(new_Jinkela_wire_8066),
        .dout(new_Jinkela_wire_8067)
    );

    bfr new_Jinkela_buffer_6679 (
        .din(new_Jinkela_wire_8200),
        .dout(new_Jinkela_wire_8201)
    );

    bfr new_Jinkela_buffer_6601 (
        .din(new_Jinkela_wire_8067),
        .dout(new_Jinkela_wire_8068)
    );

    spl3L new_Jinkela_splitter_602 (
        .a(new_Jinkela_wire_8192),
        .d(new_Jinkela_wire_8193),
        .b(new_Jinkela_wire_8194),
        .c(new_Jinkela_wire_8195)
    );

    bfr new_Jinkela_buffer_6635 (
        .din(new_Jinkela_wire_8120),
        .dout(new_Jinkela_wire_8121)
    );

    bfr new_Jinkela_buffer_6602 (
        .din(new_Jinkela_wire_8068),
        .dout(new_Jinkela_wire_8069)
    );

    bfr new_Jinkela_buffer_4104 (
        .din(new_Jinkela_wire_4804),
        .dout(new_Jinkela_wire_4805)
    );

    bfr new_Jinkela_buffer_28 (
        .din(new_Jinkela_wire_29),
        .dout(new_Jinkela_wire_30)
    );

    spl4L new_Jinkela_splitter_53 (
        .a(new_Jinkela_wire_1228),
        .d(new_Jinkela_wire_1229),
        .b(new_Jinkela_wire_1230),
        .e(new_Jinkela_wire_1231),
        .c(new_Jinkela_wire_1232)
    );

    bfr new_Jinkela_buffer_4190 (
        .din(new_Jinkela_wire_4919),
        .dout(new_Jinkela_wire_4920)
    );

    bfr new_Jinkela_buffer_91 (
        .din(new_Jinkela_wire_98),
        .dout(new_Jinkela_wire_99)
    );

    bfr new_Jinkela_buffer_1070 (
        .din(new_Jinkela_wire_1146),
        .dout(new_Jinkela_wire_1147)
    );

    bfr new_Jinkela_buffer_4128 (
        .din(new_Jinkela_wire_4828),
        .dout(new_Jinkela_wire_4829)
    );

    bfr new_Jinkela_buffer_4105 (
        .din(new_Jinkela_wire_4805),
        .dout(new_Jinkela_wire_4806)
    );

    bfr new_Jinkela_buffer_29 (
        .din(new_Jinkela_wire_30),
        .dout(new_Jinkela_wire_31)
    );

    spl4L new_Jinkela_splitter_56 (
        .a(new_Jinkela_wire_1243),
        .d(new_Jinkela_wire_1244),
        .b(new_Jinkela_wire_1249),
        .e(new_Jinkela_wire_1254),
        .c(new_Jinkela_wire_1259)
    );

    bfr new_Jinkela_buffer_94 (
        .din(new_Jinkela_wire_101),
        .dout(new_Jinkela_wire_102)
    );

    bfr new_Jinkela_buffer_1071 (
        .din(new_Jinkela_wire_1147),
        .dout(new_Jinkela_wire_1148)
    );

    bfr new_Jinkela_buffer_4154 (
        .din(new_Jinkela_wire_4866),
        .dout(new_Jinkela_wire_4867)
    );

    bfr new_Jinkela_buffer_4106 (
        .din(new_Jinkela_wire_4806),
        .dout(new_Jinkela_wire_4807)
    );

    bfr new_Jinkela_buffer_30 (
        .din(new_Jinkela_wire_31),
        .dout(new_Jinkela_wire_32)
    );

    spl4L new_Jinkela_splitter_51 (
        .a(new_Jinkela_wire_1222),
        .d(new_Jinkela_wire_1223),
        .b(new_Jinkela_wire_1228),
        .e(new_Jinkela_wire_1233),
        .c(new_Jinkela_wire_1238)
    );

    bfr new_Jinkela_buffer_92 (
        .din(new_Jinkela_wire_99),
        .dout(new_Jinkela_wire_100)
    );

    bfr new_Jinkela_buffer_1072 (
        .din(new_Jinkela_wire_1148),
        .dout(new_Jinkela_wire_1149)
    );

    bfr new_Jinkela_buffer_4129 (
        .din(new_Jinkela_wire_4829),
        .dout(new_Jinkela_wire_4830)
    );

    bfr new_Jinkela_buffer_4107 (
        .din(new_Jinkela_wire_4807),
        .dout(new_Jinkela_wire_4808)
    );

    bfr new_Jinkela_buffer_31 (
        .din(new_Jinkela_wire_32),
        .dout(new_Jinkela_wire_33)
    );

    spl4L new_Jinkela_splitter_52 (
        .a(new_Jinkela_wire_1223),
        .d(new_Jinkela_wire_1224),
        .b(new_Jinkela_wire_1225),
        .e(new_Jinkela_wire_1226),
        .c(new_Jinkela_wire_1227)
    );

    bfr new_Jinkela_buffer_97 (
        .din(new_Jinkela_wire_106),
        .dout(new_Jinkela_wire_107)
    );

    bfr new_Jinkela_buffer_1073 (
        .din(new_Jinkela_wire_1149),
        .dout(new_Jinkela_wire_1150)
    );

    bfr new_Jinkela_buffer_4108 (
        .din(new_Jinkela_wire_4808),
        .dout(new_Jinkela_wire_4809)
    );

    bfr new_Jinkela_buffer_32 (
        .din(new_Jinkela_wire_33),
        .dout(new_Jinkela_wire_34)
    );

    spl4L new_Jinkela_splitter_57 (
        .a(new_Jinkela_wire_1244),
        .d(new_Jinkela_wire_1245),
        .b(new_Jinkela_wire_1246),
        .e(new_Jinkela_wire_1247),
        .c(new_Jinkela_wire_1248)
    );

    bfr new_Jinkela_buffer_95 (
        .din(new_Jinkela_wire_102),
        .dout(new_Jinkela_wire_103)
    );

    bfr new_Jinkela_buffer_1074 (
        .din(new_Jinkela_wire_1150),
        .dout(new_Jinkela_wire_1151)
    );

    bfr new_Jinkela_buffer_4130 (
        .din(new_Jinkela_wire_4830),
        .dout(new_Jinkela_wire_4831)
    );

    bfr new_Jinkela_buffer_4109 (
        .din(new_Jinkela_wire_4809),
        .dout(new_Jinkela_wire_4810)
    );

    bfr new_Jinkela_buffer_33 (
        .din(new_Jinkela_wire_34),
        .dout(new_Jinkela_wire_35)
    );

    spl4L new_Jinkela_splitter_54 (
        .a(new_Jinkela_wire_1233),
        .d(new_Jinkela_wire_1234),
        .b(new_Jinkela_wire_1235),
        .e(new_Jinkela_wire_1236),
        .c(new_Jinkela_wire_1237)
    );

    bfr new_Jinkela_buffer_162 (
        .din(new_Jinkela_wire_173),
        .dout(new_Jinkela_wire_174)
    );

    bfr new_Jinkela_buffer_165 (
        .din(N41),
        .dout(new_Jinkela_wire_177)
    );

    bfr new_Jinkela_buffer_1075 (
        .din(new_Jinkela_wire_1151),
        .dout(new_Jinkela_wire_1152)
    );

    bfr new_Jinkela_buffer_4155 (
        .din(new_Jinkela_wire_4867),
        .dout(new_Jinkela_wire_4868)
    );

    bfr new_Jinkela_buffer_4110 (
        .din(new_Jinkela_wire_4810),
        .dout(new_Jinkela_wire_4811)
    );

    bfr new_Jinkela_buffer_34 (
        .din(new_Jinkela_wire_35),
        .dout(new_Jinkela_wire_36)
    );

    spl4L new_Jinkela_splitter_55 (
        .a(new_Jinkela_wire_1238),
        .d(new_Jinkela_wire_1239),
        .b(new_Jinkela_wire_1240),
        .e(new_Jinkela_wire_1241),
        .c(new_Jinkela_wire_1242)
    );

    bfr new_Jinkela_buffer_96 (
        .din(new_Jinkela_wire_103),
        .dout(new_Jinkela_wire_104)
    );

    bfr new_Jinkela_buffer_1076 (
        .din(new_Jinkela_wire_1152),
        .dout(new_Jinkela_wire_1153)
    );

    bfr new_Jinkela_buffer_4131 (
        .din(new_Jinkela_wire_4831),
        .dout(new_Jinkela_wire_4832)
    );

    bfr new_Jinkela_buffer_4111 (
        .din(new_Jinkela_wire_4811),
        .dout(new_Jinkela_wire_4812)
    );

    bfr new_Jinkela_buffer_35 (
        .din(new_Jinkela_wire_36),
        .dout(new_Jinkela_wire_37)
    );

    spl4L new_Jinkela_splitter_61 (
        .a(new_Jinkela_wire_1264),
        .d(new_Jinkela_wire_1265),
        .b(new_Jinkela_wire_1270),
        .e(new_Jinkela_wire_1275),
        .c(new_Jinkela_wire_1280)
    );

    bfr new_Jinkela_buffer_168 (
        .din(N151),
        .dout(new_Jinkela_wire_182)
    );

    bfr new_Jinkela_buffer_1077 (
        .din(new_Jinkela_wire_1153),
        .dout(new_Jinkela_wire_1154)
    );

    spl3L new_Jinkela_splitter_270 (
        .a(n_1366_),
        .d(new_Jinkela_wire_4917),
        .b(new_Jinkela_wire_4918),
        .c(new_Jinkela_wire_4919)
    );

    bfr new_Jinkela_buffer_4112 (
        .din(new_Jinkela_wire_4812),
        .dout(new_Jinkela_wire_4813)
    );

    bfr new_Jinkela_buffer_36 (
        .din(new_Jinkela_wire_37),
        .dout(new_Jinkela_wire_38)
    );

    spl4L new_Jinkela_splitter_58 (
        .a(new_Jinkela_wire_1249),
        .d(new_Jinkela_wire_1250),
        .b(new_Jinkela_wire_1251),
        .e(new_Jinkela_wire_1252),
        .c(new_Jinkela_wire_1253)
    );

    spl3L new_Jinkela_splitter_267 (
        .a(new_Jinkela_wire_4875),
        .d(new_Jinkela_wire_4876),
        .b(new_Jinkela_wire_4877),
        .c(new_Jinkela_wire_4878)
    );

    bfr new_Jinkela_buffer_1078 (
        .din(new_Jinkela_wire_1154),
        .dout(new_Jinkela_wire_1155)
    );

    bfr new_Jinkela_buffer_4132 (
        .din(new_Jinkela_wire_4832),
        .dout(new_Jinkela_wire_4833)
    );

    bfr new_Jinkela_buffer_4113 (
        .din(new_Jinkela_wire_4813),
        .dout(new_Jinkela_wire_4814)
    );

    bfr new_Jinkela_buffer_37 (
        .din(new_Jinkela_wire_38),
        .dout(new_Jinkela_wire_39)
    );

    spl4L new_Jinkela_splitter_62 (
        .a(new_Jinkela_wire_1265),
        .d(new_Jinkela_wire_1266),
        .b(new_Jinkela_wire_1267),
        .e(new_Jinkela_wire_1268),
        .c(new_Jinkela_wire_1269)
    );

    bfr new_Jinkela_buffer_98 (
        .din(new_Jinkela_wire_107),
        .dout(new_Jinkela_wire_108)
    );

    bfr new_Jinkela_buffer_1079 (
        .din(new_Jinkela_wire_1155),
        .dout(new_Jinkela_wire_1156)
    );

    spl2 new_Jinkela_splitter_265 (
        .a(new_Jinkela_wire_4868),
        .b(new_Jinkela_wire_4869),
        .c(new_Jinkela_wire_4870)
    );

    bfr new_Jinkela_buffer_4114 (
        .din(new_Jinkela_wire_4814),
        .dout(new_Jinkela_wire_4815)
    );

    bfr new_Jinkela_buffer_38 (
        .din(new_Jinkela_wire_39),
        .dout(new_Jinkela_wire_40)
    );

    spl4L new_Jinkela_splitter_59 (
        .a(new_Jinkela_wire_1254),
        .d(new_Jinkela_wire_1255),
        .b(new_Jinkela_wire_1256),
        .e(new_Jinkela_wire_1257),
        .c(new_Jinkela_wire_1258)
    );

    bfr new_Jinkela_buffer_1080 (
        .din(new_Jinkela_wire_1156),
        .dout(new_Jinkela_wire_1157)
    );

    bfr new_Jinkela_buffer_4133 (
        .din(new_Jinkela_wire_4833),
        .dout(new_Jinkela_wire_4834)
    );

    bfr new_Jinkela_buffer_4115 (
        .din(new_Jinkela_wire_4815),
        .dout(new_Jinkela_wire_4816)
    );

    bfr new_Jinkela_buffer_39 (
        .din(new_Jinkela_wire_40),
        .dout(new_Jinkela_wire_41)
    );

    spl4L new_Jinkela_splitter_60 (
        .a(new_Jinkela_wire_1259),
        .d(new_Jinkela_wire_1260),
        .b(new_Jinkela_wire_1261),
        .e(new_Jinkela_wire_1262),
        .c(new_Jinkela_wire_1263)
    );

    spl2 new_Jinkela_splitter_4 (
        .a(new_Jinkela_wire_108),
        .b(new_Jinkela_wire_109),
        .c(new_Jinkela_wire_110)
    );

    bfr new_Jinkela_buffer_1081 (
        .din(new_Jinkela_wire_1157),
        .dout(new_Jinkela_wire_1158)
    );

    bfr new_Jinkela_buffer_4116 (
        .din(new_Jinkela_wire_4816),
        .dout(new_Jinkela_wire_4817)
    );

    bfr new_Jinkela_buffer_40 (
        .din(new_Jinkela_wire_41),
        .dout(new_Jinkela_wire_42)
    );

    spl4L new_Jinkela_splitter_66 (
        .a(new_Jinkela_wire_1285),
        .d(new_Jinkela_wire_1286),
        .b(new_Jinkela_wire_1291),
        .e(new_Jinkela_wire_1296),
        .c(new_Jinkela_wire_1301)
    );

    bfr new_Jinkela_buffer_99 (
        .din(new_Jinkela_wire_110),
        .dout(new_Jinkela_wire_111)
    );

    bfr new_Jinkela_buffer_1082 (
        .din(new_Jinkela_wire_1158),
        .dout(new_Jinkela_wire_1159)
    );

    bfr new_Jinkela_buffer_4134 (
        .din(new_Jinkela_wire_4834),
        .dout(new_Jinkela_wire_4835)
    );

    bfr new_Jinkela_buffer_41 (
        .din(new_Jinkela_wire_42),
        .dout(new_Jinkela_wire_43)
    );

    spl4L new_Jinkela_splitter_63 (
        .a(new_Jinkela_wire_1270),
        .d(new_Jinkela_wire_1271),
        .b(new_Jinkela_wire_1272),
        .e(new_Jinkela_wire_1273),
        .c(new_Jinkela_wire_1274)
    );

    spl2 new_Jinkela_splitter_274 (
        .a(n_0747_),
        .b(new_Jinkela_wire_4963),
        .c(new_Jinkela_wire_4964)
    );

    bfr new_Jinkela_buffer_4157 (
        .din(new_Jinkela_wire_4878),
        .dout(new_Jinkela_wire_4879)
    );

    bfr new_Jinkela_buffer_163 (
        .din(new_Jinkela_wire_174),
        .dout(new_Jinkela_wire_175)
    );

    bfr new_Jinkela_buffer_1083 (
        .din(new_Jinkela_wire_1159),
        .dout(new_Jinkela_wire_1160)
    );

    bfr new_Jinkela_buffer_4135 (
        .din(new_Jinkela_wire_4835),
        .dout(new_Jinkela_wire_4836)
    );

    bfr new_Jinkela_buffer_42 (
        .din(new_Jinkela_wire_43),
        .dout(new_Jinkela_wire_44)
    );

    spl4L new_Jinkela_splitter_67 (
        .a(new_Jinkela_wire_1286),
        .d(new_Jinkela_wire_1287),
        .b(new_Jinkela_wire_1288),
        .e(new_Jinkela_wire_1289),
        .c(new_Jinkela_wire_1290)
    );

    bfr new_Jinkela_buffer_4158 (
        .din(new_Jinkela_wire_4879),
        .dout(new_Jinkela_wire_4880)
    );

    spl2 new_Jinkela_splitter_6 (
        .a(N211),
        .b(new_Jinkela_wire_186),
        .c(new_Jinkela_wire_187)
    );

    bfr new_Jinkela_buffer_166 (
        .din(new_Jinkela_wire_177),
        .dout(new_Jinkela_wire_178)
    );

    bfr new_Jinkela_buffer_1084 (
        .din(new_Jinkela_wire_1160),
        .dout(new_Jinkela_wire_1161)
    );

    bfr new_Jinkela_buffer_4136 (
        .din(new_Jinkela_wire_4836),
        .dout(new_Jinkela_wire_4837)
    );

    bfr new_Jinkela_buffer_43 (
        .din(new_Jinkela_wire_44),
        .dout(new_Jinkela_wire_45)
    );

    spl4L new_Jinkela_splitter_64 (
        .a(new_Jinkela_wire_1275),
        .d(new_Jinkela_wire_1276),
        .b(new_Jinkela_wire_1277),
        .e(new_Jinkela_wire_1278),
        .c(new_Jinkela_wire_1279)
    );

    bfr new_Jinkela_buffer_100 (
        .din(new_Jinkela_wire_111),
        .dout(new_Jinkela_wire_112)
    );

    bfr new_Jinkela_buffer_1085 (
        .din(new_Jinkela_wire_1161),
        .dout(new_Jinkela_wire_1162)
    );

    bfr new_Jinkela_buffer_4137 (
        .din(new_Jinkela_wire_4837),
        .dout(new_Jinkela_wire_4838)
    );

    bfr new_Jinkela_buffer_44 (
        .din(new_Jinkela_wire_45),
        .dout(new_Jinkela_wire_46)
    );

    spl4L new_Jinkela_splitter_65 (
        .a(new_Jinkela_wire_1280),
        .d(new_Jinkela_wire_1281),
        .b(new_Jinkela_wire_1282),
        .e(new_Jinkela_wire_1283),
        .c(new_Jinkela_wire_1284)
    );

    spl4L new_Jinkela_splitter_271 (
        .a(n_0178_),
        .d(new_Jinkela_wire_4921),
        .b(new_Jinkela_wire_4922),
        .e(new_Jinkela_wire_4923),
        .c(new_Jinkela_wire_4924)
    );

    bfr new_Jinkela_buffer_4159 (
        .din(new_Jinkela_wire_4880),
        .dout(new_Jinkela_wire_4881)
    );

    bfr new_Jinkela_buffer_164 (
        .din(new_Jinkela_wire_175),
        .dout(new_Jinkela_wire_176)
    );

    bfr new_Jinkela_buffer_1086 (
        .din(new_Jinkela_wire_1162),
        .dout(new_Jinkela_wire_1163)
    );

    bfr new_Jinkela_buffer_4138 (
        .din(new_Jinkela_wire_4838),
        .dout(new_Jinkela_wire_4839)
    );

    bfr new_Jinkela_buffer_45 (
        .din(new_Jinkela_wire_46),
        .dout(new_Jinkela_wire_47)
    );

    bfr new_Jinkela_buffer_1164 (
        .din(new_Jinkela_wire_1477),
        .dout(new_Jinkela_wire_1478)
    );

    bfr new_Jinkela_buffer_101 (
        .din(new_Jinkela_wire_112),
        .dout(new_Jinkela_wire_113)
    );

    bfr new_Jinkela_buffer_4191 (
        .din(new_net_2541),
        .dout(new_Jinkela_wire_4925)
    );

    bfr new_Jinkela_buffer_1087 (
        .din(new_Jinkela_wire_1163),
        .dout(new_Jinkela_wire_1164)
    );

    bfr new_Jinkela_buffer_4139 (
        .din(new_Jinkela_wire_4839),
        .dout(new_Jinkela_wire_4840)
    );

    bfr new_Jinkela_buffer_46 (
        .din(new_Jinkela_wire_47),
        .dout(new_Jinkela_wire_48)
    );

    spl4L new_Jinkela_splitter_68 (
        .a(new_Jinkela_wire_1291),
        .d(new_Jinkela_wire_1292),
        .b(new_Jinkela_wire_1293),
        .e(new_Jinkela_wire_1294),
        .c(new_Jinkela_wire_1295)
    );

    bfr new_Jinkela_buffer_4192 (
        .din(new_Jinkela_wire_4925),
        .dout(new_Jinkela_wire_4926)
    );

    bfr new_Jinkela_buffer_4160 (
        .din(new_Jinkela_wire_4881),
        .dout(new_Jinkela_wire_4882)
    );

    bfr new_Jinkela_buffer_172 (
        .din(N175),
        .dout(new_Jinkela_wire_188)
    );

    bfr new_Jinkela_buffer_4140 (
        .din(new_Jinkela_wire_4840),
        .dout(new_Jinkela_wire_4841)
    );

    spl4L new_Jinkela_splitter_74 (
        .a(new_Jinkela_wire_1313),
        .d(new_Jinkela_wire_1314),
        .b(new_Jinkela_wire_1315),
        .e(new_Jinkela_wire_1316),
        .c(new_Jinkela_wire_1317)
    );

    bfr new_Jinkela_buffer_47 (
        .din(new_Jinkela_wire_48),
        .dout(new_Jinkela_wire_49)
    );

    spl4L new_Jinkela_splitter_69 (
        .a(new_Jinkela_wire_1296),
        .d(new_Jinkela_wire_1297),
        .b(new_Jinkela_wire_1298),
        .e(new_Jinkela_wire_1299),
        .c(new_Jinkela_wire_1300)
    );

    bfr new_Jinkela_buffer_102 (
        .din(new_Jinkela_wire_113),
        .dout(new_Jinkela_wire_114)
    );

    spl4L new_Jinkela_splitter_70 (
        .a(new_Jinkela_wire_1301),
        .d(new_Jinkela_wire_1302),
        .b(new_Jinkela_wire_1303),
        .e(new_Jinkela_wire_1304),
        .c(new_Jinkela_wire_1305)
    );

    bfr new_Jinkela_buffer_4141 (
        .din(new_Jinkela_wire_4841),
        .dout(new_Jinkela_wire_4842)
    );

    bfr new_Jinkela_buffer_48 (
        .din(new_Jinkela_wire_49),
        .dout(new_Jinkela_wire_50)
    );

    spl4L new_Jinkela_splitter_77 (
        .a(new_Jinkela_wire_1328),
        .d(new_Jinkela_wire_1329),
        .b(new_Jinkela_wire_1334),
        .e(new_Jinkela_wire_1339),
        .c(new_Jinkela_wire_1344)
    );

    spl3L new_Jinkela_splitter_272 (
        .a(n_0621_),
        .d(new_Jinkela_wire_4957),
        .b(new_Jinkela_wire_4958),
        .c(new_Jinkela_wire_4959)
    );

    bfr new_Jinkela_buffer_4161 (
        .din(new_Jinkela_wire_4882),
        .dout(new_Jinkela_wire_4883)
    );

    bfr new_Jinkela_buffer_169 (
        .din(new_Jinkela_wire_182),
        .dout(new_Jinkela_wire_183)
    );

    bfr new_Jinkela_buffer_167 (
        .din(new_Jinkela_wire_178),
        .dout(new_Jinkela_wire_179)
    );

    spl4L new_Jinkela_splitter_72 (
        .a(new_Jinkela_wire_1307),
        .d(new_Jinkela_wire_1308),
        .b(new_Jinkela_wire_1313),
        .e(new_Jinkela_wire_1318),
        .c(new_Jinkela_wire_1323)
    );

    bfr new_Jinkela_buffer_4142 (
        .din(new_Jinkela_wire_4842),
        .dout(new_Jinkela_wire_4843)
    );

    bfr new_Jinkela_buffer_4967 (
        .din(new_Jinkela_wire_5916),
        .dout(new_Jinkela_wire_5917)
    );

    bfr new_Jinkela_buffer_4931 (
        .din(new_Jinkela_wire_5867),
        .dout(new_Jinkela_wire_5868)
    );

    bfr new_Jinkela_buffer_5783 (
        .din(new_Jinkela_wire_6976),
        .dout(new_Jinkela_wire_6977)
    );

    spl3L new_Jinkela_splitter_367 (
        .a(n_1334_),
        .d(new_Jinkela_wire_5979),
        .b(new_Jinkela_wire_5980),
        .c(new_Jinkela_wire_5981)
    );

    spl3L new_Jinkela_splitter_357 (
        .a(new_Jinkela_wire_5868),
        .d(new_Jinkela_wire_5869),
        .b(new_Jinkela_wire_5870),
        .c(new_Jinkela_wire_5871)
    );

    bfr new_Jinkela_buffer_5784 (
        .din(new_Jinkela_wire_6977),
        .dout(new_Jinkela_wire_6978)
    );

    spl3L new_Jinkela_splitter_370 (
        .a(n_0975_),
        .d(new_Jinkela_wire_6008),
        .b(new_Jinkela_wire_6009),
        .c(new_Jinkela_wire_6010)
    );

    bfr new_Jinkela_buffer_5831 (
        .din(new_Jinkela_wire_7035),
        .dout(new_Jinkela_wire_7036)
    );

    bfr new_Jinkela_buffer_4983 (
        .din(new_Jinkela_wire_5940),
        .dout(new_Jinkela_wire_5941)
    );

    bfr new_Jinkela_buffer_5785 (
        .din(new_Jinkela_wire_6978),
        .dout(new_Jinkela_wire_6979)
    );

    bfr new_Jinkela_buffer_5013 (
        .din(new_Jinkela_wire_5972),
        .dout(new_Jinkela_wire_5973)
    );

    bfr new_Jinkela_buffer_5865 (
        .din(new_Jinkela_wire_7087),
        .dout(new_Jinkela_wire_7088)
    );

    bfr new_Jinkela_buffer_5864 (
        .din(new_Jinkela_wire_7084),
        .dout(new_Jinkela_wire_7085)
    );

    bfr new_Jinkela_buffer_4984 (
        .din(new_Jinkela_wire_5941),
        .dout(new_Jinkela_wire_5942)
    );

    bfr new_Jinkela_buffer_5786 (
        .din(new_Jinkela_wire_6979),
        .dout(new_Jinkela_wire_6980)
    );

    bfr new_Jinkela_buffer_5832 (
        .din(new_Jinkela_wire_7036),
        .dout(new_Jinkela_wire_7037)
    );

    bfr new_Jinkela_buffer_4985 (
        .din(new_Jinkela_wire_5942),
        .dout(new_Jinkela_wire_5943)
    );

    bfr new_Jinkela_buffer_5787 (
        .din(new_Jinkela_wire_6980),
        .dout(new_Jinkela_wire_6981)
    );

    bfr new_Jinkela_buffer_5014 (
        .din(new_Jinkela_wire_5973),
        .dout(new_Jinkela_wire_5974)
    );

    bfr new_Jinkela_buffer_4986 (
        .din(new_Jinkela_wire_5943),
        .dout(new_Jinkela_wire_5944)
    );

    bfr new_Jinkela_buffer_5788 (
        .din(new_Jinkela_wire_6981),
        .dout(new_Jinkela_wire_6982)
    );

    spl2 new_Jinkela_splitter_373 (
        .a(n_0106_),
        .b(new_Jinkela_wire_6016),
        .c(new_Jinkela_wire_6017)
    );

    bfr new_Jinkela_buffer_5833 (
        .din(new_Jinkela_wire_7037),
        .dout(new_Jinkela_wire_7038)
    );

    bfr new_Jinkela_buffer_4987 (
        .din(new_Jinkela_wire_5944),
        .dout(new_Jinkela_wire_5945)
    );

    bfr new_Jinkela_buffer_5789 (
        .din(new_Jinkela_wire_6982),
        .dout(new_Jinkela_wire_6983)
    );

    bfr new_Jinkela_buffer_5015 (
        .din(new_Jinkela_wire_5974),
        .dout(new_Jinkela_wire_5975)
    );

    spl3L new_Jinkela_splitter_478 (
        .a(n_1075_),
        .d(new_Jinkela_wire_7092),
        .b(new_Jinkela_wire_7093),
        .c(new_Jinkela_wire_7094)
    );

    bfr new_Jinkela_buffer_4988 (
        .din(new_Jinkela_wire_5945),
        .dout(new_Jinkela_wire_5946)
    );

    bfr new_Jinkela_buffer_5790 (
        .din(new_Jinkela_wire_6983),
        .dout(new_Jinkela_wire_6984)
    );

    bfr new_Jinkela_buffer_5019 (
        .din(new_Jinkela_wire_5981),
        .dout(new_Jinkela_wire_5982)
    );

    bfr new_Jinkela_buffer_5834 (
        .din(new_Jinkela_wire_7038),
        .dout(new_Jinkela_wire_7039)
    );

    bfr new_Jinkela_buffer_4989 (
        .din(new_Jinkela_wire_5946),
        .dout(new_Jinkela_wire_5947)
    );

    bfr new_Jinkela_buffer_5791 (
        .din(new_Jinkela_wire_6984),
        .dout(new_Jinkela_wire_6985)
    );

    bfr new_Jinkela_buffer_5016 (
        .din(new_Jinkela_wire_5975),
        .dout(new_Jinkela_wire_5976)
    );

    spl2 new_Jinkela_splitter_480 (
        .a(n_0044_),
        .b(new_Jinkela_wire_7097),
        .c(new_Jinkela_wire_7098)
    );

    spl2 new_Jinkela_splitter_479 (
        .a(new_Jinkela_wire_7094),
        .b(new_Jinkela_wire_7095),
        .c(new_Jinkela_wire_7096)
    );

    bfr new_Jinkela_buffer_4990 (
        .din(new_Jinkela_wire_5947),
        .dout(new_Jinkela_wire_5948)
    );

    bfr new_Jinkela_buffer_5792 (
        .din(new_Jinkela_wire_6985),
        .dout(new_Jinkela_wire_6986)
    );

    bfr new_Jinkela_buffer_5020 (
        .din(new_Jinkela_wire_5982),
        .dout(new_Jinkela_wire_5983)
    );

    bfr new_Jinkela_buffer_5835 (
        .din(new_Jinkela_wire_7039),
        .dout(new_Jinkela_wire_7040)
    );

    bfr new_Jinkela_buffer_4991 (
        .din(new_Jinkela_wire_5948),
        .dout(new_Jinkela_wire_5949)
    );

    bfr new_Jinkela_buffer_5793 (
        .din(new_Jinkela_wire_6986),
        .dout(new_Jinkela_wire_6987)
    );

    spl2 new_Jinkela_splitter_371 (
        .a(new_Jinkela_wire_6010),
        .b(new_Jinkela_wire_6011),
        .c(new_Jinkela_wire_6012)
    );

    spl3L new_Jinkela_splitter_482 (
        .a(n_1090_),
        .d(new_Jinkela_wire_7116),
        .b(new_Jinkela_wire_7117),
        .c(new_Jinkela_wire_7118)
    );

    spl2 new_Jinkela_splitter_481 (
        .a(n_1345_),
        .b(new_Jinkela_wire_7114),
        .c(new_Jinkela_wire_7115)
    );

    bfr new_Jinkela_buffer_4992 (
        .din(new_Jinkela_wire_5949),
        .dout(new_Jinkela_wire_5950)
    );

    bfr new_Jinkela_buffer_5794 (
        .din(new_Jinkela_wire_6987),
        .dout(new_Jinkela_wire_6988)
    );

    spl2 new_Jinkela_splitter_372 (
        .a(n_0296_),
        .b(new_Jinkela_wire_6013),
        .c(new_Jinkela_wire_6014)
    );

    bfr new_Jinkela_buffer_5041 (
        .din(new_Jinkela_wire_6014),
        .dout(new_Jinkela_wire_6015)
    );

    bfr new_Jinkela_buffer_5836 (
        .din(new_Jinkela_wire_7040),
        .dout(new_Jinkela_wire_7041)
    );

    bfr new_Jinkela_buffer_4993 (
        .din(new_Jinkela_wire_5950),
        .dout(new_Jinkela_wire_5951)
    );

    bfr new_Jinkela_buffer_5795 (
        .din(new_Jinkela_wire_6988),
        .dout(new_Jinkela_wire_6989)
    );

    spl2 new_Jinkela_splitter_368 (
        .a(new_Jinkela_wire_5983),
        .b(new_Jinkela_wire_5984),
        .c(new_Jinkela_wire_5985)
    );

    bfr new_Jinkela_buffer_4994 (
        .din(new_Jinkela_wire_5951),
        .dout(new_Jinkela_wire_5952)
    );

    bfr new_Jinkela_buffer_5796 (
        .din(new_Jinkela_wire_6989),
        .dout(new_Jinkela_wire_6990)
    );

    bfr new_Jinkela_buffer_5021 (
        .din(new_Jinkela_wire_5985),
        .dout(new_Jinkela_wire_5986)
    );

    bfr new_Jinkela_buffer_5837 (
        .din(new_Jinkela_wire_7041),
        .dout(new_Jinkela_wire_7042)
    );

    bfr new_Jinkela_buffer_4995 (
        .din(new_Jinkela_wire_5952),
        .dout(new_Jinkela_wire_5953)
    );

    bfr new_Jinkela_buffer_5797 (
        .din(new_Jinkela_wire_6990),
        .dout(new_Jinkela_wire_6991)
    );

    bfr new_Jinkela_buffer_4996 (
        .din(new_Jinkela_wire_5953),
        .dout(new_Jinkela_wire_5954)
    );

    bfr new_Jinkela_buffer_5798 (
        .din(new_Jinkela_wire_6991),
        .dout(new_Jinkela_wire_6992)
    );

    spl2 new_Jinkela_splitter_374 (
        .a(n_0456_),
        .b(new_Jinkela_wire_6059),
        .c(new_Jinkela_wire_6060)
    );

    bfr new_Jinkela_buffer_5042 (
        .din(new_Jinkela_wire_6017),
        .dout(new_Jinkela_wire_6018)
    );

    bfr new_Jinkela_buffer_5838 (
        .din(new_Jinkela_wire_7042),
        .dout(new_Jinkela_wire_7043)
    );

    bfr new_Jinkela_buffer_4997 (
        .din(new_Jinkela_wire_5954),
        .dout(new_Jinkela_wire_5955)
    );

    bfr new_Jinkela_buffer_5799 (
        .din(new_Jinkela_wire_6992),
        .dout(new_Jinkela_wire_6993)
    );

    bfr new_Jinkela_buffer_5022 (
        .din(new_Jinkela_wire_5986),
        .dout(new_Jinkela_wire_5987)
    );

    bfr new_Jinkela_buffer_5866 (
        .din(new_Jinkela_wire_7098),
        .dout(new_Jinkela_wire_7099)
    );

    bfr new_Jinkela_buffer_4998 (
        .din(new_Jinkela_wire_5955),
        .dout(new_Jinkela_wire_5956)
    );

    bfr new_Jinkela_buffer_5800 (
        .din(new_Jinkela_wire_6993),
        .dout(new_Jinkela_wire_6994)
    );

    bfr new_Jinkela_buffer_5083 (
        .din(n_0497_),
        .dout(new_Jinkela_wire_6061)
    );

    bfr new_Jinkela_buffer_5839 (
        .din(new_Jinkela_wire_7043),
        .dout(new_Jinkela_wire_7044)
    );

    bfr new_Jinkela_buffer_4999 (
        .din(new_Jinkela_wire_5956),
        .dout(new_Jinkela_wire_5957)
    );

    bfr new_Jinkela_buffer_5801 (
        .din(new_Jinkela_wire_6994),
        .dout(new_Jinkela_wire_6995)
    );

    bfr new_Jinkela_buffer_5023 (
        .din(new_Jinkela_wire_5987),
        .dout(new_Jinkela_wire_5988)
    );

    bfr new_Jinkela_buffer_5881 (
        .din(new_net_2562),
        .dout(new_Jinkela_wire_7121)
    );

    bfr new_Jinkela_buffer_5000 (
        .din(new_Jinkela_wire_5957),
        .dout(new_Jinkela_wire_5958)
    );

    bfr new_Jinkela_buffer_5802 (
        .din(new_Jinkela_wire_6995),
        .dout(new_Jinkela_wire_6996)
    );

    spl2 new_Jinkela_splitter_375 (
        .a(n_1328_),
        .b(new_Jinkela_wire_6087),
        .c(new_Jinkela_wire_6088)
    );

    bfr new_Jinkela_buffer_5840 (
        .din(new_Jinkela_wire_7044),
        .dout(new_Jinkela_wire_7045)
    );

    bfr new_Jinkela_buffer_5001 (
        .din(new_Jinkela_wire_5958),
        .dout(new_Jinkela_wire_5959)
    );

    bfr new_Jinkela_buffer_5803 (
        .din(new_Jinkela_wire_6996),
        .dout(new_Jinkela_wire_6997)
    );

    bfr new_Jinkela_buffer_5024 (
        .din(new_Jinkela_wire_5988),
        .dout(new_Jinkela_wire_5989)
    );

    bfr new_Jinkela_buffer_5867 (
        .din(new_Jinkela_wire_7099),
        .dout(new_Jinkela_wire_7100)
    );

    bfr new_Jinkela_buffer_1585 (
        .din(new_Jinkela_wire_1928),
        .dout(new_Jinkela_wire_1929)
    );

    bfr new_Jinkela_buffer_2427 (
        .din(new_Jinkela_wire_2828),
        .dout(new_Jinkela_wire_2829)
    );

    spl2 new_Jinkela_splitter_178 (
        .a(n_1205_),
        .b(new_Jinkela_wire_3838),
        .c(new_Jinkela_wire_3839)
    );

    bfr new_Jinkela_buffer_1543 (
        .din(new_Jinkela_wire_1880),
        .dout(new_Jinkela_wire_1881)
    );

    bfr new_Jinkela_buffer_2373 (
        .din(new_Jinkela_wire_2769),
        .dout(new_Jinkela_wire_2770)
    );

    bfr new_Jinkela_buffer_3268 (
        .din(new_Jinkela_wire_3756),
        .dout(new_Jinkela_wire_3757)
    );

    bfr new_Jinkela_buffer_1649 (
        .din(new_Jinkela_wire_1992),
        .dout(new_Jinkela_wire_1993)
    );

    bfr new_Jinkela_buffer_2491 (
        .din(new_Jinkela_wire_2892),
        .dout(new_Jinkela_wire_2893)
    );

    bfr new_Jinkela_buffer_3316 (
        .din(new_Jinkela_wire_3824),
        .dout(new_Jinkela_wire_3825)
    );

    bfr new_Jinkela_buffer_3290 (
        .din(new_Jinkela_wire_3798),
        .dout(new_Jinkela_wire_3799)
    );

    bfr new_Jinkela_buffer_1544 (
        .din(new_Jinkela_wire_1881),
        .dout(new_Jinkela_wire_1882)
    );

    bfr new_Jinkela_buffer_2374 (
        .din(new_Jinkela_wire_2770),
        .dout(new_Jinkela_wire_2771)
    );

    bfr new_Jinkela_buffer_3269 (
        .din(new_Jinkela_wire_3757),
        .dout(new_Jinkela_wire_3758)
    );

    bfr new_Jinkela_buffer_1586 (
        .din(new_Jinkela_wire_1929),
        .dout(new_Jinkela_wire_1930)
    );

    bfr new_Jinkela_buffer_2428 (
        .din(new_Jinkela_wire_2829),
        .dout(new_Jinkela_wire_2830)
    );

    bfr new_Jinkela_buffer_1545 (
        .din(new_Jinkela_wire_1882),
        .dout(new_Jinkela_wire_1883)
    );

    bfr new_Jinkela_buffer_2375 (
        .din(new_Jinkela_wire_2771),
        .dout(new_Jinkela_wire_2772)
    );

    bfr new_Jinkela_buffer_3270 (
        .din(new_Jinkela_wire_3758),
        .dout(new_Jinkela_wire_3759)
    );

    bfr new_Jinkela_buffer_2500 (
        .din(N241_I),
        .dout(new_Jinkela_wire_2902)
    );

    bfr new_Jinkela_buffer_3291 (
        .din(new_Jinkela_wire_3799),
        .dout(new_Jinkela_wire_3800)
    );

    bfr new_Jinkela_buffer_1546 (
        .din(new_Jinkela_wire_1883),
        .dout(new_Jinkela_wire_1884)
    );

    bfr new_Jinkela_buffer_2376 (
        .din(new_Jinkela_wire_2772),
        .dout(new_Jinkela_wire_2773)
    );

    bfr new_Jinkela_buffer_3271 (
        .din(new_Jinkela_wire_3759),
        .dout(new_Jinkela_wire_3760)
    );

    bfr new_Jinkela_buffer_1587 (
        .din(new_Jinkela_wire_1930),
        .dout(new_Jinkela_wire_1931)
    );

    bfr new_Jinkela_buffer_2429 (
        .din(new_Jinkela_wire_2830),
        .dout(new_Jinkela_wire_2831)
    );

    bfr new_Jinkela_buffer_1547 (
        .din(new_Jinkela_wire_1884),
        .dout(new_Jinkela_wire_1885)
    );

    bfr new_Jinkela_buffer_2377 (
        .din(new_Jinkela_wire_2773),
        .dout(new_Jinkela_wire_2774)
    );

    bfr new_Jinkela_buffer_3272 (
        .din(new_Jinkela_wire_3760),
        .dout(new_Jinkela_wire_3761)
    );

    bfr new_Jinkela_buffer_1652 (
        .din(new_Jinkela_wire_1995),
        .dout(new_Jinkela_wire_1996)
    );

    bfr new_Jinkela_buffer_2494 (
        .din(new_Jinkela_wire_2895),
        .dout(new_Jinkela_wire_2896)
    );

    bfr new_Jinkela_buffer_3317 (
        .din(new_Jinkela_wire_3825),
        .dout(new_Jinkela_wire_3826)
    );

    bfr new_Jinkela_buffer_3292 (
        .din(new_Jinkela_wire_3800),
        .dout(new_Jinkela_wire_3801)
    );

    bfr new_Jinkela_buffer_1548 (
        .din(new_Jinkela_wire_1885),
        .dout(new_Jinkela_wire_1886)
    );

    bfr new_Jinkela_buffer_2378 (
        .din(new_Jinkela_wire_2774),
        .dout(new_Jinkela_wire_2775)
    );

    bfr new_Jinkela_buffer_3273 (
        .din(new_Jinkela_wire_3761),
        .dout(new_Jinkela_wire_3762)
    );

    bfr new_Jinkela_buffer_1588 (
        .din(new_Jinkela_wire_1931),
        .dout(new_Jinkela_wire_1932)
    );

    bfr new_Jinkela_buffer_2430 (
        .din(new_Jinkela_wire_2831),
        .dout(new_Jinkela_wire_2832)
    );

    bfr new_Jinkela_buffer_1549 (
        .din(new_Jinkela_wire_1886),
        .dout(new_Jinkela_wire_1887)
    );

    bfr new_Jinkela_buffer_2379 (
        .din(new_Jinkela_wire_2775),
        .dout(new_Jinkela_wire_2776)
    );

    bfr new_Jinkela_buffer_3274 (
        .din(new_Jinkela_wire_3762),
        .dout(new_Jinkela_wire_3763)
    );

    bfr new_Jinkela_buffer_1723 (
        .din(N226),
        .dout(new_Jinkela_wire_2069)
    );

    bfr new_Jinkela_buffer_2497 (
        .din(new_Jinkela_wire_2898),
        .dout(new_Jinkela_wire_2899)
    );

    bfr new_Jinkela_buffer_1655 (
        .din(new_Jinkela_wire_1998),
        .dout(new_Jinkela_wire_1999)
    );

    bfr new_Jinkela_buffer_3293 (
        .din(new_Jinkela_wire_3801),
        .dout(new_Jinkela_wire_3802)
    );

    bfr new_Jinkela_buffer_1550 (
        .din(new_Jinkela_wire_1887),
        .dout(new_Jinkela_wire_1888)
    );

    bfr new_Jinkela_buffer_2380 (
        .din(new_Jinkela_wire_2776),
        .dout(new_Jinkela_wire_2777)
    );

    spl2 new_Jinkela_splitter_169 (
        .a(new_Jinkela_wire_3763),
        .b(new_Jinkela_wire_3764),
        .c(new_Jinkela_wire_3765)
    );

    bfr new_Jinkela_buffer_1589 (
        .din(new_Jinkela_wire_1932),
        .dout(new_Jinkela_wire_1933)
    );

    bfr new_Jinkela_buffer_2431 (
        .din(new_Jinkela_wire_2832),
        .dout(new_Jinkela_wire_2833)
    );

    bfr new_Jinkela_buffer_3275 (
        .din(new_Jinkela_wire_3765),
        .dout(new_Jinkela_wire_3766)
    );

    bfr new_Jinkela_buffer_1551 (
        .din(new_Jinkela_wire_1888),
        .dout(new_Jinkela_wire_1889)
    );

    bfr new_Jinkela_buffer_2381 (
        .din(new_Jinkela_wire_2777),
        .dout(new_Jinkela_wire_2778)
    );

    spl2 new_Jinkela_splitter_179 (
        .a(n_0271_),
        .b(new_Jinkela_wire_3842),
        .c(new_Jinkela_wire_3843)
    );

    bfr new_Jinkela_buffer_1653 (
        .din(new_Jinkela_wire_1996),
        .dout(new_Jinkela_wire_1997)
    );

    bfr new_Jinkela_buffer_2495 (
        .din(new_Jinkela_wire_2896),
        .dout(new_Jinkela_wire_2897)
    );

    bfr new_Jinkela_buffer_3318 (
        .din(new_Jinkela_wire_3826),
        .dout(new_Jinkela_wire_3827)
    );

    bfr new_Jinkela_buffer_3294 (
        .din(new_Jinkela_wire_3802),
        .dout(new_Jinkela_wire_3803)
    );

    bfr new_Jinkela_buffer_1552 (
        .din(new_Jinkela_wire_1889),
        .dout(new_Jinkela_wire_1890)
    );

    bfr new_Jinkela_buffer_2382 (
        .din(new_Jinkela_wire_2778),
        .dout(new_Jinkela_wire_2779)
    );

    spl2 new_Jinkela_splitter_170 (
        .a(new_Jinkela_wire_3766),
        .b(new_Jinkela_wire_3767),
        .c(new_Jinkela_wire_3768)
    );

    bfr new_Jinkela_buffer_1590 (
        .din(new_Jinkela_wire_1933),
        .dout(new_Jinkela_wire_1934)
    );

    bfr new_Jinkela_buffer_2432 (
        .din(new_Jinkela_wire_2833),
        .dout(new_Jinkela_wire_2834)
    );

    bfr new_Jinkela_buffer_3327 (
        .din(new_Jinkela_wire_3839),
        .dout(new_Jinkela_wire_3840)
    );

    bfr new_Jinkela_buffer_3295 (
        .din(new_Jinkela_wire_3803),
        .dout(new_Jinkela_wire_3804)
    );

    bfr new_Jinkela_buffer_1553 (
        .din(new_Jinkela_wire_1890),
        .dout(new_Jinkela_wire_1891)
    );

    bfr new_Jinkela_buffer_2383 (
        .din(new_Jinkela_wire_2779),
        .dout(new_Jinkela_wire_2780)
    );

    bfr new_Jinkela_buffer_2566 (
        .din(N187),
        .dout(new_Jinkela_wire_2968)
    );

    bfr new_Jinkela_buffer_1554 (
        .din(new_Jinkela_wire_1891),
        .dout(new_Jinkela_wire_1892)
    );

    bfr new_Jinkela_buffer_2384 (
        .din(new_Jinkela_wire_2780),
        .dout(new_Jinkela_wire_2781)
    );

    bfr new_Jinkela_buffer_3319 (
        .din(new_Jinkela_wire_3827),
        .dout(new_Jinkela_wire_3828)
    );

    bfr new_Jinkela_buffer_3296 (
        .din(new_Jinkela_wire_3804),
        .dout(new_Jinkela_wire_3805)
    );

    bfr new_Jinkela_buffer_1591 (
        .din(new_Jinkela_wire_1934),
        .dout(new_Jinkela_wire_1935)
    );

    bfr new_Jinkela_buffer_2433 (
        .din(new_Jinkela_wire_2834),
        .dout(new_Jinkela_wire_2835)
    );

    bfr new_Jinkela_buffer_1555 (
        .din(new_Jinkela_wire_1892),
        .dout(new_Jinkela_wire_1893)
    );

    bfr new_Jinkela_buffer_2385 (
        .din(new_Jinkela_wire_2781),
        .dout(new_Jinkela_wire_2782)
    );

    bfr new_Jinkela_buffer_3329 (
        .din(n_0290_),
        .dout(new_Jinkela_wire_3844)
    );

    bfr new_Jinkela_buffer_3297 (
        .din(new_Jinkela_wire_3805),
        .dout(new_Jinkela_wire_3806)
    );

    bfr new_Jinkela_buffer_1720 (
        .din(new_Jinkela_wire_2065),
        .dout(new_Jinkela_wire_2066)
    );

    bfr new_Jinkela_buffer_2498 (
        .din(new_Jinkela_wire_2899),
        .dout(new_Jinkela_wire_2900)
    );

    bfr new_Jinkela_buffer_1656 (
        .din(new_Jinkela_wire_1999),
        .dout(new_Jinkela_wire_2000)
    );

    bfr new_Jinkela_buffer_3330 (
        .din(new_Jinkela_wire_3844),
        .dout(new_Jinkela_wire_3845)
    );

    bfr new_Jinkela_buffer_1556 (
        .din(new_Jinkela_wire_1893),
        .dout(new_Jinkela_wire_1894)
    );

    bfr new_Jinkela_buffer_2386 (
        .din(new_Jinkela_wire_2782),
        .dout(new_Jinkela_wire_2783)
    );

    bfr new_Jinkela_buffer_3320 (
        .din(new_Jinkela_wire_3828),
        .dout(new_Jinkela_wire_3829)
    );

    bfr new_Jinkela_buffer_3298 (
        .din(new_Jinkela_wire_3806),
        .dout(new_Jinkela_wire_3807)
    );

    bfr new_Jinkela_buffer_1592 (
        .din(new_Jinkela_wire_1935),
        .dout(new_Jinkela_wire_1936)
    );

    bfr new_Jinkela_buffer_2434 (
        .din(new_Jinkela_wire_2835),
        .dout(new_Jinkela_wire_2836)
    );

    bfr new_Jinkela_buffer_1557 (
        .din(new_Jinkela_wire_1894),
        .dout(new_Jinkela_wire_1895)
    );

    bfr new_Jinkela_buffer_2387 (
        .din(new_Jinkela_wire_2783),
        .dout(new_Jinkela_wire_2784)
    );

    bfr new_Jinkela_buffer_3299 (
        .din(new_Jinkela_wire_3807),
        .dout(new_Jinkela_wire_3808)
    );

    bfr new_Jinkela_buffer_2501 (
        .din(new_Jinkela_wire_2902),
        .dout(new_Jinkela_wire_2903)
    );

    bfr new_Jinkela_buffer_3328 (
        .din(new_Jinkela_wire_3840),
        .dout(new_Jinkela_wire_3841)
    );

    bfr new_Jinkela_buffer_1558 (
        .din(new_Jinkela_wire_1895),
        .dout(new_Jinkela_wire_1896)
    );

    bfr new_Jinkela_buffer_2388 (
        .din(new_Jinkela_wire_2784),
        .dout(new_Jinkela_wire_2785)
    );

    bfr new_Jinkela_buffer_3321 (
        .din(new_Jinkela_wire_3829),
        .dout(new_Jinkela_wire_3830)
    );

    bfr new_Jinkela_buffer_3300 (
        .din(new_Jinkela_wire_3808),
        .dout(new_Jinkela_wire_3809)
    );

    bfr new_Jinkela_buffer_1593 (
        .din(new_Jinkela_wire_1936),
        .dout(new_Jinkela_wire_1937)
    );

    bfr new_Jinkela_buffer_2435 (
        .din(new_Jinkela_wire_2836),
        .dout(new_Jinkela_wire_2837)
    );

    bfr new_Jinkela_buffer_1559 (
        .din(new_Jinkela_wire_1896),
        .dout(new_Jinkela_wire_1897)
    );

    bfr new_Jinkela_buffer_2389 (
        .din(new_Jinkela_wire_2785),
        .dout(new_Jinkela_wire_2786)
    );

    bfr new_Jinkela_buffer_3301 (
        .din(new_Jinkela_wire_3809),
        .dout(new_Jinkela_wire_3810)
    );

    bfr new_Jinkela_buffer_1727 (
        .din(N77),
        .dout(new_Jinkela_wire_2073)
    );

    bfr new_Jinkela_buffer_2499 (
        .din(new_Jinkela_wire_2900),
        .dout(new_Jinkela_wire_2901)
    );

    spl2 new_Jinkela_splitter_109 (
        .a(new_Jinkela_wire_2000),
        .b(new_Jinkela_wire_2001),
        .c(new_Jinkela_wire_2002)
    );

    spl2 new_Jinkela_splitter_181 (
        .a(n_0764_),
        .b(new_Jinkela_wire_3853),
        .c(new_Jinkela_wire_3854)
    );

    bfr new_Jinkela_buffer_1560 (
        .din(new_Jinkela_wire_1897),
        .dout(new_Jinkela_wire_1898)
    );

    bfr new_Jinkela_buffer_2390 (
        .din(new_Jinkela_wire_2786),
        .dout(new_Jinkela_wire_2787)
    );

    bfr new_Jinkela_buffer_3322 (
        .din(new_Jinkela_wire_3830),
        .dout(new_Jinkela_wire_3831)
    );

    bfr new_Jinkela_buffer_3302 (
        .din(new_Jinkela_wire_3810),
        .dout(new_Jinkela_wire_3811)
    );

    bfr new_Jinkela_buffer_1594 (
        .din(new_Jinkela_wire_1937),
        .dout(new_Jinkela_wire_1938)
    );

    bfr new_Jinkela_buffer_2436 (
        .din(new_Jinkela_wire_2837),
        .dout(new_Jinkela_wire_2838)
    );

    bfr new_Jinkela_buffer_1561 (
        .din(new_Jinkela_wire_1898),
        .dout(new_Jinkela_wire_1899)
    );

    bfr new_Jinkela_buffer_2391 (
        .din(new_Jinkela_wire_2787),
        .dout(new_Jinkela_wire_2788)
    );

    spl2 new_Jinkela_splitter_180 (
        .a(n_0899_),
        .b(new_Jinkela_wire_3851),
        .c(new_Jinkela_wire_3852)
    );

    bfr new_Jinkela_buffer_3303 (
        .din(new_Jinkela_wire_3811),
        .dout(new_Jinkela_wire_3812)
    );

    bfr new_Jinkela_buffer_2570 (
        .din(N60),
        .dout(new_Jinkela_wire_2972)
    );

    bfr new_Jinkela_buffer_1657 (
        .din(new_Jinkela_wire_2002),
        .dout(new_Jinkela_wire_2003)
    );

    bfr new_Jinkela_buffer_1595 (
        .din(new_Jinkela_wire_1938),
        .dout(new_Jinkela_wire_1939)
    );

    bfr new_Jinkela_buffer_2392 (
        .din(new_Jinkela_wire_2788),
        .dout(new_Jinkela_wire_2789)
    );

    bfr new_Jinkela_buffer_3323 (
        .din(new_Jinkela_wire_3831),
        .dout(new_Jinkela_wire_3832)
    );

    bfr new_Jinkela_buffer_3304 (
        .din(new_Jinkela_wire_3812),
        .dout(new_Jinkela_wire_3813)
    );

    bfr new_Jinkela_buffer_2437 (
        .din(new_Jinkela_wire_2838),
        .dout(new_Jinkela_wire_2839)
    );

    bfr new_Jinkela_buffer_1596 (
        .din(new_Jinkela_wire_1939),
        .dout(new_Jinkela_wire_1940)
    );

    bfr new_Jinkela_buffer_2393 (
        .din(new_Jinkela_wire_2789),
        .dout(new_Jinkela_wire_2790)
    );

    bfr new_Jinkela_buffer_3305 (
        .din(new_Jinkela_wire_3813),
        .dout(new_Jinkela_wire_3814)
    );

    bfr new_Jinkela_buffer_6603 (
        .din(new_Jinkela_wire_8069),
        .dout(new_Jinkela_wire_8070)
    );

    bfr new_Jinkela_buffer_6636 (
        .din(new_Jinkela_wire_8121),
        .dout(new_Jinkela_wire_8122)
    );

    bfr new_Jinkela_buffer_6678 (
        .din(new_Jinkela_wire_8195),
        .dout(new_Jinkela_wire_8196)
    );

    bfr new_Jinkela_buffer_6637 (
        .din(new_Jinkela_wire_8122),
        .dout(new_Jinkela_wire_8123)
    );

    spl3L new_Jinkela_splitter_606 (
        .a(n_1009_),
        .d(new_Jinkela_wire_8270),
        .b(new_Jinkela_wire_8271),
        .c(new_Jinkela_wire_8272)
    );

    bfr new_Jinkela_buffer_6638 (
        .din(new_Jinkela_wire_8123),
        .dout(new_Jinkela_wire_8124)
    );

    spl2 new_Jinkela_splitter_603 (
        .a(new_Jinkela_wire_8196),
        .b(new_Jinkela_wire_8197),
        .c(new_Jinkela_wire_8198)
    );

    bfr new_Jinkela_buffer_6639 (
        .din(new_Jinkela_wire_8124),
        .dout(new_Jinkela_wire_8125)
    );

    bfr new_Jinkela_buffer_6743 (
        .din(new_Jinkela_wire_8268),
        .dout(new_Jinkela_wire_8269)
    );

    bfr new_Jinkela_buffer_6640 (
        .din(new_Jinkela_wire_8125),
        .dout(new_Jinkela_wire_8126)
    );

    spl2 new_Jinkela_splitter_608 (
        .a(n_0871_),
        .b(new_Jinkela_wire_8275),
        .c(new_Jinkela_wire_8276)
    );

    bfr new_Jinkela_buffer_6680 (
        .din(new_Jinkela_wire_8201),
        .dout(new_Jinkela_wire_8202)
    );

    bfr new_Jinkela_buffer_6641 (
        .din(new_Jinkela_wire_8126),
        .dout(new_Jinkela_wire_8127)
    );

    bfr new_Jinkela_buffer_6681 (
        .din(new_Jinkela_wire_8202),
        .dout(new_Jinkela_wire_8203)
    );

    bfr new_Jinkela_buffer_6642 (
        .din(new_Jinkela_wire_8127),
        .dout(new_Jinkela_wire_8128)
    );

    bfr new_Jinkela_buffer_6742 (
        .din(new_Jinkela_wire_8267),
        .dout(new_Jinkela_wire_8268)
    );

    bfr new_Jinkela_buffer_6643 (
        .din(new_Jinkela_wire_8128),
        .dout(new_Jinkela_wire_8129)
    );

    spl2 new_Jinkela_splitter_607 (
        .a(new_Jinkela_wire_8272),
        .b(new_Jinkela_wire_8273),
        .c(new_Jinkela_wire_8274)
    );

    bfr new_Jinkela_buffer_6682 (
        .din(new_Jinkela_wire_8203),
        .dout(new_Jinkela_wire_8204)
    );

    bfr new_Jinkela_buffer_6644 (
        .din(new_Jinkela_wire_8129),
        .dout(new_Jinkela_wire_8130)
    );

    and_bi n_2588_ (
        .a(new_Jinkela_wire_9551),
        .b(new_Jinkela_wire_9845),
        .c(n_0447_)
    );

    and_bi n_2587_ (
        .a(new_Jinkela_wire_9846),
        .b(new_Jinkela_wire_9552),
        .c(n_0446_)
    );

    bfr new_Jinkela_buffer_6645 (
        .din(new_Jinkela_wire_8130),
        .dout(new_Jinkela_wire_8131)
    );

    bfr new_Jinkela_buffer_6683 (
        .din(new_Jinkela_wire_8204),
        .dout(new_Jinkela_wire_8205)
    );

    bfr new_Jinkela_buffer_6646 (
        .din(new_Jinkela_wire_8131),
        .dout(new_Jinkela_wire_8132)
    );

    and_ii n_2586_ (
        .a(n_0444_),
        .b(n_0443_),
        .c(n_0445_)
    );

    bfr new_Jinkela_buffer_6647 (
        .din(new_Jinkela_wire_8132),
        .dout(new_Jinkela_wire_8133)
    );

    spl3L new_Jinkela_splitter_613 (
        .a(n_0990_),
        .d(new_Jinkela_wire_8285),
        .b(new_Jinkela_wire_8286),
        .c(new_Jinkela_wire_8287)
    );

    bfr new_Jinkela_buffer_6684 (
        .din(new_Jinkela_wire_8205),
        .dout(new_Jinkela_wire_8206)
    );

    bfr new_Jinkela_buffer_6648 (
        .din(new_Jinkela_wire_8133),
        .dout(new_Jinkela_wire_8134)
    );

    bfr new_Jinkela_buffer_6649 (
        .din(new_Jinkela_wire_8134),
        .dout(new_Jinkela_wire_8135)
    );

    spl2 new_Jinkela_splitter_609 (
        .a(n_0693_),
        .b(new_Jinkela_wire_8277),
        .c(new_Jinkela_wire_8278)
    );

    bfr new_Jinkela_buffer_6685 (
        .din(new_Jinkela_wire_8206),
        .dout(new_Jinkela_wire_8207)
    );

    bfr new_Jinkela_buffer_6650 (
        .din(new_Jinkela_wire_8135),
        .dout(new_Jinkela_wire_8136)
    );

    bfr new_Jinkela_buffer_6651 (
        .din(new_Jinkela_wire_8136),
        .dout(new_Jinkela_wire_8137)
    );

    bfr new_Jinkela_buffer_6686 (
        .din(new_Jinkela_wire_8207),
        .dout(new_Jinkela_wire_8208)
    );

    bfr new_Jinkela_buffer_6652 (
        .din(new_Jinkela_wire_8137),
        .dout(new_Jinkela_wire_8138)
    );

    spl2 new_Jinkela_splitter_610 (
        .a(n_0748_),
        .b(new_Jinkela_wire_8279),
        .c(new_Jinkela_wire_8280)
    );

    bfr new_Jinkela_buffer_6653 (
        .din(new_Jinkela_wire_8138),
        .dout(new_Jinkela_wire_8139)
    );

    spl2 new_Jinkela_splitter_611 (
        .a(n_0387_),
        .b(new_Jinkela_wire_8281),
        .c(new_Jinkela_wire_8282)
    );

    bfr new_Jinkela_buffer_6687 (
        .din(new_Jinkela_wire_8208),
        .dout(new_Jinkela_wire_8209)
    );

    bfr new_Jinkela_buffer_6654 (
        .din(new_Jinkela_wire_8139),
        .dout(new_Jinkela_wire_8140)
    );

    spl2 new_Jinkela_splitter_612 (
        .a(n_0083_),
        .b(new_Jinkela_wire_8283),
        .c(new_Jinkela_wire_8284)
    );

    bfr new_Jinkela_buffer_6655 (
        .din(new_Jinkela_wire_8140),
        .dout(new_Jinkela_wire_8141)
    );

    bfr new_Jinkela_buffer_7597 (
        .din(new_net_2566),
        .dout(new_Jinkela_wire_9519)
    );

    bfr new_Jinkela_buffer_49 (
        .din(new_Jinkela_wire_50),
        .dout(new_Jinkela_wire_51)
    );

    bfr new_Jinkela_buffer_103 (
        .din(new_Jinkela_wire_114),
        .dout(new_Jinkela_wire_115)
    );

    bfr new_Jinkela_buffer_50 (
        .din(new_Jinkela_wire_51),
        .dout(new_Jinkela_wire_52)
    );

    bfr new_Jinkela_buffer_51 (
        .din(new_Jinkela_wire_52),
        .dout(new_Jinkela_wire_53)
    );

    bfr new_Jinkela_buffer_104 (
        .din(new_Jinkela_wire_115),
        .dout(new_Jinkela_wire_116)
    );

    bfr new_Jinkela_buffer_52 (
        .din(new_Jinkela_wire_53),
        .dout(new_Jinkela_wire_54)
    );

    spl2 new_Jinkela_splitter_5 (
        .a(new_Jinkela_wire_179),
        .b(new_Jinkela_wire_180),
        .c(new_Jinkela_wire_181)
    );

    bfr new_Jinkela_buffer_53 (
        .din(new_Jinkela_wire_54),
        .dout(new_Jinkela_wire_55)
    );

    bfr new_Jinkela_buffer_105 (
        .din(new_Jinkela_wire_116),
        .dout(new_Jinkela_wire_117)
    );

    bfr new_Jinkela_buffer_54 (
        .din(new_Jinkela_wire_55),
        .dout(new_Jinkela_wire_56)
    );

    bfr new_Jinkela_buffer_55 (
        .din(new_Jinkela_wire_56),
        .dout(new_Jinkela_wire_57)
    );

    bfr new_Jinkela_buffer_106 (
        .din(new_Jinkela_wire_117),
        .dout(new_Jinkela_wire_118)
    );

    bfr new_Jinkela_buffer_56 (
        .din(new_Jinkela_wire_57),
        .dout(new_Jinkela_wire_58)
    );

    bfr new_Jinkela_buffer_173 (
        .din(new_Jinkela_wire_188),
        .dout(new_Jinkela_wire_189)
    );

    bfr new_Jinkela_buffer_57 (
        .din(new_Jinkela_wire_58),
        .dout(new_Jinkela_wire_59)
    );

    bfr new_Jinkela_buffer_107 (
        .din(new_Jinkela_wire_118),
        .dout(new_Jinkela_wire_119)
    );

    bfr new_Jinkela_buffer_58 (
        .din(new_Jinkela_wire_59),
        .dout(new_Jinkela_wire_60)
    );

    bfr new_Jinkela_buffer_170 (
        .din(new_Jinkela_wire_183),
        .dout(new_Jinkela_wire_184)
    );

    bfr new_Jinkela_buffer_59 (
        .din(new_Jinkela_wire_60),
        .dout(new_Jinkela_wire_61)
    );

    bfr new_Jinkela_buffer_108 (
        .din(new_Jinkela_wire_119),
        .dout(new_Jinkela_wire_120)
    );

    bfr new_Jinkela_buffer_60 (
        .din(new_Jinkela_wire_61),
        .dout(new_Jinkela_wire_62)
    );

    bfr new_Jinkela_buffer_171 (
        .din(new_Jinkela_wire_184),
        .dout(new_Jinkela_wire_185)
    );

    bfr new_Jinkela_buffer_61 (
        .din(new_Jinkela_wire_62),
        .dout(new_Jinkela_wire_63)
    );

    bfr new_Jinkela_buffer_109 (
        .din(new_Jinkela_wire_120),
        .dout(new_Jinkela_wire_121)
    );

    bfr new_Jinkela_buffer_62 (
        .din(new_Jinkela_wire_63),
        .dout(new_Jinkela_wire_64)
    );

    bfr new_Jinkela_buffer_176 (
        .din(N207),
        .dout(new_Jinkela_wire_192)
    );

    bfr new_Jinkela_buffer_63 (
        .din(new_Jinkela_wire_64),
        .dout(new_Jinkela_wire_65)
    );

    bfr new_Jinkela_buffer_110 (
        .din(new_Jinkela_wire_121),
        .dout(new_Jinkela_wire_122)
    );

    spl4L new_Jinkela_splitter_1 (
        .a(new_Jinkela_wire_65),
        .d(new_Jinkela_wire_66),
        .b(new_Jinkela_wire_67),
        .e(new_Jinkela_wire_68),
        .c(new_Jinkela_wire_69)
    );

    bfr new_Jinkela_buffer_111 (
        .din(new_Jinkela_wire_122),
        .dout(new_Jinkela_wire_123)
    );

    bfr new_Jinkela_buffer_180 (
        .din(N26),
        .dout(new_Jinkela_wire_196)
    );

    bfr new_Jinkela_buffer_174 (
        .din(new_Jinkela_wire_189),
        .dout(new_Jinkela_wire_190)
    );

    bfr new_Jinkela_buffer_112 (
        .din(new_Jinkela_wire_123),
        .dout(new_Jinkela_wire_124)
    );

    bfr new_Jinkela_buffer_177 (
        .din(new_Jinkela_wire_192),
        .dout(new_Jinkela_wire_193)
    );

    bfr new_Jinkela_buffer_113 (
        .din(new_Jinkela_wire_124),
        .dout(new_Jinkela_wire_125)
    );

    bfr new_Jinkela_buffer_175 (
        .din(new_Jinkela_wire_190),
        .dout(new_Jinkela_wire_191)
    );

    bfr new_Jinkela_buffer_114 (
        .din(new_Jinkela_wire_125),
        .dout(new_Jinkela_wire_126)
    );

    spl2 new_Jinkela_splitter_7 (
        .a(N346),
        .b(new_Jinkela_wire_200),
        .c(new_Jinkela_wire_201)
    );

    bfr new_Jinkela_buffer_248 (
        .din(N166),
        .dout(new_Jinkela_wire_268)
    );

    bfr new_Jinkela_buffer_115 (
        .din(new_Jinkela_wire_126),
        .dout(new_Jinkela_wire_127)
    );

    bfr new_Jinkela_buffer_178 (
        .din(new_Jinkela_wire_193),
        .dout(new_Jinkela_wire_194)
    );

    and_ii n_1863_ (
        .a(n_1128_),
        .b(n_1126_),
        .c(n_1129_)
    );

    and_ii n_2577_ (
        .a(new_Jinkela_wire_9749),
        .b(new_Jinkela_wire_8567),
        .c(n_0436_)
    );

    bfr new_Jinkela_buffer_5804 (
        .din(new_Jinkela_wire_6997),
        .dout(new_Jinkela_wire_6998)
    );

    and_ii n_1864_ (
        .a(new_Jinkela_wire_8869),
        .b(new_Jinkela_wire_6833),
        .c(n_1130_)
    );

    and_bi n_2578_ (
        .a(new_Jinkela_wire_6823),
        .b(new_Jinkela_wire_4443),
        .c(n_0437_)
    );

    bfr new_Jinkela_buffer_4143 (
        .din(new_Jinkela_wire_4843),
        .dout(new_Jinkela_wire_4844)
    );

    bfr new_Jinkela_buffer_5841 (
        .din(new_Jinkela_wire_7045),
        .dout(new_Jinkela_wire_7046)
    );

    and_bb n_1865_ (
        .a(new_Jinkela_wire_8868),
        .b(new_Jinkela_wire_6832),
        .c(n_1131_)
    );

    and_bi n_2579_ (
        .a(new_Jinkela_wire_9163),
        .b(new_Jinkela_wire_5594),
        .c(n_0438_)
    );

    spl3L new_Jinkela_splitter_275 (
        .a(n_0730_),
        .d(new_Jinkela_wire_4965),
        .b(new_Jinkela_wire_4966),
        .c(new_Jinkela_wire_4967)
    );

    bfr new_Jinkela_buffer_5805 (
        .din(new_Jinkela_wire_6998),
        .dout(new_Jinkela_wire_6999)
    );

    bfr new_Jinkela_buffer_4162 (
        .din(new_Jinkela_wire_4883),
        .dout(new_Jinkela_wire_4884)
    );

    or_bb n_1866_ (
        .a(n_1131_),
        .b(n_1130_),
        .c(n_1132_)
    );

    or_bb n_2580_ (
        .a(n_0438_),
        .b(n_0437_),
        .c(n_0439_)
    );

    bfr new_Jinkela_buffer_4144 (
        .din(new_Jinkela_wire_4844),
        .dout(new_Jinkela_wire_4845)
    );

    bfr new_Jinkela_buffer_5947 (
        .din(n_0311_),
        .dout(new_Jinkela_wire_7189)
    );

    and_bi n_1867_ (
        .a(new_Jinkela_wire_1237),
        .b(new_Jinkela_wire_3531),
        .c(n_1133_)
    );

    and_bi n_2581_ (
        .a(new_Jinkela_wire_6843),
        .b(new_Jinkela_wire_6794),
        .c(n_0440_)
    );

    bfr new_Jinkela_buffer_5806 (
        .din(new_Jinkela_wire_6999),
        .dout(new_Jinkela_wire_7000)
    );

    bfr new_Jinkela_buffer_4193 (
        .din(new_Jinkela_wire_4926),
        .dout(new_Jinkela_wire_4927)
    );

    and_ii n_1868_ (
        .a(new_Jinkela_wire_6887),
        .b(new_Jinkela_wire_9443),
        .c(n_1134_)
    );

    and_bi n_2582_ (
        .a(new_Jinkela_wire_6792),
        .b(new_Jinkela_wire_6844),
        .c(n_0441_)
    );

    bfr new_Jinkela_buffer_4145 (
        .din(new_Jinkela_wire_4845),
        .dout(new_Jinkela_wire_4846)
    );

    bfr new_Jinkela_buffer_5842 (
        .din(new_Jinkela_wire_7046),
        .dout(new_Jinkela_wire_7047)
    );

    and_bi n_1869_ (
        .a(new_Jinkela_wire_1242),
        .b(new_Jinkela_wire_775),
        .c(n_1135_)
    );

    or_bb n_2583_ (
        .a(n_0441_),
        .b(n_0440_),
        .c(n_0442_)
    );

    bfr new_Jinkela_buffer_5807 (
        .din(new_Jinkela_wire_7000),
        .dout(new_Jinkela_wire_7001)
    );

    bfr new_Jinkela_buffer_4163 (
        .din(new_Jinkela_wire_4884),
        .dout(new_Jinkela_wire_4885)
    );

    and_bb n_1870_ (
        .a(new_Jinkela_wire_5062),
        .b(new_Jinkela_wire_7746),
        .c(n_1136_)
    );

    and_ii n_2584_ (
        .a(new_Jinkela_wire_4533),
        .b(new_Jinkela_wire_7407),
        .c(n_0443_)
    );

    bfr new_Jinkela_buffer_4146 (
        .din(new_Jinkela_wire_4846),
        .dout(new_Jinkela_wire_4847)
    );

    bfr new_Jinkela_buffer_5868 (
        .din(new_Jinkela_wire_7100),
        .dout(new_Jinkela_wire_7101)
    );

    and_ii n_1871_ (
        .a(new_Jinkela_wire_5059),
        .b(new_Jinkela_wire_9464),
        .c(n_1137_)
    );

    and_bb n_2585_ (
        .a(new_Jinkela_wire_4532),
        .b(new_Jinkela_wire_7406),
        .c(n_0444_)
    );

    bfr new_Jinkela_buffer_5808 (
        .din(new_Jinkela_wire_7001),
        .dout(new_Jinkela_wire_7002)
    );

    and_bb n_1872_ (
        .a(new_Jinkela_wire_7844),
        .b(new_Jinkela_wire_6890),
        .c(n_1138_)
    );

    bfr new_Jinkela_buffer_4147 (
        .din(new_Jinkela_wire_4847),
        .dout(new_Jinkela_wire_4848)
    );

    bfr new_Jinkela_buffer_5843 (
        .din(new_Jinkela_wire_7047),
        .dout(new_Jinkela_wire_7048)
    );

    and_ii n_2590_ (
        .a(new_Jinkela_wire_8566),
        .b(new_Jinkela_wire_9579),
        .c(n_0449_)
    );

    and_ii n_1873_ (
        .a(n_1138_),
        .b(n_1136_),
        .c(n_1139_)
    );

    bfr new_Jinkela_buffer_5809 (
        .din(new_Jinkela_wire_7002),
        .dout(new_Jinkela_wire_7003)
    );

    and_bi n_2591_ (
        .a(new_Jinkela_wire_9158),
        .b(new_Jinkela_wire_4439),
        .c(n_0450_)
    );

    bfr new_Jinkela_buffer_4164 (
        .din(new_Jinkela_wire_4885),
        .dout(new_Jinkela_wire_4886)
    );

    or_bi n_1874_ (
        .a(new_Jinkela_wire_71),
        .b(new_Jinkela_wire_1701),
        .c(n_1140_)
    );

    bfr new_Jinkela_buffer_4148 (
        .din(new_Jinkela_wire_4848),
        .dout(new_Jinkela_wire_4849)
    );

    bfr new_Jinkela_buffer_5946 (
        .din(new_Jinkela_wire_7185),
        .dout(new_Jinkela_wire_7186)
    );

    and_ii n_2592_ (
        .a(new_Jinkela_wire_3778),
        .b(new_Jinkela_wire_6822),
        .c(n_0451_)
    );

    bfr new_Jinkela_buffer_5945 (
        .din(n_0577_),
        .dout(new_Jinkela_wire_7185)
    );

    and_bi n_1875_ (
        .a(new_Jinkela_wire_70),
        .b(new_Jinkela_wire_1700),
        .c(n_1141_)
    );

    bfr new_Jinkela_buffer_5810 (
        .din(new_Jinkela_wire_7003),
        .dout(new_Jinkela_wire_7004)
    );

    and_bi n_2593_ (
        .a(new_Jinkela_wire_7805),
        .b(new_Jinkela_wire_6798),
        .c(n_0452_)
    );

    bfr new_Jinkela_buffer_4194 (
        .din(new_Jinkela_wire_4927),
        .dout(new_Jinkela_wire_4928)
    );

    and_bi n_1876_ (
        .a(n_1140_),
        .b(n_1141_),
        .c(n_1142_)
    );

    bfr new_Jinkela_buffer_4149 (
        .din(new_Jinkela_wire_4849),
        .dout(new_Jinkela_wire_4850)
    );

    bfr new_Jinkela_buffer_5844 (
        .din(new_Jinkela_wire_7048),
        .dout(new_Jinkela_wire_7049)
    );

    and_bi n_2594_ (
        .a(new_Jinkela_wire_6797),
        .b(new_Jinkela_wire_7804),
        .c(n_0453_)
    );

    and_ii n_1877_ (
        .a(new_Jinkela_wire_4989),
        .b(new_Jinkela_wire_6262),
        .c(n_1143_)
    );

    bfr new_Jinkela_buffer_5811 (
        .din(new_Jinkela_wire_7004),
        .dout(new_Jinkela_wire_7005)
    );

    and_ii n_2595_ (
        .a(n_0453_),
        .b(n_0452_),
        .c(n_0454_)
    );

    bfr new_Jinkela_buffer_4165 (
        .din(new_Jinkela_wire_4886),
        .dout(new_Jinkela_wire_4887)
    );

    and_bi n_1878_ (
        .a(new_Jinkela_wire_9756),
        .b(new_Jinkela_wire_7823),
        .c(n_1144_)
    );

    bfr new_Jinkela_buffer_4150 (
        .din(new_Jinkela_wire_4850),
        .dout(new_Jinkela_wire_4851)
    );

    bfr new_Jinkela_buffer_5869 (
        .din(new_Jinkela_wire_7101),
        .dout(new_Jinkela_wire_7102)
    );

    and_ii n_2596_ (
        .a(new_Jinkela_wire_7503),
        .b(new_Jinkela_wire_5593),
        .c(n_0455_)
    );

    and_bi n_1879_ (
        .a(new_Jinkela_wire_7822),
        .b(new_Jinkela_wire_9755),
        .c(n_1145_)
    );

    bfr new_Jinkela_buffer_5812 (
        .din(new_Jinkela_wire_7005),
        .dout(new_Jinkela_wire_7006)
    );

    and_ii n_2597_ (
        .a(new_Jinkela_wire_9147),
        .b(new_Jinkela_wire_6604),
        .c(n_0456_)
    );

    bfr new_Jinkela_buffer_4224 (
        .din(n_0599_),
        .dout(new_Jinkela_wire_4970)
    );

    and_ii n_1880_ (
        .a(n_1145_),
        .b(n_1144_),
        .c(n_1146_)
    );

    spl2 new_Jinkela_splitter_259 (
        .a(new_Jinkela_wire_4851),
        .b(new_Jinkela_wire_4852),
        .c(new_Jinkela_wire_4853)
    );

    bfr new_Jinkela_buffer_5845 (
        .din(new_Jinkela_wire_7049),
        .dout(new_Jinkela_wire_7050)
    );

    or_ii n_2598_ (
        .a(new_Jinkela_wire_6060),
        .b(new_Jinkela_wire_6850),
        .c(n_0457_)
    );

    or_bb n_1881_ (
        .a(new_Jinkela_wire_8882),
        .b(new_Jinkela_wire_5096),
        .c(n_1147_)
    );

    bfr new_Jinkela_buffer_5813 (
        .din(new_Jinkela_wire_7006),
        .dout(new_Jinkela_wire_7007)
    );

    and_ii n_2599_ (
        .a(new_Jinkela_wire_6059),
        .b(new_Jinkela_wire_6849),
        .c(n_0458_)
    );

    bfr new_Jinkela_buffer_4195 (
        .din(new_Jinkela_wire_4928),
        .dout(new_Jinkela_wire_4929)
    );

    and_bb n_1882_ (
        .a(new_Jinkela_wire_8881),
        .b(new_Jinkela_wire_5095),
        .c(n_1148_)
    );

    and_bi n_2600_ (
        .a(n_0457_),
        .b(n_0458_),
        .c(n_0459_)
    );

    spl2 new_Jinkela_splitter_483 (
        .a(new_Jinkela_wire_7118),
        .b(new_Jinkela_wire_7119),
        .c(new_Jinkela_wire_7120)
    );

    bfr new_Jinkela_buffer_4166 (
        .din(new_Jinkela_wire_4887),
        .dout(new_Jinkela_wire_4888)
    );

    and_bi n_1883_ (
        .a(n_1147_),
        .b(n_1148_),
        .c(n_1149_)
    );

    bfr new_Jinkela_buffer_5814 (
        .din(new_Jinkela_wire_7007),
        .dout(new_Jinkela_wire_7008)
    );

    and_ii n_2601_ (
        .a(new_Jinkela_wire_7743),
        .b(new_Jinkela_wire_5419),
        .c(n_0460_)
    );

    bfr new_Jinkela_buffer_4167 (
        .din(new_Jinkela_wire_4888),
        .dout(new_Jinkela_wire_4889)
    );

    and_bb n_1884_ (
        .a(new_Jinkela_wire_1806),
        .b(new_Jinkela_wire_1362),
        .c(n_1150_)
    );

    bfr new_Jinkela_buffer_5846 (
        .din(new_Jinkela_wire_7050),
        .dout(new_Jinkela_wire_7051)
    );

    and_bb n_2602_ (
        .a(new_Jinkela_wire_7742),
        .b(new_Jinkela_wire_5418),
        .c(n_0461_)
    );

    spl2 new_Jinkela_splitter_276 (
        .a(n_0945_),
        .b(new_Jinkela_wire_4968),
        .c(new_Jinkela_wire_4969)
    );

    and_ii n_1885_ (
        .a(new_Jinkela_wire_7934),
        .b(new_Jinkela_wire_4984),
        .c(n_1151_)
    );

    bfr new_Jinkela_buffer_4223 (
        .din(new_Jinkela_wire_4959),
        .dout(new_Jinkela_wire_4960)
    );

    bfr new_Jinkela_buffer_5815 (
        .din(new_Jinkela_wire_7008),
        .dout(new_Jinkela_wire_7009)
    );

    and_ii n_2603_ (
        .a(n_0461_),
        .b(n_0460_),
        .c(n_0462_)
    );

    bfr new_Jinkela_buffer_4168 (
        .din(new_Jinkela_wire_4889),
        .dout(new_Jinkela_wire_4890)
    );

    and_bb n_1886_ (
        .a(new_Jinkela_wire_871),
        .b(new_Jinkela_wire_1300),
        .c(n_1152_)
    );

    bfr new_Jinkela_buffer_5870 (
        .din(new_Jinkela_wire_7102),
        .dout(new_Jinkela_wire_7103)
    );

    and_bi n_2604_ (
        .a(new_Jinkela_wire_5093),
        .b(new_Jinkela_wire_4077),
        .c(n_0463_)
    );

    bfr new_Jinkela_buffer_4196 (
        .din(new_Jinkela_wire_4929),
        .dout(new_Jinkela_wire_4930)
    );

    and_ii n_1887_ (
        .a(new_Jinkela_wire_8179),
        .b(new_Jinkela_wire_8327),
        .c(n_1153_)
    );

    bfr new_Jinkela_buffer_5816 (
        .din(new_Jinkela_wire_7009),
        .dout(new_Jinkela_wire_7010)
    );

    and_bi n_2605_ (
        .a(new_Jinkela_wire_4076),
        .b(new_Jinkela_wire_5092),
        .c(n_0464_)
    );

    bfr new_Jinkela_buffer_4169 (
        .din(new_Jinkela_wire_4890),
        .dout(new_Jinkela_wire_4891)
    );

    and_ii n_1888_ (
        .a(new_Jinkela_wire_3581),
        .b(new_Jinkela_wire_9005),
        .c(n_1154_)
    );

    bfr new_Jinkela_buffer_5847 (
        .din(new_Jinkela_wire_7051),
        .dout(new_Jinkela_wire_7052)
    );

    or_bb n_2606_ (
        .a(n_0464_),
        .b(n_0463_),
        .c(n_0465_)
    );

    spl2 new_Jinkela_splitter_273 (
        .a(new_Jinkela_wire_4960),
        .b(new_Jinkela_wire_4961),
        .c(new_Jinkela_wire_4962)
    );

    and_bb n_1889_ (
        .a(new_Jinkela_wire_3580),
        .b(new_Jinkela_wire_9006),
        .c(n_1155_)
    );

    and_bi n_2607_ (
        .a(new_Jinkela_wire_9574),
        .b(new_Jinkela_wire_9731),
        .c(n_0466_)
    );

    bfr new_Jinkela_buffer_5882 (
        .din(new_Jinkela_wire_7121),
        .dout(new_Jinkela_wire_7122)
    );

    bfr new_Jinkela_buffer_4170 (
        .din(new_Jinkela_wire_4891),
        .dout(new_Jinkela_wire_4892)
    );

    and_ii n_1890_ (
        .a(n_1155_),
        .b(n_1154_),
        .c(n_1156_)
    );

    bfr new_Jinkela_buffer_5848 (
        .din(new_Jinkela_wire_7052),
        .dout(new_Jinkela_wire_7053)
    );

    and_ii n_2608_ (
        .a(n_0466_),
        .b(n_0449_),
        .c(n_0467_)
    );

    bfr new_Jinkela_buffer_4197 (
        .din(new_Jinkela_wire_4930),
        .dout(new_Jinkela_wire_4931)
    );

    and_bb n_1891_ (
        .a(new_Jinkela_wire_2450),
        .b(new_Jinkela_wire_1260),
        .c(n_1157_)
    );

    bfr new_Jinkela_buffer_5871 (
        .din(new_Jinkela_wire_7103),
        .dout(new_Jinkela_wire_7104)
    );

    or_bi n_2609_ (
        .a(new_Jinkela_wire_4651),
        .b(new_Jinkela_wire_9960),
        .c(n_0468_)
    );

    bfr new_Jinkela_buffer_4171 (
        .din(new_Jinkela_wire_4892),
        .dout(new_Jinkela_wire_4893)
    );

    and_ii n_1892_ (
        .a(new_Jinkela_wire_5156),
        .b(new_Jinkela_wire_3836),
        .c(n_1158_)
    );

    bfr new_Jinkela_buffer_5849 (
        .din(new_Jinkela_wire_7053),
        .dout(new_Jinkela_wire_7054)
    );

    and_bi n_2610_ (
        .a(new_Jinkela_wire_4650),
        .b(new_Jinkela_wire_9959),
        .c(n_0469_)
    );

    spl4L new_Jinkela_splitter_277 (
        .a(n_1233_),
        .d(new_Jinkela_wire_4971),
        .b(new_Jinkela_wire_4972),
        .e(new_Jinkela_wire_4973),
        .c(new_Jinkela_wire_4974)
    );

    and_bb n_1893_ (
        .a(new_Jinkela_wire_682),
        .b(new_Jinkela_wire_1261),
        .c(n_1159_)
    );

    spl2 new_Jinkela_splitter_278 (
        .a(n_0893_),
        .b(new_Jinkela_wire_4975),
        .c(new_Jinkela_wire_4976)
    );

    and_bi n_2611_ (
        .a(n_0468_),
        .b(n_0469_),
        .c(new_net_2527)
    );

    bfr new_Jinkela_buffer_5883 (
        .din(new_Jinkela_wire_7122),
        .dout(new_Jinkela_wire_7123)
    );

    bfr new_Jinkela_buffer_4172 (
        .din(new_Jinkela_wire_4893),
        .dout(new_Jinkela_wire_4894)
    );

    and_ii n_1894_ (
        .a(new_Jinkela_wire_8443),
        .b(new_Jinkela_wire_8717),
        .c(n_1160_)
    );

    bfr new_Jinkela_buffer_5850 (
        .din(new_Jinkela_wire_7054),
        .dout(new_Jinkela_wire_7055)
    );

    and_bi n_2612_ (
        .a(new_Jinkela_wire_7018),
        .b(new_Jinkela_wire_4737),
        .c(n_0470_)
    );

    bfr new_Jinkela_buffer_4198 (
        .din(new_Jinkela_wire_4931),
        .dout(new_Jinkela_wire_4932)
    );

    and_bi n_1895_ (
        .a(new_Jinkela_wire_3724),
        .b(new_Jinkela_wire_4873),
        .c(n_1161_)
    );

    bfr new_Jinkela_buffer_5872 (
        .din(new_Jinkela_wire_7104),
        .dout(new_Jinkela_wire_7105)
    );

    or_bb n_2613_ (
        .a(n_0470_),
        .b(new_Jinkela_wire_8162),
        .c(n_0471_)
    );

    bfr new_Jinkela_buffer_4173 (
        .din(new_Jinkela_wire_4894),
        .dout(new_Jinkela_wire_4895)
    );

    and_bi n_1896_ (
        .a(new_Jinkela_wire_4871),
        .b(new_Jinkela_wire_3722),
        .c(n_1162_)
    );

    bfr new_Jinkela_buffer_5851 (
        .din(new_Jinkela_wire_7055),
        .dout(new_Jinkela_wire_7056)
    );

    and_bi n_2614_ (
        .a(new_Jinkela_wire_9040),
        .b(new_Jinkela_wire_9652),
        .c(n_0472_)
    );

    and_ii n_1897_ (
        .a(n_1162_),
        .b(n_1161_),
        .c(n_1163_)
    );

    and_bi n_2615_ (
        .a(new_Jinkela_wire_9650),
        .b(new_Jinkela_wire_9039),
        .c(n_0473_)
    );

    spl3L new_Jinkela_splitter_485 (
        .a(n_0930_),
        .d(new_Jinkela_wire_7200),
        .b(new_Jinkela_wire_7201),
        .c(new_Jinkela_wire_7202)
    );

    bfr new_Jinkela_buffer_4174 (
        .din(new_Jinkela_wire_4895),
        .dout(new_Jinkela_wire_4896)
    );

    and_bb n_1898_ (
        .a(new_Jinkela_wire_3558),
        .b(new_Jinkela_wire_1217),
        .c(n_1164_)
    );

    bfr new_Jinkela_buffer_5852 (
        .din(new_Jinkela_wire_7056),
        .dout(new_Jinkela_wire_7057)
    );

    and_ii n_2616_ (
        .a(n_0473_),
        .b(n_0472_),
        .c(n_0474_)
    );

    bfr new_Jinkela_buffer_4199 (
        .din(new_Jinkela_wire_4932),
        .dout(new_Jinkela_wire_4933)
    );

    and_ii n_1899_ (
        .a(new_Jinkela_wire_5978),
        .b(new_Jinkela_wire_4521),
        .c(n_1165_)
    );

    bfr new_Jinkela_buffer_5873 (
        .din(new_Jinkela_wire_7105),
        .dout(new_Jinkela_wire_7106)
    );

    and_bi n_2617_ (
        .a(new_Jinkela_wire_8020),
        .b(new_Jinkela_wire_6309),
        .c(n_0475_)
    );

    bfr new_Jinkela_buffer_4175 (
        .din(new_Jinkela_wire_4896),
        .dout(new_Jinkela_wire_4897)
    );

    and_bb n_1900_ (
        .a(new_Jinkela_wire_2474),
        .b(new_Jinkela_wire_1331),
        .c(n_1166_)
    );

    bfr new_Jinkela_buffer_5853 (
        .din(new_Jinkela_wire_7057),
        .dout(new_Jinkela_wire_7058)
    );

    and_bi n_2618_ (
        .a(new_Jinkela_wire_6308),
        .b(new_Jinkela_wire_8021),
        .c(n_0476_)
    );

    and_ii n_1901_ (
        .a(new_Jinkela_wire_9649),
        .b(new_Jinkela_wire_7927),
        .c(n_1167_)
    );

    or_bb n_2619_ (
        .a(n_0476_),
        .b(n_0475_),
        .c(n_0477_)
    );

    bfr new_Jinkela_buffer_5884 (
        .din(new_Jinkela_wire_7123),
        .dout(new_Jinkela_wire_7124)
    );

    bfr new_Jinkela_buffer_4176 (
        .din(new_Jinkela_wire_4897),
        .dout(new_Jinkela_wire_4898)
    );

    and_ii n_1902_ (
        .a(new_Jinkela_wire_5366),
        .b(new_Jinkela_wire_10525),
        .c(n_1168_)
    );

    bfr new_Jinkela_buffer_5854 (
        .din(new_Jinkela_wire_7058),
        .dout(new_Jinkela_wire_7059)
    );

    and_ii n_2620_ (
        .a(new_Jinkela_wire_5755),
        .b(new_Jinkela_wire_9200),
        .c(n_0478_)
    );

    bfr new_Jinkela_buffer_4200 (
        .din(new_Jinkela_wire_4933),
        .dout(new_Jinkela_wire_4934)
    );

    and_bb n_1903_ (
        .a(new_Jinkela_wire_5364),
        .b(new_Jinkela_wire_10524),
        .c(n_1169_)
    );

    bfr new_Jinkela_buffer_5874 (
        .din(new_Jinkela_wire_7106),
        .dout(new_Jinkela_wire_7107)
    );

    and_bi n_2621_ (
        .a(new_Jinkela_wire_7024),
        .b(new_Jinkela_wire_3835),
        .c(n_0479_)
    );

    bfr new_Jinkela_buffer_4177 (
        .din(new_Jinkela_wire_4898),
        .dout(new_Jinkela_wire_4899)
    );

    and_ii n_1904_ (
        .a(n_1169_),
        .b(n_1168_),
        .c(n_1170_)
    );

    bfr new_Jinkela_buffer_5855 (
        .din(new_Jinkela_wire_7059),
        .dout(new_Jinkela_wire_7060)
    );

    bfr new_Jinkela_buffer_2502 (
        .din(new_Jinkela_wire_2903),
        .dout(new_Jinkela_wire_2904)
    );

    bfr new_Jinkela_buffer_2394 (
        .din(new_Jinkela_wire_2790),
        .dout(new_Jinkela_wire_2791)
    );

    bfr new_Jinkela_buffer_2438 (
        .din(new_Jinkela_wire_2839),
        .dout(new_Jinkela_wire_2840)
    );

    bfr new_Jinkela_buffer_2395 (
        .din(new_Jinkela_wire_2791),
        .dout(new_Jinkela_wire_2792)
    );

    bfr new_Jinkela_buffer_2567 (
        .din(new_Jinkela_wire_2968),
        .dout(new_Jinkela_wire_2969)
    );

    bfr new_Jinkela_buffer_2396 (
        .din(new_Jinkela_wire_2792),
        .dout(new_Jinkela_wire_2793)
    );

    bfr new_Jinkela_buffer_2439 (
        .din(new_Jinkela_wire_2840),
        .dout(new_Jinkela_wire_2841)
    );

    bfr new_Jinkela_buffer_2397 (
        .din(new_Jinkela_wire_2793),
        .dout(new_Jinkela_wire_2794)
    );

    bfr new_Jinkela_buffer_2503 (
        .din(new_Jinkela_wire_2904),
        .dout(new_Jinkela_wire_2905)
    );

    bfr new_Jinkela_buffer_2398 (
        .din(new_Jinkela_wire_2794),
        .dout(new_Jinkela_wire_2795)
    );

    bfr new_Jinkela_buffer_2440 (
        .din(new_Jinkela_wire_2841),
        .dout(new_Jinkela_wire_2842)
    );

    bfr new_Jinkela_buffer_2399 (
        .din(new_Jinkela_wire_2795),
        .dout(new_Jinkela_wire_2796)
    );

    spl4L new_Jinkela_splitter_135 (
        .a(N267),
        .d(new_Jinkela_wire_2976),
        .b(new_Jinkela_wire_2977),
        .e(new_Jinkela_wire_2978),
        .c(new_Jinkela_wire_2979)
    );

    bfr new_Jinkela_buffer_2639 (
        .din(N204),
        .dout(new_Jinkela_wire_3045)
    );

    bfr new_Jinkela_buffer_2400 (
        .din(new_Jinkela_wire_2796),
        .dout(new_Jinkela_wire_2797)
    );

    bfr new_Jinkela_buffer_2441 (
        .din(new_Jinkela_wire_2842),
        .dout(new_Jinkela_wire_2843)
    );

    bfr new_Jinkela_buffer_2401 (
        .din(new_Jinkela_wire_2797),
        .dout(new_Jinkela_wire_2798)
    );

    bfr new_Jinkela_buffer_2504 (
        .din(new_Jinkela_wire_2905),
        .dout(new_Jinkela_wire_2906)
    );

    bfr new_Jinkela_buffer_2402 (
        .din(new_Jinkela_wire_2798),
        .dout(new_Jinkela_wire_2799)
    );

    bfr new_Jinkela_buffer_2442 (
        .din(new_Jinkela_wire_2843),
        .dout(new_Jinkela_wire_2844)
    );

    bfr new_Jinkela_buffer_2403 (
        .din(new_Jinkela_wire_2799),
        .dout(new_Jinkela_wire_2800)
    );

    bfr new_Jinkela_buffer_2568 (
        .din(new_Jinkela_wire_2969),
        .dout(new_Jinkela_wire_2970)
    );

    bfr new_Jinkela_buffer_2404 (
        .din(new_Jinkela_wire_2800),
        .dout(new_Jinkela_wire_2801)
    );

    bfr new_Jinkela_buffer_2443 (
        .din(new_Jinkela_wire_2844),
        .dout(new_Jinkela_wire_2845)
    );

    bfr new_Jinkela_buffer_2405 (
        .din(new_Jinkela_wire_2801),
        .dout(new_Jinkela_wire_2802)
    );

    bfr new_Jinkela_buffer_2505 (
        .din(new_Jinkela_wire_2906),
        .dout(new_Jinkela_wire_2907)
    );

    bfr new_Jinkela_buffer_2406 (
        .din(new_Jinkela_wire_2802),
        .dout(new_Jinkela_wire_2803)
    );

    bfr new_Jinkela_buffer_2444 (
        .din(new_Jinkela_wire_2845),
        .dout(new_Jinkela_wire_2846)
    );

    bfr new_Jinkela_buffer_2407 (
        .din(new_Jinkela_wire_2803),
        .dout(new_Jinkela_wire_2804)
    );

    bfr new_Jinkela_buffer_2571 (
        .din(new_Jinkela_wire_2972),
        .dout(new_Jinkela_wire_2973)
    );

    bfr new_Jinkela_buffer_2445 (
        .din(new_Jinkela_wire_2846),
        .dout(new_Jinkela_wire_2847)
    );

    bfr new_Jinkela_buffer_2506 (
        .din(new_Jinkela_wire_2907),
        .dout(new_Jinkela_wire_2908)
    );

    bfr new_Jinkela_buffer_2446 (
        .din(new_Jinkela_wire_2847),
        .dout(new_Jinkela_wire_2848)
    );

    bfr new_Jinkela_buffer_2569 (
        .din(new_Jinkela_wire_2970),
        .dout(new_Jinkela_wire_2971)
    );

    bfr new_Jinkela_buffer_2447 (
        .din(new_Jinkela_wire_2848),
        .dout(new_Jinkela_wire_2849)
    );

    bfr new_Jinkela_buffer_2507 (
        .din(new_Jinkela_wire_2908),
        .dout(new_Jinkela_wire_2909)
    );

    bfr new_Jinkela_buffer_2448 (
        .din(new_Jinkela_wire_2849),
        .dout(new_Jinkela_wire_2850)
    );

    bfr new_Jinkela_buffer_2574 (
        .din(new_Jinkela_wire_2979),
        .dout(new_Jinkela_wire_2980)
    );

    bfr new_Jinkela_buffer_2449 (
        .din(new_Jinkela_wire_2850),
        .dout(new_Jinkela_wire_2851)
    );

    bfr new_Jinkela_buffer_2508 (
        .din(new_Jinkela_wire_2909),
        .dout(new_Jinkela_wire_2910)
    );

    bfr new_Jinkela_buffer_2450 (
        .din(new_Jinkela_wire_2851),
        .dout(new_Jinkela_wire_2852)
    );

    bfr new_Jinkela_buffer_2572 (
        .din(new_Jinkela_wire_2973),
        .dout(new_Jinkela_wire_2974)
    );

    bfr new_Jinkela_buffer_2451 (
        .din(new_Jinkela_wire_2852),
        .dout(new_Jinkela_wire_2853)
    );

    bfr new_Jinkela_buffer_1721 (
        .din(new_Jinkela_wire_2066),
        .dout(new_Jinkela_wire_2067)
    );

    bfr new_Jinkela_buffer_3324 (
        .din(new_Jinkela_wire_3832),
        .dout(new_Jinkela_wire_3833)
    );

    bfr new_Jinkela_buffer_1597 (
        .din(new_Jinkela_wire_1940),
        .dout(new_Jinkela_wire_1941)
    );

    bfr new_Jinkela_buffer_3306 (
        .din(new_Jinkela_wire_3814),
        .dout(new_Jinkela_wire_3815)
    );

    bfr new_Jinkela_buffer_1724 (
        .din(new_Jinkela_wire_2069),
        .dout(new_Jinkela_wire_2070)
    );

    bfr new_Jinkela_buffer_1658 (
        .din(new_Jinkela_wire_2003),
        .dout(new_Jinkela_wire_2004)
    );

    bfr new_Jinkela_buffer_3331 (
        .din(new_Jinkela_wire_3845),
        .dout(new_Jinkela_wire_3846)
    );

    bfr new_Jinkela_buffer_1598 (
        .din(new_Jinkela_wire_1941),
        .dout(new_Jinkela_wire_1942)
    );

    bfr new_Jinkela_buffer_3307 (
        .din(new_Jinkela_wire_3815),
        .dout(new_Jinkela_wire_3816)
    );

    bfr new_Jinkela_buffer_3325 (
        .din(new_Jinkela_wire_3833),
        .dout(new_Jinkela_wire_3834)
    );

    bfr new_Jinkela_buffer_1599 (
        .din(new_Jinkela_wire_1942),
        .dout(new_Jinkela_wire_1943)
    );

    bfr new_Jinkela_buffer_3308 (
        .din(new_Jinkela_wire_3816),
        .dout(new_Jinkela_wire_3817)
    );

    bfr new_Jinkela_buffer_1722 (
        .din(new_Jinkela_wire_2067),
        .dout(new_Jinkela_wire_2068)
    );

    bfr new_Jinkela_buffer_1659 (
        .din(new_Jinkela_wire_2004),
        .dout(new_Jinkela_wire_2005)
    );

    bfr new_Jinkela_buffer_1600 (
        .din(new_Jinkela_wire_1943),
        .dout(new_Jinkela_wire_1944)
    );

    bfr new_Jinkela_buffer_3309 (
        .din(new_Jinkela_wire_3817),
        .dout(new_Jinkela_wire_3818)
    );

    bfr new_Jinkela_buffer_3336 (
        .din(n_0818_),
        .dout(new_Jinkela_wire_3855)
    );

    bfr new_Jinkela_buffer_3332 (
        .din(new_Jinkela_wire_3846),
        .dout(new_Jinkela_wire_3847)
    );

    bfr new_Jinkela_buffer_1601 (
        .din(new_Jinkela_wire_1944),
        .dout(new_Jinkela_wire_1945)
    );

    bfr new_Jinkela_buffer_3310 (
        .din(new_Jinkela_wire_3818),
        .dout(new_Jinkela_wire_3819)
    );

    bfr new_Jinkela_buffer_1731 (
        .din(N201),
        .dout(new_Jinkela_wire_2077)
    );

    bfr new_Jinkela_buffer_1660 (
        .din(new_Jinkela_wire_2005),
        .dout(new_Jinkela_wire_2006)
    );

    bfr new_Jinkela_buffer_1602 (
        .din(new_Jinkela_wire_1945),
        .dout(new_Jinkela_wire_1946)
    );

    bfr new_Jinkela_buffer_3311 (
        .din(new_Jinkela_wire_3819),
        .dout(new_Jinkela_wire_3820)
    );

    bfr new_Jinkela_buffer_3333 (
        .din(new_Jinkela_wire_3847),
        .dout(new_Jinkela_wire_3848)
    );

    bfr new_Jinkela_buffer_1603 (
        .din(new_Jinkela_wire_1946),
        .dout(new_Jinkela_wire_1947)
    );

    bfr new_Jinkela_buffer_3312 (
        .din(new_Jinkela_wire_3820),
        .dout(new_Jinkela_wire_3821)
    );

    bfr new_Jinkela_buffer_1725 (
        .din(new_Jinkela_wire_2070),
        .dout(new_Jinkela_wire_2071)
    );

    bfr new_Jinkela_buffer_1661 (
        .din(new_Jinkela_wire_2006),
        .dout(new_Jinkela_wire_2007)
    );

    spl2 new_Jinkela_splitter_183 (
        .a(n_1199_),
        .b(new_Jinkela_wire_3860),
        .c(new_Jinkela_wire_3861)
    );

    bfr new_Jinkela_buffer_1604 (
        .din(new_Jinkela_wire_1947),
        .dout(new_Jinkela_wire_1948)
    );

    bfr new_Jinkela_buffer_3337 (
        .din(new_Jinkela_wire_3855),
        .dout(new_Jinkela_wire_3856)
    );

    bfr new_Jinkela_buffer_3334 (
        .din(new_Jinkela_wire_3848),
        .dout(new_Jinkela_wire_3849)
    );

    bfr new_Jinkela_buffer_1605 (
        .din(new_Jinkela_wire_1948),
        .dout(new_Jinkela_wire_1949)
    );

    bfr new_Jinkela_buffer_3335 (
        .din(new_Jinkela_wire_3849),
        .dout(new_Jinkela_wire_3850)
    );

    bfr new_Jinkela_buffer_1728 (
        .din(new_Jinkela_wire_2073),
        .dout(new_Jinkela_wire_2074)
    );

    bfr new_Jinkela_buffer_1662 (
        .din(new_Jinkela_wire_2007),
        .dout(new_Jinkela_wire_2008)
    );

    spl4L new_Jinkela_splitter_184 (
        .a(n_0761_),
        .d(new_Jinkela_wire_3862),
        .b(new_Jinkela_wire_3863),
        .e(new_Jinkela_wire_3864),
        .c(new_Jinkela_wire_3865)
    );

    bfr new_Jinkela_buffer_1606 (
        .din(new_Jinkela_wire_1949),
        .dout(new_Jinkela_wire_1950)
    );

    bfr new_Jinkela_buffer_3338 (
        .din(new_Jinkela_wire_3856),
        .dout(new_Jinkela_wire_3857)
    );

    spl4L new_Jinkela_splitter_185 (
        .a(n_1262_),
        .d(new_Jinkela_wire_3866),
        .b(new_Jinkela_wire_3867),
        .e(new_Jinkela_wire_3868),
        .c(new_Jinkela_wire_3869)
    );

    bfr new_Jinkela_buffer_1607 (
        .din(new_Jinkela_wire_1950),
        .dout(new_Jinkela_wire_1951)
    );

    spl2 new_Jinkela_splitter_182 (
        .a(new_Jinkela_wire_3857),
        .b(new_Jinkela_wire_3858),
        .c(new_Jinkela_wire_3859)
    );

    bfr new_Jinkela_buffer_1726 (
        .din(new_Jinkela_wire_2071),
        .dout(new_Jinkela_wire_2072)
    );

    bfr new_Jinkela_buffer_1663 (
        .din(new_Jinkela_wire_2008),
        .dout(new_Jinkela_wire_2009)
    );

    spl2 new_Jinkela_splitter_186 (
        .a(n_0119_),
        .b(new_Jinkela_wire_3870),
        .c(new_Jinkela_wire_3871)
    );

    bfr new_Jinkela_buffer_1608 (
        .din(new_Jinkela_wire_1951),
        .dout(new_Jinkela_wire_1952)
    );

    bfr new_Jinkela_buffer_3340 (
        .din(n_1303_),
        .dout(new_Jinkela_wire_3873)
    );

    bfr new_Jinkela_buffer_3339 (
        .din(new_Jinkela_wire_3871),
        .dout(new_Jinkela_wire_3872)
    );

    bfr new_Jinkela_buffer_1609 (
        .din(new_Jinkela_wire_1952),
        .dout(new_Jinkela_wire_1953)
    );

    bfr new_Jinkela_buffer_3343 (
        .din(new_net_2535),
        .dout(new_Jinkela_wire_3878)
    );

    spl3L new_Jinkela_splitter_188 (
        .a(n_0587_),
        .d(new_Jinkela_wire_3911),
        .b(new_Jinkela_wire_3912),
        .c(new_Jinkela_wire_3913)
    );

    bfr new_Jinkela_buffer_1735 (
        .din(N286),
        .dout(new_Jinkela_wire_2081)
    );

    bfr new_Jinkela_buffer_1664 (
        .din(new_Jinkela_wire_2009),
        .dout(new_Jinkela_wire_2010)
    );

    bfr new_Jinkela_buffer_3341 (
        .din(new_Jinkela_wire_3873),
        .dout(new_Jinkela_wire_3874)
    );

    spl2 new_Jinkela_splitter_190 (
        .a(n_0663_),
        .b(new_Jinkela_wire_3921),
        .c(new_Jinkela_wire_3922)
    );

    bfr new_Jinkela_buffer_1610 (
        .din(new_Jinkela_wire_1953),
        .dout(new_Jinkela_wire_1954)
    );

    bfr new_Jinkela_buffer_3344 (
        .din(new_Jinkela_wire_3878),
        .dout(new_Jinkela_wire_3879)
    );

    bfr new_Jinkela_buffer_1799 (
        .din(N170),
        .dout(new_Jinkela_wire_2150)
    );

    spl2 new_Jinkela_splitter_187 (
        .a(new_Jinkela_wire_3874),
        .b(new_Jinkela_wire_3875),
        .c(new_Jinkela_wire_3876)
    );

    bfr new_Jinkela_buffer_1611 (
        .din(new_Jinkela_wire_1954),
        .dout(new_Jinkela_wire_1955)
    );

    bfr new_Jinkela_buffer_3342 (
        .din(new_Jinkela_wire_3876),
        .dout(new_Jinkela_wire_3877)
    );

    bfr new_Jinkela_buffer_1729 (
        .din(new_Jinkela_wire_2074),
        .dout(new_Jinkela_wire_2075)
    );

    bfr new_Jinkela_buffer_1665 (
        .din(new_Jinkela_wire_2010),
        .dout(new_Jinkela_wire_2011)
    );

    bfr new_Jinkela_buffer_1612 (
        .din(new_Jinkela_wire_1955),
        .dout(new_Jinkela_wire_1956)
    );

    bfr new_Jinkela_buffer_3345 (
        .din(new_Jinkela_wire_3879),
        .dout(new_Jinkela_wire_3880)
    );

    bfr new_Jinkela_buffer_1613 (
        .din(new_Jinkela_wire_1956),
        .dout(new_Jinkela_wire_1957)
    );

    bfr new_Jinkela_buffer_3381 (
        .din(new_Jinkela_wire_3922),
        .dout(new_Jinkela_wire_3923)
    );

    bfr new_Jinkela_buffer_3346 (
        .din(new_Jinkela_wire_3880),
        .dout(new_Jinkela_wire_3881)
    );

    bfr new_Jinkela_buffer_1732 (
        .din(new_Jinkela_wire_2077),
        .dout(new_Jinkela_wire_2078)
    );

    bfr new_Jinkela_buffer_1666 (
        .din(new_Jinkela_wire_2011),
        .dout(new_Jinkela_wire_2012)
    );

    bfr new_Jinkela_buffer_3376 (
        .din(new_Jinkela_wire_3913),
        .dout(new_Jinkela_wire_3914)
    );

    bfr new_Jinkela_buffer_1614 (
        .din(new_Jinkela_wire_1957),
        .dout(new_Jinkela_wire_1958)
    );

    bfr new_Jinkela_buffer_3347 (
        .din(new_Jinkela_wire_3881),
        .dout(new_Jinkela_wire_3882)
    );

    spl2 new_Jinkela_splitter_193 (
        .a(n_0951_),
        .b(new_Jinkela_wire_3934),
        .c(new_Jinkela_wire_3935)
    );

    bfr new_Jinkela_buffer_1615 (
        .din(new_Jinkela_wire_1958),
        .dout(new_Jinkela_wire_1959)
    );

    bfr new_Jinkela_buffer_3384 (
        .din(n_0767_),
        .dout(new_Jinkela_wire_3929)
    );

    bfr new_Jinkela_buffer_3348 (
        .din(new_Jinkela_wire_3882),
        .dout(new_Jinkela_wire_3883)
    );

    bfr new_Jinkela_buffer_1730 (
        .din(new_Jinkela_wire_2075),
        .dout(new_Jinkela_wire_2076)
    );

    bfr new_Jinkela_buffer_1667 (
        .din(new_Jinkela_wire_2012),
        .dout(new_Jinkela_wire_2013)
    );

    bfr new_Jinkela_buffer_3377 (
        .din(new_Jinkela_wire_3914),
        .dout(new_Jinkela_wire_3915)
    );

    bfr new_Jinkela_buffer_1616 (
        .din(new_Jinkela_wire_1959),
        .dout(new_Jinkela_wire_1960)
    );

    bfr new_Jinkela_buffer_3349 (
        .din(new_Jinkela_wire_3883),
        .dout(new_Jinkela_wire_3884)
    );

    bfr new_Jinkela_buffer_1617 (
        .din(new_Jinkela_wire_1960),
        .dout(new_Jinkela_wire_1961)
    );

    bfr new_Jinkela_buffer_5002 (
        .din(new_Jinkela_wire_5959),
        .dout(new_Jinkela_wire_5960)
    );

    bfr new_Jinkela_buffer_5043 (
        .din(new_Jinkela_wire_6018),
        .dout(new_Jinkela_wire_6019)
    );

    bfr new_Jinkela_buffer_5003 (
        .din(new_Jinkela_wire_5960),
        .dout(new_Jinkela_wire_5961)
    );

    bfr new_Jinkela_buffer_5025 (
        .din(new_Jinkela_wire_5989),
        .dout(new_Jinkela_wire_5990)
    );

    bfr new_Jinkela_buffer_5004 (
        .din(new_Jinkela_wire_5961),
        .dout(new_Jinkela_wire_5962)
    );

    spl2 new_Jinkela_splitter_376 (
        .a(n_0392_),
        .b(new_Jinkela_wire_6097),
        .c(new_Jinkela_wire_6098)
    );

    bfr new_Jinkela_buffer_5005 (
        .din(new_Jinkela_wire_5962),
        .dout(new_Jinkela_wire_5963)
    );

    bfr new_Jinkela_buffer_5084 (
        .din(new_Jinkela_wire_6061),
        .dout(new_Jinkela_wire_6062)
    );

    bfr new_Jinkela_buffer_5026 (
        .din(new_Jinkela_wire_5990),
        .dout(new_Jinkela_wire_5991)
    );

    bfr new_Jinkela_buffer_5006 (
        .din(new_Jinkela_wire_5963),
        .dout(new_Jinkela_wire_5964)
    );

    bfr new_Jinkela_buffer_5044 (
        .din(new_Jinkela_wire_6019),
        .dout(new_Jinkela_wire_6020)
    );

    bfr new_Jinkela_buffer_5007 (
        .din(new_Jinkela_wire_5964),
        .dout(new_Jinkela_wire_5965)
    );

    bfr new_Jinkela_buffer_5027 (
        .din(new_Jinkela_wire_5991),
        .dout(new_Jinkela_wire_5992)
    );

    bfr new_Jinkela_buffer_5008 (
        .din(new_Jinkela_wire_5965),
        .dout(new_Jinkela_wire_5966)
    );

    bfr new_Jinkela_buffer_5009 (
        .din(new_Jinkela_wire_5966),
        .dout(new_Jinkela_wire_5967)
    );

    bfr new_Jinkela_buffer_5109 (
        .din(new_Jinkela_wire_6088),
        .dout(new_Jinkela_wire_6089)
    );

    bfr new_Jinkela_buffer_5028 (
        .din(new_Jinkela_wire_5992),
        .dout(new_Jinkela_wire_5993)
    );

    spl2 new_Jinkela_splitter_366 (
        .a(new_Jinkela_wire_5967),
        .b(new_Jinkela_wire_5968),
        .c(new_Jinkela_wire_5969)
    );

    bfr new_Jinkela_buffer_5029 (
        .din(new_Jinkela_wire_5993),
        .dout(new_Jinkela_wire_5994)
    );

    bfr new_Jinkela_buffer_5045 (
        .din(new_Jinkela_wire_6020),
        .dout(new_Jinkela_wire_6021)
    );

    bfr new_Jinkela_buffer_5085 (
        .din(new_Jinkela_wire_6062),
        .dout(new_Jinkela_wire_6063)
    );

    bfr new_Jinkela_buffer_5030 (
        .din(new_Jinkela_wire_5994),
        .dout(new_Jinkela_wire_5995)
    );

    bfr new_Jinkela_buffer_5046 (
        .din(new_Jinkela_wire_6021),
        .dout(new_Jinkela_wire_6022)
    );

    bfr new_Jinkela_buffer_5031 (
        .din(new_Jinkela_wire_5995),
        .dout(new_Jinkela_wire_5996)
    );

    bfr new_Jinkela_buffer_5032 (
        .din(new_Jinkela_wire_5996),
        .dout(new_Jinkela_wire_5997)
    );

    bfr new_Jinkela_buffer_5047 (
        .din(new_Jinkela_wire_6022),
        .dout(new_Jinkela_wire_6023)
    );

    bfr new_Jinkela_buffer_5033 (
        .din(new_Jinkela_wire_5997),
        .dout(new_Jinkela_wire_5998)
    );

    bfr new_Jinkela_buffer_5086 (
        .din(new_Jinkela_wire_6063),
        .dout(new_Jinkela_wire_6064)
    );

    bfr new_Jinkela_buffer_5034 (
        .din(new_Jinkela_wire_5998),
        .dout(new_Jinkela_wire_5999)
    );

    bfr new_Jinkela_buffer_5048 (
        .din(new_Jinkela_wire_6023),
        .dout(new_Jinkela_wire_6024)
    );

    bfr new_Jinkela_buffer_5035 (
        .din(new_Jinkela_wire_5999),
        .dout(new_Jinkela_wire_6000)
    );

    spl3L new_Jinkela_splitter_377 (
        .a(n_0666_),
        .d(new_Jinkela_wire_6099),
        .b(new_Jinkela_wire_6100),
        .c(new_Jinkela_wire_6101)
    );

    bfr new_Jinkela_buffer_5036 (
        .din(new_Jinkela_wire_6000),
        .dout(new_Jinkela_wire_6001)
    );

    bfr new_Jinkela_buffer_5049 (
        .din(new_Jinkela_wire_6024),
        .dout(new_Jinkela_wire_6025)
    );

    bfr new_Jinkela_buffer_5037 (
        .din(new_Jinkela_wire_6001),
        .dout(new_Jinkela_wire_6002)
    );

    bfr new_Jinkela_buffer_5087 (
        .din(new_Jinkela_wire_6064),
        .dout(new_Jinkela_wire_6065)
    );

    bfr new_Jinkela_buffer_5038 (
        .din(new_Jinkela_wire_6002),
        .dout(new_Jinkela_wire_6003)
    );

    bfr new_Jinkela_buffer_5050 (
        .din(new_Jinkela_wire_6025),
        .dout(new_Jinkela_wire_6026)
    );

    bfr new_Jinkela_buffer_5039 (
        .din(new_Jinkela_wire_6003),
        .dout(new_Jinkela_wire_6004)
    );

    spl3L new_Jinkela_splitter_379 (
        .a(n_1228_),
        .d(new_Jinkela_wire_6105),
        .b(new_Jinkela_wire_6106),
        .c(new_Jinkela_wire_6107)
    );

    bfr new_Jinkela_buffer_5040 (
        .din(new_Jinkela_wire_6004),
        .dout(new_Jinkela_wire_6005)
    );

    bfr new_Jinkela_buffer_5051 (
        .din(new_Jinkela_wire_6026),
        .dout(new_Jinkela_wire_6027)
    );

    bfr new_Jinkela_buffer_6688 (
        .din(new_Jinkela_wire_8209),
        .dout(new_Jinkela_wire_8210)
    );

    bfr new_Jinkela_buffer_6656 (
        .din(new_Jinkela_wire_8141),
        .dout(new_Jinkela_wire_8142)
    );

    bfr new_Jinkela_buffer_6657 (
        .din(new_Jinkela_wire_8142),
        .dout(new_Jinkela_wire_8143)
    );

    bfr new_Jinkela_buffer_6689 (
        .din(new_Jinkela_wire_8210),
        .dout(new_Jinkela_wire_8211)
    );

    bfr new_Jinkela_buffer_6658 (
        .din(new_Jinkela_wire_8143),
        .dout(new_Jinkela_wire_8144)
    );

    spl4L new_Jinkela_splitter_615 (
        .a(n_1273_),
        .d(new_Jinkela_wire_8290),
        .b(new_Jinkela_wire_8291),
        .e(new_Jinkela_wire_8292),
        .c(new_Jinkela_wire_8293)
    );

    bfr new_Jinkela_buffer_6659 (
        .din(new_Jinkela_wire_8144),
        .dout(new_Jinkela_wire_8145)
    );

    spl2 new_Jinkela_splitter_616 (
        .a(n_0777_),
        .b(new_Jinkela_wire_8294),
        .c(new_Jinkela_wire_8295)
    );

    bfr new_Jinkela_buffer_6690 (
        .din(new_Jinkela_wire_8211),
        .dout(new_Jinkela_wire_8212)
    );

    bfr new_Jinkela_buffer_6660 (
        .din(new_Jinkela_wire_8145),
        .dout(new_Jinkela_wire_8146)
    );

    bfr new_Jinkela_buffer_6744 (
        .din(new_Jinkela_wire_8299),
        .dout(new_Jinkela_wire_8300)
    );

    bfr new_Jinkela_buffer_6661 (
        .din(new_Jinkela_wire_8146),
        .dout(new_Jinkela_wire_8147)
    );

    spl2 new_Jinkela_splitter_614 (
        .a(new_Jinkela_wire_8287),
        .b(new_Jinkela_wire_8288),
        .c(new_Jinkela_wire_8289)
    );

    bfr new_Jinkela_buffer_6691 (
        .din(new_Jinkela_wire_8212),
        .dout(new_Jinkela_wire_8213)
    );

    bfr new_Jinkela_buffer_6662 (
        .din(new_Jinkela_wire_8147),
        .dout(new_Jinkela_wire_8148)
    );

    spl2 new_Jinkela_splitter_619 (
        .a(n_0978_),
        .b(new_Jinkela_wire_8301),
        .c(new_Jinkela_wire_8302)
    );

    bfr new_Jinkela_buffer_6663 (
        .din(new_Jinkela_wire_8148),
        .dout(new_Jinkela_wire_8149)
    );

    bfr new_Jinkela_buffer_6692 (
        .din(new_Jinkela_wire_8213),
        .dout(new_Jinkela_wire_8214)
    );

    bfr new_Jinkela_buffer_6664 (
        .din(new_Jinkela_wire_8149),
        .dout(new_Jinkela_wire_8150)
    );

    bfr new_Jinkela_buffer_6665 (
        .din(new_Jinkela_wire_8150),
        .dout(new_Jinkela_wire_8151)
    );

    spl2 new_Jinkela_splitter_617 (
        .a(n_1002_),
        .b(new_Jinkela_wire_8296),
        .c(new_Jinkela_wire_8297)
    );

    bfr new_Jinkela_buffer_6693 (
        .din(new_Jinkela_wire_8214),
        .dout(new_Jinkela_wire_8215)
    );

    bfr new_Jinkela_buffer_6666 (
        .din(new_Jinkela_wire_8151),
        .dout(new_Jinkela_wire_8152)
    );

    bfr new_Jinkela_buffer_6667 (
        .din(new_Jinkela_wire_8152),
        .dout(new_Jinkela_wire_8153)
    );

    bfr new_Jinkela_buffer_6694 (
        .din(new_Jinkela_wire_8215),
        .dout(new_Jinkela_wire_8216)
    );

    bfr new_Jinkela_buffer_6668 (
        .din(new_Jinkela_wire_8153),
        .dout(new_Jinkela_wire_8154)
    );

    spl2 new_Jinkela_splitter_618 (
        .a(n_0226_),
        .b(new_Jinkela_wire_8298),
        .c(new_Jinkela_wire_8299)
    );

    bfr new_Jinkela_buffer_6669 (
        .din(new_Jinkela_wire_8154),
        .dout(new_Jinkela_wire_8155)
    );

    bfr new_Jinkela_buffer_6695 (
        .din(new_Jinkela_wire_8216),
        .dout(new_Jinkela_wire_8217)
    );

    bfr new_Jinkela_buffer_6670 (
        .din(new_Jinkela_wire_8155),
        .dout(new_Jinkela_wire_8156)
    );

    bfr new_Jinkela_buffer_6671 (
        .din(new_Jinkela_wire_8156),
        .dout(new_Jinkela_wire_8157)
    );

    bfr new_Jinkela_buffer_6745 (
        .din(n_0050_),
        .dout(new_Jinkela_wire_8303)
    );

    bfr new_Jinkela_buffer_6696 (
        .din(new_Jinkela_wire_8217),
        .dout(new_Jinkela_wire_8218)
    );

    bfr new_Jinkela_buffer_6672 (
        .din(new_Jinkela_wire_8157),
        .dout(new_Jinkela_wire_8158)
    );

    bfr new_Jinkela_buffer_6746 (
        .din(new_Jinkela_wire_8303),
        .dout(new_Jinkela_wire_8304)
    );

    bfr new_Jinkela_buffer_6673 (
        .din(new_Jinkela_wire_8158),
        .dout(new_Jinkela_wire_8159)
    );

    bfr new_Jinkela_buffer_6697 (
        .din(new_Jinkela_wire_8218),
        .dout(new_Jinkela_wire_8219)
    );

    spl2 new_Jinkela_splitter_590 (
        .a(new_Jinkela_wire_8159),
        .b(new_Jinkela_wire_8160),
        .c(new_Jinkela_wire_8161)
    );

    bfr new_Jinkela_buffer_6674 (
        .din(new_Jinkela_wire_8161),
        .dout(new_Jinkela_wire_8162)
    );

    bfr new_Jinkela_buffer_6749 (
        .din(n_0567_),
        .dout(new_Jinkela_wire_8309)
    );

    spl2 new_Jinkela_splitter_620 (
        .a(n_0535_),
        .b(new_Jinkela_wire_8307),
        .c(new_Jinkela_wire_8308)
    );

    bfr new_Jinkela_buffer_6698 (
        .din(new_Jinkela_wire_8219),
        .dout(new_Jinkela_wire_8220)
    );

    bfr new_Jinkela_buffer_1668 (
        .din(new_Jinkela_wire_2013),
        .dout(new_Jinkela_wire_2014)
    );

    bfr new_Jinkela_buffer_1618 (
        .din(new_Jinkela_wire_1961),
        .dout(new_Jinkela_wire_1962)
    );

    bfr new_Jinkela_buffer_1619 (
        .din(new_Jinkela_wire_1962),
        .dout(new_Jinkela_wire_1963)
    );

    bfr new_Jinkela_buffer_1733 (
        .din(new_Jinkela_wire_2078),
        .dout(new_Jinkela_wire_2079)
    );

    bfr new_Jinkela_buffer_1669 (
        .din(new_Jinkela_wire_2014),
        .dout(new_Jinkela_wire_2015)
    );

    bfr new_Jinkela_buffer_1620 (
        .din(new_Jinkela_wire_1963),
        .dout(new_Jinkela_wire_1964)
    );

    bfr new_Jinkela_buffer_1621 (
        .din(new_Jinkela_wire_1964),
        .dout(new_Jinkela_wire_1965)
    );

    bfr new_Jinkela_buffer_1806 (
        .din(N227),
        .dout(new_Jinkela_wire_2157)
    );

    bfr new_Jinkela_buffer_1670 (
        .din(new_Jinkela_wire_2015),
        .dout(new_Jinkela_wire_2016)
    );

    bfr new_Jinkela_buffer_1622 (
        .din(new_Jinkela_wire_1965),
        .dout(new_Jinkela_wire_1966)
    );

    bfr new_Jinkela_buffer_1623 (
        .din(new_Jinkela_wire_1966),
        .dout(new_Jinkela_wire_1967)
    );

    bfr new_Jinkela_buffer_1734 (
        .din(new_Jinkela_wire_2079),
        .dout(new_Jinkela_wire_2080)
    );

    bfr new_Jinkela_buffer_1671 (
        .din(new_Jinkela_wire_2016),
        .dout(new_Jinkela_wire_2017)
    );

    bfr new_Jinkela_buffer_1624 (
        .din(new_Jinkela_wire_1967),
        .dout(new_Jinkela_wire_1968)
    );

    bfr new_Jinkela_buffer_1625 (
        .din(new_Jinkela_wire_1968),
        .dout(new_Jinkela_wire_1969)
    );

    bfr new_Jinkela_buffer_1672 (
        .din(new_Jinkela_wire_2017),
        .dout(new_Jinkela_wire_2018)
    );

    bfr new_Jinkela_buffer_1626 (
        .din(new_Jinkela_wire_1969),
        .dout(new_Jinkela_wire_1970)
    );

    bfr new_Jinkela_buffer_1810 (
        .din(N236),
        .dout(new_Jinkela_wire_2161)
    );

    bfr new_Jinkela_buffer_1627 (
        .din(new_Jinkela_wire_1970),
        .dout(new_Jinkela_wire_1971)
    );

    bfr new_Jinkela_buffer_1737 (
        .din(new_Jinkela_wire_2082),
        .dout(new_Jinkela_wire_2083)
    );

    bfr new_Jinkela_buffer_1673 (
        .din(new_Jinkela_wire_2018),
        .dout(new_Jinkela_wire_2019)
    );

    bfr new_Jinkela_buffer_1628 (
        .din(new_Jinkela_wire_1971),
        .dout(new_Jinkela_wire_1972)
    );

    bfr new_Jinkela_buffer_1800 (
        .din(new_Jinkela_wire_2150),
        .dout(new_Jinkela_wire_2151)
    );

    bfr new_Jinkela_buffer_1629 (
        .din(new_Jinkela_wire_1972),
        .dout(new_Jinkela_wire_1973)
    );

    bfr new_Jinkela_buffer_1674 (
        .din(new_Jinkela_wire_2019),
        .dout(new_Jinkela_wire_2020)
    );

    bfr new_Jinkela_buffer_1736 (
        .din(new_Jinkela_wire_2081),
        .dout(new_Jinkela_wire_2082)
    );

    spl2 new_Jinkela_splitter_110 (
        .a(new_Jinkela_wire_2083),
        .b(new_Jinkela_wire_2084),
        .c(new_Jinkela_wire_2085)
    );

    bfr new_Jinkela_buffer_1675 (
        .din(new_Jinkela_wire_2020),
        .dout(new_Jinkela_wire_2021)
    );

    bfr new_Jinkela_buffer_1738 (
        .din(new_Jinkela_wire_2085),
        .dout(new_Jinkela_wire_2086)
    );

    bfr new_Jinkela_buffer_1676 (
        .din(new_Jinkela_wire_2021),
        .dout(new_Jinkela_wire_2022)
    );

    bfr new_Jinkela_buffer_1677 (
        .din(new_Jinkela_wire_2022),
        .dout(new_Jinkela_wire_2023)
    );

    bfr new_Jinkela_buffer_1801 (
        .din(new_Jinkela_wire_2151),
        .dout(new_Jinkela_wire_2152)
    );

    bfr new_Jinkela_buffer_1678 (
        .din(new_Jinkela_wire_2023),
        .dout(new_Jinkela_wire_2024)
    );

    bfr new_Jinkela_buffer_1807 (
        .din(new_Jinkela_wire_2157),
        .dout(new_Jinkela_wire_2158)
    );

    bfr new_Jinkela_buffer_1679 (
        .din(new_Jinkela_wire_2024),
        .dout(new_Jinkela_wire_2025)
    );

    bfr new_Jinkela_buffer_1739 (
        .din(new_Jinkela_wire_2086),
        .dout(new_Jinkela_wire_2087)
    );

    bfr new_Jinkela_buffer_1680 (
        .din(new_Jinkela_wire_2025),
        .dout(new_Jinkela_wire_2026)
    );

    bfr new_Jinkela_buffer_1802 (
        .din(new_Jinkela_wire_2152),
        .dout(new_Jinkela_wire_2153)
    );

    bfr new_Jinkela_buffer_1681 (
        .din(new_Jinkela_wire_2026),
        .dout(new_Jinkela_wire_2027)
    );

    bfr new_Jinkela_buffer_1740 (
        .din(new_Jinkela_wire_2087),
        .dout(new_Jinkela_wire_2088)
    );

    bfr new_Jinkela_buffer_1682 (
        .din(new_Jinkela_wire_2027),
        .dout(new_Jinkela_wire_2028)
    );

    bfr new_Jinkela_buffer_116 (
        .din(new_Jinkela_wire_127),
        .dout(new_Jinkela_wire_128)
    );

    spl2 new_Jinkela_splitter_280 (
        .a(n_0856_),
        .b(new_Jinkela_wire_4984),
        .c(new_Jinkela_wire_4985)
    );

    bfr new_Jinkela_buffer_181 (
        .din(new_Jinkela_wire_196),
        .dout(new_Jinkela_wire_197)
    );

    bfr new_Jinkela_buffer_4178 (
        .din(new_Jinkela_wire_4899),
        .dout(new_Jinkela_wire_4900)
    );

    bfr new_Jinkela_buffer_117 (
        .din(new_Jinkela_wire_128),
        .dout(new_Jinkela_wire_129)
    );

    bfr new_Jinkela_buffer_4201 (
        .din(new_Jinkela_wire_4934),
        .dout(new_Jinkela_wire_4935)
    );

    bfr new_Jinkela_buffer_179 (
        .din(new_Jinkela_wire_194),
        .dout(new_Jinkela_wire_195)
    );

    bfr new_Jinkela_buffer_4179 (
        .din(new_Jinkela_wire_4900),
        .dout(new_Jinkela_wire_4901)
    );

    bfr new_Jinkela_buffer_118 (
        .din(new_Jinkela_wire_129),
        .dout(new_Jinkela_wire_130)
    );

    bfr new_Jinkela_buffer_4230 (
        .din(n_1142_),
        .dout(new_Jinkela_wire_4986)
    );

    bfr new_Jinkela_buffer_4180 (
        .din(new_Jinkela_wire_4901),
        .dout(new_Jinkela_wire_4902)
    );

    bfr new_Jinkela_buffer_184 (
        .din(new_Jinkela_wire_201),
        .dout(new_Jinkela_wire_202)
    );

    bfr new_Jinkela_buffer_119 (
        .din(new_Jinkela_wire_130),
        .dout(new_Jinkela_wire_131)
    );

    bfr new_Jinkela_buffer_4202 (
        .din(new_Jinkela_wire_4935),
        .dout(new_Jinkela_wire_4936)
    );

    bfr new_Jinkela_buffer_182 (
        .din(new_Jinkela_wire_197),
        .dout(new_Jinkela_wire_198)
    );

    bfr new_Jinkela_buffer_4181 (
        .din(new_Jinkela_wire_4902),
        .dout(new_Jinkela_wire_4903)
    );

    bfr new_Jinkela_buffer_120 (
        .din(new_Jinkela_wire_131),
        .dout(new_Jinkela_wire_132)
    );

    bfr new_Jinkela_buffer_4225 (
        .din(n_1350_),
        .dout(new_Jinkela_wire_4977)
    );

    bfr new_Jinkela_buffer_4226 (
        .din(new_Jinkela_wire_4977),
        .dout(new_Jinkela_wire_4978)
    );

    bfr new_Jinkela_buffer_249 (
        .din(new_Jinkela_wire_268),
        .dout(new_Jinkela_wire_269)
    );

    bfr new_Jinkela_buffer_4182 (
        .din(new_Jinkela_wire_4903),
        .dout(new_Jinkela_wire_4904)
    );

    bfr new_Jinkela_buffer_252 (
        .din(N319),
        .dout(new_Jinkela_wire_272)
    );

    bfr new_Jinkela_buffer_121 (
        .din(new_Jinkela_wire_132),
        .dout(new_Jinkela_wire_133)
    );

    bfr new_Jinkela_buffer_4203 (
        .din(new_Jinkela_wire_4936),
        .dout(new_Jinkela_wire_4937)
    );

    bfr new_Jinkela_buffer_183 (
        .din(new_Jinkela_wire_198),
        .dout(new_Jinkela_wire_199)
    );

    bfr new_Jinkela_buffer_4183 (
        .din(new_Jinkela_wire_4904),
        .dout(new_Jinkela_wire_4905)
    );

    bfr new_Jinkela_buffer_122 (
        .din(new_Jinkela_wire_133),
        .dout(new_Jinkela_wire_134)
    );

    bfr new_Jinkela_buffer_4231 (
        .din(new_Jinkela_wire_4986),
        .dout(new_Jinkela_wire_4987)
    );

    bfr new_Jinkela_buffer_4184 (
        .din(new_Jinkela_wire_4905),
        .dout(new_Jinkela_wire_4906)
    );

    bfr new_Jinkela_buffer_123 (
        .din(new_Jinkela_wire_134),
        .dout(new_Jinkela_wire_135)
    );

    bfr new_Jinkela_buffer_4204 (
        .din(new_Jinkela_wire_4937),
        .dout(new_Jinkela_wire_4938)
    );

    bfr new_Jinkela_buffer_4185 (
        .din(new_Jinkela_wire_4906),
        .dout(new_Jinkela_wire_4907)
    );

    bfr new_Jinkela_buffer_124 (
        .din(new_Jinkela_wire_135),
        .dout(new_Jinkela_wire_136)
    );

    bfr new_Jinkela_buffer_4227 (
        .din(new_Jinkela_wire_4978),
        .dout(new_Jinkela_wire_4979)
    );

    bfr new_Jinkela_buffer_185 (
        .din(new_Jinkela_wire_202),
        .dout(new_Jinkela_wire_203)
    );

    bfr new_Jinkela_buffer_4186 (
        .din(new_Jinkela_wire_4907),
        .dout(new_Jinkela_wire_4908)
    );

    bfr new_Jinkela_buffer_125 (
        .din(new_Jinkela_wire_136),
        .dout(new_Jinkela_wire_137)
    );

    bfr new_Jinkela_buffer_4205 (
        .din(new_Jinkela_wire_4938),
        .dout(new_Jinkela_wire_4939)
    );

    bfr new_Jinkela_buffer_4187 (
        .din(new_Jinkela_wire_4908),
        .dout(new_Jinkela_wire_4909)
    );

    bfr new_Jinkela_buffer_126 (
        .din(new_Jinkela_wire_137),
        .dout(new_Jinkela_wire_138)
    );

    spl2 new_Jinkela_splitter_282 (
        .a(n_0921_),
        .b(new_Jinkela_wire_4997),
        .c(new_Jinkela_wire_4998)
    );

    spl2 new_Jinkela_splitter_8 (
        .a(new_Jinkela_wire_203),
        .b(new_Jinkela_wire_204),
        .c(new_Jinkela_wire_205)
    );

    bfr new_Jinkela_buffer_4188 (
        .din(new_Jinkela_wire_4909),
        .dout(new_Jinkela_wire_4910)
    );

    bfr new_Jinkela_buffer_127 (
        .din(new_Jinkela_wire_138),
        .dout(new_Jinkela_wire_139)
    );

    bfr new_Jinkela_buffer_4206 (
        .din(new_Jinkela_wire_4939),
        .dout(new_Jinkela_wire_4940)
    );

    bfr new_Jinkela_buffer_186 (
        .din(new_Jinkela_wire_205),
        .dout(new_Jinkela_wire_206)
    );

    bfr new_Jinkela_buffer_4189 (
        .din(new_Jinkela_wire_4910),
        .dout(new_Jinkela_wire_4911)
    );

    bfr new_Jinkela_buffer_128 (
        .din(new_Jinkela_wire_139),
        .dout(new_Jinkela_wire_140)
    );

    bfr new_Jinkela_buffer_4234 (
        .din(n_0670_),
        .dout(new_Jinkela_wire_4990)
    );

    bfr new_Jinkela_buffer_4228 (
        .din(new_Jinkela_wire_4979),
        .dout(new_Jinkela_wire_4980)
    );

    bfr new_Jinkela_buffer_250 (
        .din(new_Jinkela_wire_269),
        .dout(new_Jinkela_wire_270)
    );

    spl2 new_Jinkela_splitter_268 (
        .a(new_Jinkela_wire_4911),
        .b(new_Jinkela_wire_4912),
        .c(new_Jinkela_wire_4913)
    );

    bfr new_Jinkela_buffer_129 (
        .din(new_Jinkela_wire_140),
        .dout(new_Jinkela_wire_141)
    );

    bfr new_Jinkela_buffer_253 (
        .din(new_Jinkela_wire_272),
        .dout(new_Jinkela_wire_273)
    );

    bfr new_Jinkela_buffer_4207 (
        .din(new_Jinkela_wire_4940),
        .dout(new_Jinkela_wire_4941)
    );

    bfr new_Jinkela_buffer_130 (
        .din(new_Jinkela_wire_141),
        .dout(new_Jinkela_wire_142)
    );

    bfr new_Jinkela_buffer_4208 (
        .din(new_Jinkela_wire_4941),
        .dout(new_Jinkela_wire_4942)
    );

    bfr new_Jinkela_buffer_187 (
        .din(new_Jinkela_wire_206),
        .dout(new_Jinkela_wire_207)
    );

    bfr new_Jinkela_buffer_4229 (
        .din(new_Jinkela_wire_4980),
        .dout(new_Jinkela_wire_4981)
    );

    bfr new_Jinkela_buffer_131 (
        .din(new_Jinkela_wire_142),
        .dout(new_Jinkela_wire_143)
    );

    bfr new_Jinkela_buffer_4209 (
        .din(new_Jinkela_wire_4942),
        .dout(new_Jinkela_wire_4943)
    );

    bfr new_Jinkela_buffer_251 (
        .din(new_Jinkela_wire_270),
        .dout(new_Jinkela_wire_271)
    );

    bfr new_Jinkela_buffer_4239 (
        .din(new_net_2529),
        .dout(new_Jinkela_wire_4999)
    );

    bfr new_Jinkela_buffer_132 (
        .din(new_Jinkela_wire_143),
        .dout(new_Jinkela_wire_144)
    );

    bfr new_Jinkela_buffer_4210 (
        .din(new_Jinkela_wire_4943),
        .dout(new_Jinkela_wire_4944)
    );

    bfr new_Jinkela_buffer_188 (
        .din(new_Jinkela_wire_207),
        .dout(new_Jinkela_wire_208)
    );

    bfr new_Jinkela_buffer_4232 (
        .din(new_Jinkela_wire_4987),
        .dout(new_Jinkela_wire_4988)
    );

    spl2 new_Jinkela_splitter_279 (
        .a(new_Jinkela_wire_4981),
        .b(new_Jinkela_wire_4982),
        .c(new_Jinkela_wire_4983)
    );

    bfr new_Jinkela_buffer_133 (
        .din(new_Jinkela_wire_144),
        .dout(new_Jinkela_wire_145)
    );

    bfr new_Jinkela_buffer_4211 (
        .din(new_Jinkela_wire_4944),
        .dout(new_Jinkela_wire_4945)
    );

    bfr new_Jinkela_buffer_320 (
        .din(N156),
        .dout(new_Jinkela_wire_345)
    );

    bfr new_Jinkela_buffer_4235 (
        .din(new_Jinkela_wire_4990),
        .dout(new_Jinkela_wire_4991)
    );

    bfr new_Jinkela_buffer_134 (
        .din(new_Jinkela_wire_145),
        .dout(new_Jinkela_wire_146)
    );

    bfr new_Jinkela_buffer_4212 (
        .din(new_Jinkela_wire_4945),
        .dout(new_Jinkela_wire_4946)
    );

    bfr new_Jinkela_buffer_189 (
        .din(new_Jinkela_wire_208),
        .dout(new_Jinkela_wire_209)
    );

    bfr new_Jinkela_buffer_4233 (
        .din(new_Jinkela_wire_4988),
        .dout(new_Jinkela_wire_4989)
    );

    bfr new_Jinkela_buffer_135 (
        .din(new_Jinkela_wire_146),
        .dout(new_Jinkela_wire_147)
    );

    bfr new_Jinkela_buffer_4213 (
        .din(new_Jinkela_wire_4946),
        .dout(new_Jinkela_wire_4947)
    );

    bfr new_Jinkela_buffer_317 (
        .din(new_Jinkela_wire_341),
        .dout(new_Jinkela_wire_342)
    );

    bfr new_Jinkela_buffer_316 (
        .din(N59),
        .dout(new_Jinkela_wire_341)
    );

    bfr new_Jinkela_buffer_136 (
        .din(new_Jinkela_wire_147),
        .dout(new_Jinkela_wire_148)
    );

    bfr new_Jinkela_buffer_4214 (
        .din(new_Jinkela_wire_4947),
        .dout(new_Jinkela_wire_4948)
    );

    bfr new_Jinkela_buffer_190 (
        .din(new_Jinkela_wire_209),
        .dout(new_Jinkela_wire_210)
    );

    and_bi n_2622_ (
        .a(new_Jinkela_wire_4239),
        .b(new_Jinkela_wire_4870),
        .c(n_0480_)
    );

    bfr new_Jinkela_buffer_2509 (
        .din(new_Jinkela_wire_2910),
        .dout(new_Jinkela_wire_2911)
    );

    and_bb n_1905_ (
        .a(new_Jinkela_wire_4653),
        .b(new_Jinkela_wire_7073),
        .c(n_1171_)
    );

    and_bi n_2623_ (
        .a(new_Jinkela_wire_4869),
        .b(new_Jinkela_wire_4238),
        .c(n_0481_)
    );

    bfr new_Jinkela_buffer_2452 (
        .din(new_Jinkela_wire_2853),
        .dout(new_Jinkela_wire_2854)
    );

    and_ii n_1906_ (
        .a(new_Jinkela_wire_4652),
        .b(new_Jinkela_wire_7072),
        .c(n_1172_)
    );

    bfr new_Jinkela_buffer_5856 (
        .din(new_Jinkela_wire_7060),
        .dout(new_Jinkela_wire_7061)
    );

    and_ii n_2624_ (
        .a(n_0481_),
        .b(n_0480_),
        .c(n_0482_)
    );

    and_ii n_1907_ (
        .a(n_1172_),
        .b(n_1171_),
        .c(n_1173_)
    );

    bfr new_Jinkela_buffer_2640 (
        .din(new_Jinkela_wire_3045),
        .dout(new_Jinkela_wire_3046)
    );

    bfr new_Jinkela_buffer_5875 (
        .din(new_Jinkela_wire_7107),
        .dout(new_Jinkela_wire_7108)
    );

    and_bb n_2625_ (
        .a(new_Jinkela_wire_9657),
        .b(new_Jinkela_wire_7545),
        .c(n_0483_)
    );

    bfr new_Jinkela_buffer_2453 (
        .din(new_Jinkela_wire_2854),
        .dout(new_Jinkela_wire_2855)
    );

    and_bi n_1908_ (
        .a(new_Jinkela_wire_7833),
        .b(new_Jinkela_wire_7298),
        .c(n_1174_)
    );

    bfr new_Jinkela_buffer_5857 (
        .din(new_Jinkela_wire_7061),
        .dout(new_Jinkela_wire_7062)
    );

    and_ii n_2626_ (
        .a(new_Jinkela_wire_8539),
        .b(new_Jinkela_wire_9140),
        .c(n_0484_)
    );

    bfr new_Jinkela_buffer_2510 (
        .din(new_Jinkela_wire_2911),
        .dout(new_Jinkela_wire_2912)
    );

    and_bi n_1909_ (
        .a(new_Jinkela_wire_7297),
        .b(new_Jinkela_wire_7832),
        .c(n_1175_)
    );

    spl2 new_Jinkela_splitter_487 (
        .a(n_0344_),
        .b(new_Jinkela_wire_7205),
        .c(new_Jinkela_wire_7206)
    );

    and_bi n_2627_ (
        .a(new_Jinkela_wire_6197),
        .b(new_Jinkela_wire_7548),
        .c(n_0485_)
    );

    bfr new_Jinkela_buffer_2454 (
        .din(new_Jinkela_wire_2855),
        .dout(new_Jinkela_wire_2856)
    );

    bfr new_Jinkela_buffer_5885 (
        .din(new_Jinkela_wire_7124),
        .dout(new_Jinkela_wire_7125)
    );

    and_ii n_1910_ (
        .a(n_1175_),
        .b(n_1174_),
        .c(n_1176_)
    );

    bfr new_Jinkela_buffer_5858 (
        .din(new_Jinkela_wire_7062),
        .dout(new_Jinkela_wire_7063)
    );

    and_ii n_2628_ (
        .a(new_Jinkela_wire_8265),
        .b(new_Jinkela_wire_9582),
        .c(n_0486_)
    );

    bfr new_Jinkela_buffer_2573 (
        .din(new_Jinkela_wire_2974),
        .dout(new_Jinkela_wire_2975)
    );

    and_bb n_1911_ (
        .a(new_Jinkela_wire_3346),
        .b(new_Jinkela_wire_1210),
        .c(n_1177_)
    );

    bfr new_Jinkela_buffer_5876 (
        .din(new_Jinkela_wire_7108),
        .dout(new_Jinkela_wire_7109)
    );

    and_bi n_2629_ (
        .a(new_Jinkela_wire_9583),
        .b(new_Jinkela_wire_5569),
        .c(n_0487_)
    );

    bfr new_Jinkela_buffer_2455 (
        .din(new_Jinkela_wire_2856),
        .dout(new_Jinkela_wire_2857)
    );

    and_ii n_1912_ (
        .a(new_Jinkela_wire_5287),
        .b(new_Jinkela_wire_8998),
        .c(n_1178_)
    );

    bfr new_Jinkela_buffer_5859 (
        .din(new_Jinkela_wire_7063),
        .dout(new_Jinkela_wire_7064)
    );

    or_bb n_2630_ (
        .a(n_0487_),
        .b(n_0486_),
        .c(n_0488_)
    );

    bfr new_Jinkela_buffer_2511 (
        .din(new_Jinkela_wire_2912),
        .dout(new_Jinkela_wire_2913)
    );

    and_bb n_1913_ (
        .a(new_Jinkela_wire_1778),
        .b(new_Jinkela_wire_1304),
        .c(n_1179_)
    );

    and_bi n_2631_ (
        .a(new_Jinkela_wire_5678),
        .b(new_Jinkela_wire_4542),
        .c(n_0489_)
    );

    bfr new_Jinkela_buffer_2456 (
        .din(new_Jinkela_wire_2857),
        .dout(new_Jinkela_wire_2858)
    );

    bfr new_Jinkela_buffer_5948 (
        .din(new_Jinkela_wire_7189),
        .dout(new_Jinkela_wire_7190)
    );

    and_ii n_1914_ (
        .a(new_Jinkela_wire_9394),
        .b(new_Jinkela_wire_6517),
        .c(n_1180_)
    );

    bfr new_Jinkela_buffer_5860 (
        .din(new_Jinkela_wire_7064),
        .dout(new_Jinkela_wire_7065)
    );

    and_bi n_2632_ (
        .a(new_Jinkela_wire_4541),
        .b(new_Jinkela_wire_5679),
        .c(n_0490_)
    );

    bfr new_Jinkela_buffer_2707 (
        .din(N75),
        .dout(new_Jinkela_wire_3117)
    );

    and_ii n_1915_ (
        .a(new_Jinkela_wire_8186),
        .b(new_Jinkela_wire_7278),
        .c(n_1181_)
    );

    spl2 new_Jinkela_splitter_136 (
        .a(N325),
        .b(new_Jinkela_wire_3049),
        .c(new_Jinkela_wire_3050)
    );

    bfr new_Jinkela_buffer_5877 (
        .din(new_Jinkela_wire_7109),
        .dout(new_Jinkela_wire_7110)
    );

    or_bb n_2633_ (
        .a(n_0490_),
        .b(n_0489_),
        .c(n_0491_)
    );

    bfr new_Jinkela_buffer_2457 (
        .din(new_Jinkela_wire_2858),
        .dout(new_Jinkela_wire_2859)
    );

    and_bb n_1916_ (
        .a(new_Jinkela_wire_8185),
        .b(new_Jinkela_wire_7279),
        .c(n_1182_)
    );

    bfr new_Jinkela_buffer_5861 (
        .din(new_Jinkela_wire_7065),
        .dout(new_Jinkela_wire_7066)
    );

    and_ii n_2634_ (
        .a(new_Jinkela_wire_9892),
        .b(new_Jinkela_wire_9600),
        .c(n_0492_)
    );

    bfr new_Jinkela_buffer_2512 (
        .din(new_Jinkela_wire_2913),
        .dout(new_Jinkela_wire_2914)
    );

    and_ii n_1917_ (
        .a(n_1182_),
        .b(n_1181_),
        .c(n_1183_)
    );

    spl2 new_Jinkela_splitter_484 (
        .a(new_Jinkela_wire_7186),
        .b(new_Jinkela_wire_7187),
        .c(new_Jinkela_wire_7188)
    );

    and_bb n_2635_ (
        .a(new_Jinkela_wire_9891),
        .b(new_Jinkela_wire_9599),
        .c(n_0493_)
    );

    bfr new_Jinkela_buffer_2458 (
        .din(new_Jinkela_wire_2859),
        .dout(new_Jinkela_wire_2860)
    );

    bfr new_Jinkela_buffer_5886 (
        .din(new_Jinkela_wire_7125),
        .dout(new_Jinkela_wire_7126)
    );

    and_bb n_1918_ (
        .a(new_Jinkela_wire_1798),
        .b(new_Jinkela_wire_1246),
        .c(n_1184_)
    );

    bfr new_Jinkela_buffer_5878 (
        .din(new_Jinkela_wire_7110),
        .dout(new_Jinkela_wire_7111)
    );

    and_ii n_2636_ (
        .a(n_0493_),
        .b(n_0492_),
        .c(n_0494_)
    );

    and_ii n_1919_ (
        .a(new_Jinkela_wire_9385),
        .b(new_Jinkela_wire_4534),
        .c(n_1185_)
    );

    bfr new_Jinkela_buffer_2575 (
        .din(new_Jinkela_wire_2980),
        .dout(new_Jinkela_wire_2981)
    );

    and_bb n_2637_ (
        .a(new_Jinkela_wire_5416),
        .b(new_Jinkela_wire_6789),
        .c(n_0495_)
    );

    bfr new_Jinkela_buffer_2459 (
        .din(new_Jinkela_wire_2860),
        .dout(new_Jinkela_wire_2861)
    );

    and_bb n_1920_ (
        .a(new_Jinkela_wire_2971),
        .b(new_Jinkela_wire_1198),
        .c(n_1186_)
    );

    bfr new_Jinkela_buffer_5879 (
        .din(new_Jinkela_wire_7111),
        .dout(new_Jinkela_wire_7112)
    );

    and_ii n_2638_ (
        .a(new_Jinkela_wire_5415),
        .b(new_Jinkela_wire_6788),
        .c(n_0496_)
    );

    bfr new_Jinkela_buffer_2513 (
        .din(new_Jinkela_wire_2914),
        .dout(new_Jinkela_wire_2915)
    );

    and_ii n_1921_ (
        .a(new_Jinkela_wire_8450),
        .b(new_Jinkela_wire_8275),
        .c(n_1187_)
    );

    bfr new_Jinkela_buffer_5968 (
        .din(n_1321_),
        .dout(new_Jinkela_wire_7217)
    );

    or_bb n_2639_ (
        .a(n_0496_),
        .b(n_0495_),
        .c(n_0497_)
    );

    bfr new_Jinkela_buffer_2460 (
        .din(new_Jinkela_wire_2861),
        .dout(new_Jinkela_wire_2862)
    );

    bfr new_Jinkela_buffer_5887 (
        .din(new_Jinkela_wire_7126),
        .dout(new_Jinkela_wire_7127)
    );

    and_bb n_1922_ (
        .a(new_Jinkela_wire_6392),
        .b(new_Jinkela_wire_6673),
        .c(n_1188_)
    );

    bfr new_Jinkela_buffer_5880 (
        .din(new_Jinkela_wire_7112),
        .dout(new_Jinkela_wire_7113)
    );

    and_bi n_2640_ (
        .a(new_Jinkela_wire_5143),
        .b(new_Jinkela_wire_6086),
        .c(n_0498_)
    );

    and_ii n_1923_ (
        .a(new_Jinkela_wire_6390),
        .b(new_Jinkela_wire_6672),
        .c(n_1189_)
    );

    and_bi n_2641_ (
        .a(new_Jinkela_wire_6435),
        .b(new_Jinkela_wire_8264),
        .c(n_0499_)
    );

    bfr new_Jinkela_buffer_2461 (
        .din(new_Jinkela_wire_2862),
        .dout(new_Jinkela_wire_2863)
    );

    bfr new_Jinkela_buffer_5949 (
        .din(new_Jinkela_wire_7190),
        .dout(new_Jinkela_wire_7191)
    );

    and_ii n_1924_ (
        .a(n_1189_),
        .b(n_1188_),
        .c(n_1190_)
    );

    and_ii n_2642_ (
        .a(new_Jinkela_wire_9141),
        .b(new_Jinkela_wire_8945),
        .c(n_0500_)
    );

    bfr new_Jinkela_buffer_2514 (
        .din(new_Jinkela_wire_2915),
        .dout(new_Jinkela_wire_2916)
    );

    bfr new_Jinkela_buffer_5888 (
        .din(new_Jinkela_wire_7127),
        .dout(new_Jinkela_wire_7128)
    );

    and_bi n_1925_ (
        .a(new_Jinkela_wire_6430),
        .b(new_Jinkela_wire_7384),
        .c(n_1191_)
    );

    and_bi n_2643_ (
        .a(new_Jinkela_wire_9605),
        .b(new_Jinkela_wire_5681),
        .c(n_0501_)
    );

    bfr new_Jinkela_buffer_2462 (
        .din(new_Jinkela_wire_2863),
        .dout(new_Jinkela_wire_2864)
    );

    and_bi n_1926_ (
        .a(new_Jinkela_wire_7383),
        .b(new_Jinkela_wire_6429),
        .c(n_1192_)
    );

    and_bi n_2644_ (
        .a(new_Jinkela_wire_5682),
        .b(new_Jinkela_wire_9604),
        .c(n_0502_)
    );

    bfr new_Jinkela_buffer_5889 (
        .din(new_Jinkela_wire_7128),
        .dout(new_Jinkela_wire_7129)
    );

    and_ii n_1927_ (
        .a(n_1192_),
        .b(n_1191_),
        .c(n_1193_)
    );

    bfr new_Jinkela_buffer_2576 (
        .din(new_Jinkela_wire_2981),
        .dout(new_Jinkela_wire_2982)
    );

    and_ii n_2645_ (
        .a(n_0502_),
        .b(n_0501_),
        .c(n_0503_)
    );

    bfr new_Jinkela_buffer_2463 (
        .din(new_Jinkela_wire_2864),
        .dout(new_Jinkela_wire_2865)
    );

    and_bi n_1928_ (
        .a(new_Jinkela_wire_6838),
        .b(new_Jinkela_wire_3717),
        .c(n_1194_)
    );

    bfr new_Jinkela_buffer_5973 (
        .din(n_1326_),
        .dout(new_Jinkela_wire_7224)
    );

    and_bi n_2646_ (
        .a(new_Jinkela_wire_6538),
        .b(new_Jinkela_wire_6198),
        .c(n_0504_)
    );

    bfr new_Jinkela_buffer_2515 (
        .din(new_Jinkela_wire_2916),
        .dout(new_Jinkela_wire_2917)
    );

    bfr new_Jinkela_buffer_5890 (
        .din(new_Jinkela_wire_7129),
        .dout(new_Jinkela_wire_7130)
    );

    and_bi n_1929_ (
        .a(new_Jinkela_wire_3716),
        .b(new_Jinkela_wire_6837),
        .c(n_1195_)
    );

    and_bi n_2647_ (
        .a(new_Jinkela_wire_6193),
        .b(new_Jinkela_wire_6537),
        .c(n_0505_)
    );

    bfr new_Jinkela_buffer_2464 (
        .din(new_Jinkela_wire_2865),
        .dout(new_Jinkela_wire_2866)
    );

    bfr new_Jinkela_buffer_5950 (
        .din(new_Jinkela_wire_7191),
        .dout(new_Jinkela_wire_7192)
    );

    or_bb n_1930_ (
        .a(n_1195_),
        .b(n_1194_),
        .c(n_1196_)
    );

    and_ii n_2648_ (
        .a(n_0505_),
        .b(n_0504_),
        .c(n_0506_)
    );

    bfr new_Jinkela_buffer_5891 (
        .din(new_Jinkela_wire_7130),
        .dout(new_Jinkela_wire_7131)
    );

    or_bb n_1931_ (
        .a(n_1196_),
        .b(new_Jinkela_wire_3592),
        .c(n_1197_)
    );

    bfr new_Jinkela_buffer_2643 (
        .din(new_Jinkela_wire_3050),
        .dout(new_Jinkela_wire_3051)
    );

    and_bi n_2649_ (
        .a(new_Jinkela_wire_10145),
        .b(new_Jinkela_wire_9138),
        .c(n_0507_)
    );

    bfr new_Jinkela_buffer_2465 (
        .din(new_Jinkela_wire_2866),
        .dout(new_Jinkela_wire_2867)
    );

    spl2 new_Jinkela_splitter_486 (
        .a(new_Jinkela_wire_7202),
        .b(new_Jinkela_wire_7203),
        .c(new_Jinkela_wire_7204)
    );

    and_bb n_1932_ (
        .a(new_Jinkela_wire_1802),
        .b(new_Jinkela_wire_1272),
        .c(n_1198_)
    );

    bfr new_Jinkela_buffer_5958 (
        .din(new_Jinkela_wire_7206),
        .dout(new_Jinkela_wire_7207)
    );

    and_bi n_2650_ (
        .a(new_Jinkela_wire_9139),
        .b(new_Jinkela_wire_10144),
        .c(n_0508_)
    );

    bfr new_Jinkela_buffer_2516 (
        .din(new_Jinkela_wire_2917),
        .dout(new_Jinkela_wire_2918)
    );

    bfr new_Jinkela_buffer_5892 (
        .din(new_Jinkela_wire_7131),
        .dout(new_Jinkela_wire_7132)
    );

    and_ii n_1933_ (
        .a(new_Jinkela_wire_5554),
        .b(new_Jinkela_wire_7340),
        .c(n_1199_)
    );

    or_bb n_2651_ (
        .a(n_0508_),
        .b(n_0507_),
        .c(n_0509_)
    );

    bfr new_Jinkela_buffer_2466 (
        .din(new_Jinkela_wire_2867),
        .dout(new_Jinkela_wire_2868)
    );

    bfr new_Jinkela_buffer_5951 (
        .din(new_Jinkela_wire_7192),
        .dout(new_Jinkela_wire_7193)
    );

    and_bb n_1934_ (
        .a(new_Jinkela_wire_3197),
        .b(new_Jinkela_wire_1369),
        .c(n_1200_)
    );

    and_bi n_2652_ (
        .a(new_Jinkela_wire_4530),
        .b(new_Jinkela_wire_9831),
        .c(n_0510_)
    );

    bfr new_Jinkela_buffer_2641 (
        .din(new_Jinkela_wire_3046),
        .dout(new_Jinkela_wire_3047)
    );

    bfr new_Jinkela_buffer_5893 (
        .din(new_Jinkela_wire_7132),
        .dout(new_Jinkela_wire_7133)
    );

    and_ii n_1935_ (
        .a(new_Jinkela_wire_10342),
        .b(new_Jinkela_wire_6515),
        .c(n_1201_)
    );

    bfr new_Jinkela_buffer_2577 (
        .din(new_Jinkela_wire_2982),
        .dout(new_Jinkela_wire_2983)
    );

    or_bb n_2653_ (
        .a(n_0510_),
        .b(n_0498_),
        .c(n_0511_)
    );

    bfr new_Jinkela_buffer_2467 (
        .din(new_Jinkela_wire_2868),
        .dout(new_Jinkela_wire_2869)
    );

    and_bi n_1936_ (
        .a(new_Jinkela_wire_3861),
        .b(new_Jinkela_wire_3714),
        .c(n_1202_)
    );

    or_bb n_2654_ (
        .a(new_Jinkela_wire_9481),
        .b(new_Jinkela_wire_7727),
        .c(n_0512_)
    );

    bfr new_Jinkela_buffer_2517 (
        .din(new_Jinkela_wire_2918),
        .dout(new_Jinkela_wire_2919)
    );

    bfr new_Jinkela_buffer_5894 (
        .din(new_Jinkela_wire_7133),
        .dout(new_Jinkela_wire_7134)
    );

    and_bi n_1937_ (
        .a(new_Jinkela_wire_3712),
        .b(new_Jinkela_wire_3860),
        .c(n_1203_)
    );

    and_bb n_2655_ (
        .a(new_Jinkela_wire_9480),
        .b(new_Jinkela_wire_7726),
        .c(n_0513_)
    );

    bfr new_Jinkela_buffer_2468 (
        .din(new_Jinkela_wire_2869),
        .dout(new_Jinkela_wire_2870)
    );

    bfr new_Jinkela_buffer_5952 (
        .din(new_Jinkela_wire_7193),
        .dout(new_Jinkela_wire_7194)
    );

    or_bb n_1938_ (
        .a(n_1203_),
        .b(n_1202_),
        .c(n_1204_)
    );

    and_bi n_2656_ (
        .a(n_0512_),
        .b(n_0513_),
        .c(n_0514_)
    );

    bfr new_Jinkela_buffer_5895 (
        .din(new_Jinkela_wire_7134),
        .dout(new_Jinkela_wire_7135)
    );

    and_bi n_1939_ (
        .a(new_Jinkela_wire_1299),
        .b(new_Jinkela_wire_87),
        .c(n_1205_)
    );

    or_bi n_2657_ (
        .a(new_Jinkela_wire_5934),
        .b(new_Jinkela_wire_7740),
        .c(n_0515_)
    );

    bfr new_Jinkela_buffer_2469 (
        .din(new_Jinkela_wire_2870),
        .dout(new_Jinkela_wire_2871)
    );

    and_ii n_1940_ (
        .a(new_Jinkela_wire_3838),
        .b(new_Jinkela_wire_9452),
        .c(n_1206_)
    );

    and_bi n_2658_ (
        .a(new_Jinkela_wire_5933),
        .b(new_Jinkela_wire_7739),
        .c(n_0516_)
    );

    bfr new_Jinkela_buffer_2518 (
        .din(new_Jinkela_wire_2919),
        .dout(new_Jinkela_wire_2920)
    );

    bfr new_Jinkela_buffer_5896 (
        .din(new_Jinkela_wire_7135),
        .dout(new_Jinkela_wire_7136)
    );

    and_bi n_1941_ (
        .a(new_Jinkela_wire_1214),
        .b(new_Jinkela_wire_2377),
        .c(n_1207_)
    );

    and_bi n_2659_ (
        .a(n_0515_),
        .b(n_0516_),
        .c(new_net_2529)
    );

    bfr new_Jinkela_buffer_2470 (
        .din(new_Jinkela_wire_2871),
        .dout(new_Jinkela_wire_2872)
    );

    bfr new_Jinkela_buffer_5953 (
        .din(new_Jinkela_wire_7194),
        .dout(new_Jinkela_wire_7195)
    );

    and_bb n_1942_ (
        .a(new_Jinkela_wire_3786),
        .b(new_Jinkela_wire_6314),
        .c(n_1208_)
    );

    and_bb n_2660_ (
        .a(new_Jinkela_wire_4307),
        .b(new_Jinkela_wire_3779),
        .c(n_0517_)
    );

    bfr new_Jinkela_buffer_5897 (
        .din(new_Jinkela_wire_7136),
        .dout(new_Jinkela_wire_7137)
    );

    and_ii n_1943_ (
        .a(new_Jinkela_wire_3783),
        .b(new_Jinkela_wire_9449),
        .c(n_1209_)
    );

    bfr new_Jinkela_buffer_2578 (
        .din(new_Jinkela_wire_2983),
        .dout(new_Jinkela_wire_2984)
    );

    and_ii n_2661_ (
        .a(new_Jinkela_wire_5559),
        .b(new_Jinkela_wire_8707),
        .c(n_0518_)
    );

    bfr new_Jinkela_buffer_2471 (
        .din(new_Jinkela_wire_2872),
        .dout(new_Jinkela_wire_2873)
    );

    bfr new_Jinkela_buffer_5974 (
        .din(n_1300_),
        .dout(new_Jinkela_wire_7227)
    );

    and_bb n_1944_ (
        .a(new_Jinkela_wire_9475),
        .b(new_Jinkela_wire_3841),
        .c(n_1210_)
    );

    bfr new_Jinkela_buffer_5959 (
        .din(new_Jinkela_wire_7207),
        .dout(new_Jinkela_wire_7208)
    );

    and_bb n_2662_ (
        .a(new_Jinkela_wire_9776),
        .b(new_Jinkela_wire_3792),
        .c(n_0519_)
    );

    bfr new_Jinkela_buffer_2519 (
        .din(new_Jinkela_wire_2920),
        .dout(new_Jinkela_wire_2921)
    );

    bfr new_Jinkela_buffer_5898 (
        .din(new_Jinkela_wire_7137),
        .dout(new_Jinkela_wire_7138)
    );

    and_ii n_1945_ (
        .a(n_1210_),
        .b(n_1208_),
        .c(n_1211_)
    );

    or_bb n_2663_ (
        .a(n_0519_),
        .b(n_0518_),
        .c(n_0520_)
    );

    bfr new_Jinkela_buffer_2472 (
        .din(new_Jinkela_wire_2873),
        .dout(new_Jinkela_wire_2874)
    );

    bfr new_Jinkela_buffer_5954 (
        .din(new_Jinkela_wire_7195),
        .dout(new_Jinkela_wire_7196)
    );

    and_bi n_1946_ (
        .a(new_Jinkela_wire_1337),
        .b(new_Jinkela_wire_2236),
        .c(n_1212_)
    );

    bfr new_Jinkela_buffer_3350 (
        .din(new_Jinkela_wire_3884),
        .dout(new_Jinkela_wire_3885)
    );

    bfr new_Jinkela_buffer_137 (
        .din(new_Jinkela_wire_148),
        .dout(new_Jinkela_wire_149)
    );

    spl2 new_Jinkela_splitter_369 (
        .a(new_Jinkela_wire_6005),
        .b(new_Jinkela_wire_6006),
        .c(new_Jinkela_wire_6007)
    );

    bfr new_Jinkela_buffer_3378 (
        .din(new_Jinkela_wire_3915),
        .dout(new_Jinkela_wire_3916)
    );

    bfr new_Jinkela_buffer_254 (
        .din(new_Jinkela_wire_273),
        .dout(new_Jinkela_wire_274)
    );

    bfr new_Jinkela_buffer_5052 (
        .din(new_Jinkela_wire_6027),
        .dout(new_Jinkela_wire_6028)
    );

    bfr new_Jinkela_buffer_3351 (
        .din(new_Jinkela_wire_3885),
        .dout(new_Jinkela_wire_3886)
    );

    bfr new_Jinkela_buffer_138 (
        .din(new_Jinkela_wire_149),
        .dout(new_Jinkela_wire_150)
    );

    bfr new_Jinkela_buffer_5110 (
        .din(new_Jinkela_wire_6089),
        .dout(new_Jinkela_wire_6090)
    );

    bfr new_Jinkela_buffer_3385 (
        .din(new_Jinkela_wire_3929),
        .dout(new_Jinkela_wire_3930)
    );

    bfr new_Jinkela_buffer_191 (
        .din(new_Jinkela_wire_210),
        .dout(new_Jinkela_wire_211)
    );

    bfr new_Jinkela_buffer_5088 (
        .din(new_Jinkela_wire_6065),
        .dout(new_Jinkela_wire_6066)
    );

    spl3L new_Jinkela_splitter_191 (
        .a(new_Jinkela_wire_3923),
        .d(new_Jinkela_wire_3924),
        .b(new_Jinkela_wire_3925),
        .c(new_Jinkela_wire_3926)
    );

    bfr new_Jinkela_buffer_3352 (
        .din(new_Jinkela_wire_3886),
        .dout(new_Jinkela_wire_3887)
    );

    bfr new_Jinkela_buffer_139 (
        .din(new_Jinkela_wire_150),
        .dout(new_Jinkela_wire_151)
    );

    bfr new_Jinkela_buffer_5053 (
        .din(new_Jinkela_wire_6028),
        .dout(new_Jinkela_wire_6029)
    );

    bfr new_Jinkela_buffer_3379 (
        .din(new_Jinkela_wire_3916),
        .dout(new_Jinkela_wire_3917)
    );

    bfr new_Jinkela_buffer_326 (
        .din(N115),
        .dout(new_Jinkela_wire_356)
    );

    spl2 new_Jinkela_splitter_9 (
        .a(new_Jinkela_wire_274),
        .b(new_Jinkela_wire_275),
        .c(new_Jinkela_wire_276)
    );

    bfr new_Jinkela_buffer_5118 (
        .din(n_0139_),
        .dout(new_Jinkela_wire_6110)
    );

    bfr new_Jinkela_buffer_3353 (
        .din(new_Jinkela_wire_3887),
        .dout(new_Jinkela_wire_3888)
    );

    bfr new_Jinkela_buffer_140 (
        .din(new_Jinkela_wire_151),
        .dout(new_Jinkela_wire_152)
    );

    bfr new_Jinkela_buffer_5089 (
        .din(new_Jinkela_wire_6066),
        .dout(new_Jinkela_wire_6067)
    );

    bfr new_Jinkela_buffer_5054 (
        .din(new_Jinkela_wire_6029),
        .dout(new_Jinkela_wire_6030)
    );

    bfr new_Jinkela_buffer_192 (
        .din(new_Jinkela_wire_211),
        .dout(new_Jinkela_wire_212)
    );

    spl2 new_Jinkela_splitter_195 (
        .a(n_0252_),
        .b(new_Jinkela_wire_3942),
        .c(new_Jinkela_wire_3943)
    );

    bfr new_Jinkela_buffer_3354 (
        .din(new_Jinkela_wire_3888),
        .dout(new_Jinkela_wire_3889)
    );

    bfr new_Jinkela_buffer_141 (
        .din(new_Jinkela_wire_152),
        .dout(new_Jinkela_wire_153)
    );

    bfr new_Jinkela_buffer_5055 (
        .din(new_Jinkela_wire_6030),
        .dout(new_Jinkela_wire_6031)
    );

    bfr new_Jinkela_buffer_3380 (
        .din(new_Jinkela_wire_3917),
        .dout(new_Jinkela_wire_3918)
    );

    bfr new_Jinkela_buffer_255 (
        .din(new_Jinkela_wire_276),
        .dout(new_Jinkela_wire_277)
    );

    bfr new_Jinkela_buffer_5111 (
        .din(new_Jinkela_wire_6090),
        .dout(new_Jinkela_wire_6091)
    );

    bfr new_Jinkela_buffer_3355 (
        .din(new_Jinkela_wire_3889),
        .dout(new_Jinkela_wire_3890)
    );

    bfr new_Jinkela_buffer_142 (
        .din(new_Jinkela_wire_153),
        .dout(new_Jinkela_wire_154)
    );

    bfr new_Jinkela_buffer_5090 (
        .din(new_Jinkela_wire_6067),
        .dout(new_Jinkela_wire_6068)
    );

    bfr new_Jinkela_buffer_5056 (
        .din(new_Jinkela_wire_6031),
        .dout(new_Jinkela_wire_6032)
    );

    bfr new_Jinkela_buffer_193 (
        .din(new_Jinkela_wire_212),
        .dout(new_Jinkela_wire_213)
    );

    spl4L new_Jinkela_splitter_194 (
        .a(n_0812_),
        .d(new_Jinkela_wire_3936),
        .b(new_Jinkela_wire_3937),
        .e(new_Jinkela_wire_3938),
        .c(new_Jinkela_wire_3939)
    );

    bfr new_Jinkela_buffer_3356 (
        .din(new_Jinkela_wire_3890),
        .dout(new_Jinkela_wire_3891)
    );

    bfr new_Jinkela_buffer_143 (
        .din(new_Jinkela_wire_154),
        .dout(new_Jinkela_wire_155)
    );

    bfr new_Jinkela_buffer_5057 (
        .din(new_Jinkela_wire_6032),
        .dout(new_Jinkela_wire_6033)
    );

    spl2 new_Jinkela_splitter_189 (
        .a(new_Jinkela_wire_3918),
        .b(new_Jinkela_wire_3919),
        .c(new_Jinkela_wire_3920)
    );

    spl3L new_Jinkela_splitter_11 (
        .a(N38),
        .d(new_Jinkela_wire_349),
        .b(new_Jinkela_wire_350),
        .c(new_Jinkela_wire_351)
    );

    bfr new_Jinkela_buffer_3357 (
        .din(new_Jinkela_wire_3891),
        .dout(new_Jinkela_wire_3892)
    );

    bfr new_Jinkela_buffer_144 (
        .din(new_Jinkela_wire_155),
        .dout(new_Jinkela_wire_156)
    );

    bfr new_Jinkela_buffer_5091 (
        .din(new_Jinkela_wire_6068),
        .dout(new_Jinkela_wire_6069)
    );

    bfr new_Jinkela_buffer_5058 (
        .din(new_Jinkela_wire_6033),
        .dout(new_Jinkela_wire_6034)
    );

    bfr new_Jinkela_buffer_194 (
        .din(new_Jinkela_wire_213),
        .dout(new_Jinkela_wire_214)
    );

    bfr new_Jinkela_buffer_3386 (
        .din(new_Jinkela_wire_3930),
        .dout(new_Jinkela_wire_3931)
    );

    bfr new_Jinkela_buffer_3358 (
        .din(new_Jinkela_wire_3892),
        .dout(new_Jinkela_wire_3893)
    );

    bfr new_Jinkela_buffer_145 (
        .din(new_Jinkela_wire_156),
        .dout(new_Jinkela_wire_157)
    );

    bfr new_Jinkela_buffer_5059 (
        .din(new_Jinkela_wire_6034),
        .dout(new_Jinkela_wire_6035)
    );

    bfr new_Jinkela_buffer_3382 (
        .din(new_Jinkela_wire_3926),
        .dout(new_Jinkela_wire_3927)
    );

    bfr new_Jinkela_buffer_318 (
        .din(new_Jinkela_wire_342),
        .dout(new_Jinkela_wire_343)
    );

    bfr new_Jinkela_buffer_5112 (
        .din(new_Jinkela_wire_6091),
        .dout(new_Jinkela_wire_6092)
    );

    bfr new_Jinkela_buffer_3359 (
        .din(new_Jinkela_wire_3893),
        .dout(new_Jinkela_wire_3894)
    );

    bfr new_Jinkela_buffer_146 (
        .din(new_Jinkela_wire_157),
        .dout(new_Jinkela_wire_158)
    );

    bfr new_Jinkela_buffer_5092 (
        .din(new_Jinkela_wire_6069),
        .dout(new_Jinkela_wire_6070)
    );

    bfr new_Jinkela_buffer_5060 (
        .din(new_Jinkela_wire_6035),
        .dout(new_Jinkela_wire_6036)
    );

    bfr new_Jinkela_buffer_3383 (
        .din(new_Jinkela_wire_3927),
        .dout(new_Jinkela_wire_3928)
    );

    bfr new_Jinkela_buffer_195 (
        .din(new_Jinkela_wire_214),
        .dout(new_Jinkela_wire_215)
    );

    bfr new_Jinkela_buffer_3360 (
        .din(new_Jinkela_wire_3894),
        .dout(new_Jinkela_wire_3895)
    );

    bfr new_Jinkela_buffer_147 (
        .din(new_Jinkela_wire_158),
        .dout(new_Jinkela_wire_159)
    );

    bfr new_Jinkela_buffer_5061 (
        .din(new_Jinkela_wire_6036),
        .dout(new_Jinkela_wire_6037)
    );

    bfr new_Jinkela_buffer_321 (
        .din(new_Jinkela_wire_345),
        .dout(new_Jinkela_wire_346)
    );

    bfr new_Jinkela_buffer_3388 (
        .din(new_Jinkela_wire_3940),
        .dout(new_Jinkela_wire_3941)
    );

    spl2 new_Jinkela_splitter_382 (
        .a(n_0624_),
        .b(new_Jinkela_wire_6130),
        .c(new_Jinkela_wire_6131)
    );

    bfr new_Jinkela_buffer_3361 (
        .din(new_Jinkela_wire_3895),
        .dout(new_Jinkela_wire_3896)
    );

    bfr new_Jinkela_buffer_148 (
        .din(new_Jinkela_wire_159),
        .dout(new_Jinkela_wire_160)
    );

    bfr new_Jinkela_buffer_5093 (
        .din(new_Jinkela_wire_6070),
        .dout(new_Jinkela_wire_6071)
    );

    bfr new_Jinkela_buffer_5062 (
        .din(new_Jinkela_wire_6037),
        .dout(new_Jinkela_wire_6038)
    );

    bfr new_Jinkela_buffer_3387 (
        .din(n_0199_),
        .dout(new_Jinkela_wire_3940)
    );

    bfr new_Jinkela_buffer_196 (
        .din(new_Jinkela_wire_215),
        .dout(new_Jinkela_wire_216)
    );

    spl2 new_Jinkela_splitter_192 (
        .a(new_Jinkela_wire_3931),
        .b(new_Jinkela_wire_3932),
        .c(new_Jinkela_wire_3933)
    );

    bfr new_Jinkela_buffer_3362 (
        .din(new_Jinkela_wire_3896),
        .dout(new_Jinkela_wire_3897)
    );

    bfr new_Jinkela_buffer_149 (
        .din(new_Jinkela_wire_160),
        .dout(new_Jinkela_wire_161)
    );

    spl2 new_Jinkela_splitter_380 (
        .a(new_Jinkela_wire_6107),
        .b(new_Jinkela_wire_6108),
        .c(new_Jinkela_wire_6109)
    );

    bfr new_Jinkela_buffer_5063 (
        .din(new_Jinkela_wire_6038),
        .dout(new_Jinkela_wire_6039)
    );

    bfr new_Jinkela_buffer_256 (
        .din(new_Jinkela_wire_277),
        .dout(new_Jinkela_wire_278)
    );

    bfr new_Jinkela_buffer_3389 (
        .din(n_1204_),
        .dout(new_Jinkela_wire_3944)
    );

    bfr new_Jinkela_buffer_5113 (
        .din(new_Jinkela_wire_6092),
        .dout(new_Jinkela_wire_6093)
    );

    bfr new_Jinkela_buffer_3363 (
        .din(new_Jinkela_wire_3897),
        .dout(new_Jinkela_wire_3898)
    );

    bfr new_Jinkela_buffer_150 (
        .din(new_Jinkela_wire_161),
        .dout(new_Jinkela_wire_162)
    );

    bfr new_Jinkela_buffer_5094 (
        .din(new_Jinkela_wire_6071),
        .dout(new_Jinkela_wire_6072)
    );

    bfr new_Jinkela_buffer_5064 (
        .din(new_Jinkela_wire_6039),
        .dout(new_Jinkela_wire_6040)
    );

    bfr new_Jinkela_buffer_197 (
        .din(new_Jinkela_wire_216),
        .dout(new_Jinkela_wire_217)
    );

    bfr new_Jinkela_buffer_3392 (
        .din(new_net_2531),
        .dout(new_Jinkela_wire_3954)
    );

    bfr new_Jinkela_buffer_3364 (
        .din(new_Jinkela_wire_3898),
        .dout(new_Jinkela_wire_3899)
    );

    bfr new_Jinkela_buffer_151 (
        .din(new_Jinkela_wire_162),
        .dout(new_Jinkela_wire_163)
    );

    bfr new_Jinkela_buffer_5065 (
        .din(new_Jinkela_wire_6040),
        .dout(new_Jinkela_wire_6041)
    );

    bfr new_Jinkela_buffer_319 (
        .din(new_Jinkela_wire_343),
        .dout(new_Jinkela_wire_344)
    );

    spl2 new_Jinkela_splitter_198 (
        .a(new_Jinkela_wire_3951),
        .b(new_Jinkela_wire_3952),
        .c(new_Jinkela_wire_3953)
    );

    bfr new_Jinkela_buffer_5117 (
        .din(new_Jinkela_wire_6101),
        .dout(new_Jinkela_wire_6102)
    );

    bfr new_Jinkela_buffer_3365 (
        .din(new_Jinkela_wire_3899),
        .dout(new_Jinkela_wire_3900)
    );

    bfr new_Jinkela_buffer_152 (
        .din(new_Jinkela_wire_163),
        .dout(new_Jinkela_wire_164)
    );

    bfr new_Jinkela_buffer_5095 (
        .din(new_Jinkela_wire_6072),
        .dout(new_Jinkela_wire_6073)
    );

    bfr new_Jinkela_buffer_5066 (
        .din(new_Jinkela_wire_6041),
        .dout(new_Jinkela_wire_6042)
    );

    bfr new_Jinkela_buffer_198 (
        .din(new_Jinkela_wire_217),
        .dout(new_Jinkela_wire_218)
    );

    bfr new_Jinkela_buffer_3366 (
        .din(new_Jinkela_wire_3900),
        .dout(new_Jinkela_wire_3901)
    );

    bfr new_Jinkela_buffer_153 (
        .din(new_Jinkela_wire_164),
        .dout(new_Jinkela_wire_165)
    );

    spl2 new_Jinkela_splitter_378 (
        .a(new_Jinkela_wire_6102),
        .b(new_Jinkela_wire_6103),
        .c(new_Jinkela_wire_6104)
    );

    bfr new_Jinkela_buffer_5067 (
        .din(new_Jinkela_wire_6042),
        .dout(new_Jinkela_wire_6043)
    );

    spl3L new_Jinkela_splitter_197 (
        .a(n_1018_),
        .d(new_Jinkela_wire_3949),
        .b(new_Jinkela_wire_3950),
        .c(new_Jinkela_wire_3951)
    );

    bfr new_Jinkela_buffer_257 (
        .din(new_Jinkela_wire_278),
        .dout(new_Jinkela_wire_279)
    );

    bfr new_Jinkela_buffer_3390 (
        .din(new_Jinkela_wire_3944),
        .dout(new_Jinkela_wire_3945)
    );

    bfr new_Jinkela_buffer_5114 (
        .din(new_Jinkela_wire_6093),
        .dout(new_Jinkela_wire_6094)
    );

    bfr new_Jinkela_buffer_3367 (
        .din(new_Jinkela_wire_3901),
        .dout(new_Jinkela_wire_3902)
    );

    bfr new_Jinkela_buffer_154 (
        .din(new_Jinkela_wire_165),
        .dout(new_Jinkela_wire_166)
    );

    bfr new_Jinkela_buffer_5096 (
        .din(new_Jinkela_wire_6073),
        .dout(new_Jinkela_wire_6074)
    );

    bfr new_Jinkela_buffer_5068 (
        .din(new_Jinkela_wire_6043),
        .dout(new_Jinkela_wire_6044)
    );

    bfr new_Jinkela_buffer_199 (
        .din(new_Jinkela_wire_218),
        .dout(new_Jinkela_wire_219)
    );

    bfr new_Jinkela_buffer_3368 (
        .din(new_Jinkela_wire_3902),
        .dout(new_Jinkela_wire_3903)
    );

    bfr new_Jinkela_buffer_155 (
        .din(new_Jinkela_wire_166),
        .dout(new_Jinkela_wire_167)
    );

    bfr new_Jinkela_buffer_5069 (
        .din(new_Jinkela_wire_6044),
        .dout(new_Jinkela_wire_6045)
    );

    bfr new_Jinkela_buffer_3391 (
        .din(new_Jinkela_wire_3945),
        .dout(new_Jinkela_wire_3946)
    );

    bfr new_Jinkela_buffer_3369 (
        .din(new_Jinkela_wire_3903),
        .dout(new_Jinkela_wire_3904)
    );

    bfr new_Jinkela_buffer_156 (
        .din(new_Jinkela_wire_167),
        .dout(new_Jinkela_wire_168)
    );

    bfr new_Jinkela_buffer_5097 (
        .din(new_Jinkela_wire_6074),
        .dout(new_Jinkela_wire_6075)
    );

    bfr new_Jinkela_buffer_5070 (
        .din(new_Jinkela_wire_6045),
        .dout(new_Jinkela_wire_6046)
    );

    bfr new_Jinkela_buffer_200 (
        .din(new_Jinkela_wire_219),
        .dout(new_Jinkela_wire_220)
    );

    spl3L new_Jinkela_splitter_199 (
        .a(n_0963_),
        .d(new_Jinkela_wire_4007),
        .b(new_Jinkela_wire_4008),
        .c(new_Jinkela_wire_4009)
    );

    bfr new_Jinkela_buffer_3370 (
        .din(new_Jinkela_wire_3904),
        .dout(new_Jinkela_wire_3905)
    );

    bfr new_Jinkela_buffer_157 (
        .din(new_Jinkela_wire_168),
        .dout(new_Jinkela_wire_169)
    );

    bfr new_Jinkela_buffer_5071 (
        .din(new_Jinkela_wire_6046),
        .dout(new_Jinkela_wire_6047)
    );

    spl2 new_Jinkela_splitter_201 (
        .a(n_0075_),
        .b(new_Jinkela_wire_4012),
        .c(new_Jinkela_wire_4013)
    );

    spl3L new_Jinkela_splitter_10 (
        .a(new_Jinkela_wire_279),
        .d(new_Jinkela_wire_280),
        .b(new_Jinkela_wire_281),
        .c(new_Jinkela_wire_282)
    );

    spl2 new_Jinkela_splitter_196 (
        .a(new_Jinkela_wire_3946),
        .b(new_Jinkela_wire_3947),
        .c(new_Jinkela_wire_3948)
    );

    bfr new_Jinkela_buffer_5115 (
        .din(new_Jinkela_wire_6094),
        .dout(new_Jinkela_wire_6095)
    );

    spl2 new_Jinkela_splitter_112 (
        .a(N331),
        .b(new_Jinkela_wire_2165),
        .c(new_Jinkela_wire_2166)
    );

    bfr new_Jinkela_buffer_1683 (
        .din(new_Jinkela_wire_2028),
        .dout(new_Jinkela_wire_2029)
    );

    bfr new_Jinkela_buffer_1878 (
        .din(N176),
        .dout(new_Jinkela_wire_2233)
    );

    spl3L new_Jinkela_splitter_111 (
        .a(new_Jinkela_wire_2088),
        .d(new_Jinkela_wire_2089),
        .b(new_Jinkela_wire_2090),
        .c(new_Jinkela_wire_2091)
    );

    bfr new_Jinkela_buffer_1684 (
        .din(new_Jinkela_wire_2029),
        .dout(new_Jinkela_wire_2030)
    );

    bfr new_Jinkela_buffer_1803 (
        .din(new_Jinkela_wire_2153),
        .dout(new_Jinkela_wire_2154)
    );

    bfr new_Jinkela_buffer_1685 (
        .din(new_Jinkela_wire_2030),
        .dout(new_Jinkela_wire_2031)
    );

    bfr new_Jinkela_buffer_1741 (
        .din(new_Jinkela_wire_2091),
        .dout(new_Jinkela_wire_2092)
    );

    bfr new_Jinkela_buffer_1686 (
        .din(new_Jinkela_wire_2031),
        .dout(new_Jinkela_wire_2032)
    );

    bfr new_Jinkela_buffer_1808 (
        .din(new_Jinkela_wire_2158),
        .dout(new_Jinkela_wire_2159)
    );

    bfr new_Jinkela_buffer_1687 (
        .din(new_Jinkela_wire_2032),
        .dout(new_Jinkela_wire_2033)
    );

    bfr new_Jinkela_buffer_1742 (
        .din(new_Jinkela_wire_2092),
        .dout(new_Jinkela_wire_2093)
    );

    bfr new_Jinkela_buffer_1688 (
        .din(new_Jinkela_wire_2033),
        .dout(new_Jinkela_wire_2034)
    );

    bfr new_Jinkela_buffer_1804 (
        .din(new_Jinkela_wire_2154),
        .dout(new_Jinkela_wire_2155)
    );

    bfr new_Jinkela_buffer_1689 (
        .din(new_Jinkela_wire_2034),
        .dout(new_Jinkela_wire_2035)
    );

    bfr new_Jinkela_buffer_1743 (
        .din(new_Jinkela_wire_2093),
        .dout(new_Jinkela_wire_2094)
    );

    bfr new_Jinkela_buffer_1690 (
        .din(new_Jinkela_wire_2035),
        .dout(new_Jinkela_wire_2036)
    );

    bfr new_Jinkela_buffer_1811 (
        .din(new_Jinkela_wire_2161),
        .dout(new_Jinkela_wire_2162)
    );

    bfr new_Jinkela_buffer_1691 (
        .din(new_Jinkela_wire_2036),
        .dout(new_Jinkela_wire_2037)
    );

    bfr new_Jinkela_buffer_1744 (
        .din(new_Jinkela_wire_2094),
        .dout(new_Jinkela_wire_2095)
    );

    bfr new_Jinkela_buffer_1692 (
        .din(new_Jinkela_wire_2037),
        .dout(new_Jinkela_wire_2038)
    );

    bfr new_Jinkela_buffer_1805 (
        .din(new_Jinkela_wire_2155),
        .dout(new_Jinkela_wire_2156)
    );

    bfr new_Jinkela_buffer_1693 (
        .din(new_Jinkela_wire_2038),
        .dout(new_Jinkela_wire_2039)
    );

    bfr new_Jinkela_buffer_1745 (
        .din(new_Jinkela_wire_2095),
        .dout(new_Jinkela_wire_2096)
    );

    bfr new_Jinkela_buffer_1694 (
        .din(new_Jinkela_wire_2039),
        .dout(new_Jinkela_wire_2040)
    );

    bfr new_Jinkela_buffer_1809 (
        .din(new_Jinkela_wire_2159),
        .dout(new_Jinkela_wire_2160)
    );

    bfr new_Jinkela_buffer_1695 (
        .din(new_Jinkela_wire_2040),
        .dout(new_Jinkela_wire_2041)
    );

    bfr new_Jinkela_buffer_1746 (
        .din(new_Jinkela_wire_2096),
        .dout(new_Jinkela_wire_2097)
    );

    bfr new_Jinkela_buffer_1696 (
        .din(new_Jinkela_wire_2041),
        .dout(new_Jinkela_wire_2042)
    );

    bfr new_Jinkela_buffer_1697 (
        .din(new_Jinkela_wire_2042),
        .dout(new_Jinkela_wire_2043)
    );

    bfr new_Jinkela_buffer_1814 (
        .din(new_Jinkela_wire_2166),
        .dout(new_Jinkela_wire_2167)
    );

    bfr new_Jinkela_buffer_1747 (
        .din(new_Jinkela_wire_2097),
        .dout(new_Jinkela_wire_2098)
    );

    bfr new_Jinkela_buffer_1698 (
        .din(new_Jinkela_wire_2043),
        .dout(new_Jinkela_wire_2044)
    );

    bfr new_Jinkela_buffer_1812 (
        .din(new_Jinkela_wire_2162),
        .dout(new_Jinkela_wire_2163)
    );

    bfr new_Jinkela_buffer_1699 (
        .din(new_Jinkela_wire_2044),
        .dout(new_Jinkela_wire_2045)
    );

    bfr new_Jinkela_buffer_1748 (
        .din(new_Jinkela_wire_2098),
        .dout(new_Jinkela_wire_2099)
    );

    bfr new_Jinkela_buffer_1700 (
        .din(new_Jinkela_wire_2045),
        .dout(new_Jinkela_wire_2046)
    );

    bfr new_Jinkela_buffer_1701 (
        .din(new_Jinkela_wire_2046),
        .dout(new_Jinkela_wire_2047)
    );

    bfr new_Jinkela_buffer_1749 (
        .din(new_Jinkela_wire_2099),
        .dout(new_Jinkela_wire_2100)
    );

    bfr new_Jinkela_buffer_1702 (
        .din(new_Jinkela_wire_2047),
        .dout(new_Jinkela_wire_2048)
    );

    bfr new_Jinkela_buffer_1813 (
        .din(new_Jinkela_wire_2163),
        .dout(new_Jinkela_wire_2164)
    );

    bfr new_Jinkela_buffer_1703 (
        .din(new_Jinkela_wire_2048),
        .dout(new_Jinkela_wire_2049)
    );

    bfr new_Jinkela_buffer_4215 (
        .din(new_Jinkela_wire_4948),
        .dout(new_Jinkela_wire_4949)
    );

    bfr new_Jinkela_buffer_4246 (
        .din(n_0218_),
        .dout(new_Jinkela_wire_5012)
    );

    bfr new_Jinkela_buffer_4236 (
        .din(new_Jinkela_wire_4991),
        .dout(new_Jinkela_wire_4992)
    );

    bfr new_Jinkela_buffer_4216 (
        .din(new_Jinkela_wire_4949),
        .dout(new_Jinkela_wire_4950)
    );

    spl2 new_Jinkela_splitter_283 (
        .a(n_1024_),
        .b(new_Jinkela_wire_5000),
        .c(new_Jinkela_wire_5001)
    );

    bfr new_Jinkela_buffer_4217 (
        .din(new_Jinkela_wire_4950),
        .dout(new_Jinkela_wire_4951)
    );

    bfr new_Jinkela_buffer_4240 (
        .din(n_0551_),
        .dout(new_Jinkela_wire_5002)
    );

    bfr new_Jinkela_buffer_4237 (
        .din(new_Jinkela_wire_4992),
        .dout(new_Jinkela_wire_4993)
    );

    bfr new_Jinkela_buffer_4218 (
        .din(new_Jinkela_wire_4951),
        .dout(new_Jinkela_wire_4952)
    );

    spl2 new_Jinkela_splitter_285 (
        .a(n_0996_),
        .b(new_Jinkela_wire_5010),
        .c(new_Jinkela_wire_5011)
    );

    bfr new_Jinkela_buffer_4219 (
        .din(new_Jinkela_wire_4952),
        .dout(new_Jinkela_wire_4953)
    );

    bfr new_Jinkela_buffer_4238 (
        .din(new_Jinkela_wire_4993),
        .dout(new_Jinkela_wire_4994)
    );

    bfr new_Jinkela_buffer_4220 (
        .din(new_Jinkela_wire_4953),
        .dout(new_Jinkela_wire_4954)
    );

    bfr new_Jinkela_buffer_4221 (
        .din(new_Jinkela_wire_4954),
        .dout(new_Jinkela_wire_4955)
    );

    bfr new_Jinkela_buffer_4243 (
        .din(n_0237_),
        .dout(new_Jinkela_wire_5007)
    );

    spl2 new_Jinkela_splitter_281 (
        .a(new_Jinkela_wire_4994),
        .b(new_Jinkela_wire_4995),
        .c(new_Jinkela_wire_4996)
    );

    bfr new_Jinkela_buffer_4222 (
        .din(new_Jinkela_wire_4955),
        .dout(new_Jinkela_wire_4956)
    );

    bfr new_Jinkela_buffer_4244 (
        .din(new_Jinkela_wire_5007),
        .dout(new_Jinkela_wire_5008)
    );

    bfr new_Jinkela_buffer_4241 (
        .din(new_Jinkela_wire_5002),
        .dout(new_Jinkela_wire_5003)
    );

    bfr new_Jinkela_buffer_4242 (
        .din(new_Jinkela_wire_5003),
        .dout(new_Jinkela_wire_5004)
    );

    bfr new_Jinkela_buffer_4285 (
        .din(n_1274_),
        .dout(new_Jinkela_wire_5054)
    );

    spl2 new_Jinkela_splitter_284 (
        .a(new_Jinkela_wire_5004),
        .b(new_Jinkela_wire_5005),
        .c(new_Jinkela_wire_5006)
    );

    bfr new_Jinkela_buffer_4245 (
        .din(new_Jinkela_wire_5008),
        .dout(new_Jinkela_wire_5009)
    );

    spl3L new_Jinkela_splitter_286 (
        .a(n_0032_),
        .d(new_Jinkela_wire_5013),
        .b(new_Jinkela_wire_5014),
        .c(new_Jinkela_wire_5015)
    );

    spl4L new_Jinkela_splitter_287 (
        .a(n_0738_),
        .d(new_Jinkela_wire_5055),
        .b(new_Jinkela_wire_5056),
        .e(new_Jinkela_wire_5057),
        .c(new_Jinkela_wire_5058)
    );

    bfr new_Jinkela_buffer_4247 (
        .din(new_Jinkela_wire_5015),
        .dout(new_Jinkela_wire_5016)
    );

    spl2 new_Jinkela_splitter_288 (
        .a(n_1135_),
        .b(new_Jinkela_wire_5059),
        .c(new_Jinkela_wire_5060)
    );

    bfr new_Jinkela_buffer_4248 (
        .din(new_Jinkela_wire_5016),
        .dout(new_Jinkela_wire_5017)
    );

    spl2 new_Jinkela_splitter_289 (
        .a(n_0326_),
        .b(new_Jinkela_wire_5063),
        .c(new_Jinkela_wire_5064)
    );

    bfr new_Jinkela_buffer_4288 (
        .din(new_Jinkela_wire_5064),
        .dout(new_Jinkela_wire_5065)
    );

    bfr new_Jinkela_buffer_4249 (
        .din(new_Jinkela_wire_5017),
        .dout(new_Jinkela_wire_5018)
    );

    bfr new_Jinkela_buffer_4250 (
        .din(new_Jinkela_wire_5018),
        .dout(new_Jinkela_wire_5019)
    );

    bfr new_Jinkela_buffer_4286 (
        .din(new_Jinkela_wire_5060),
        .dout(new_Jinkela_wire_5061)
    );

    spl2 new_Jinkela_splitter_290 (
        .a(n_0832_),
        .b(new_Jinkela_wire_5067),
        .c(new_Jinkela_wire_5068)
    );

    bfr new_Jinkela_buffer_4251 (
        .din(new_Jinkela_wire_5019),
        .dout(new_Jinkela_wire_5020)
    );

    bfr new_Jinkela_buffer_4252 (
        .din(new_Jinkela_wire_5020),
        .dout(new_Jinkela_wire_5021)
    );

    bfr new_Jinkela_buffer_4287 (
        .din(new_Jinkela_wire_5061),
        .dout(new_Jinkela_wire_5062)
    );

    bfr new_Jinkela_buffer_4253 (
        .din(new_Jinkela_wire_5021),
        .dout(new_Jinkela_wire_5022)
    );

    spl2 new_Jinkela_splitter_291 (
        .a(n_1361_),
        .b(new_Jinkela_wire_5069),
        .c(new_Jinkela_wire_5070)
    );

    spl2 new_Jinkela_splitter_292 (
        .a(n_0933_),
        .b(new_Jinkela_wire_5071),
        .c(new_Jinkela_wire_5072)
    );

    bfr new_Jinkela_buffer_4254 (
        .din(new_Jinkela_wire_5022),
        .dout(new_Jinkela_wire_5023)
    );

    bfr new_Jinkela_buffer_4255 (
        .din(new_Jinkela_wire_5023),
        .dout(new_Jinkela_wire_5024)
    );

    bfr new_Jinkela_buffer_4289 (
        .din(new_Jinkela_wire_5065),
        .dout(new_Jinkela_wire_5066)
    );

    bfr new_Jinkela_buffer_158 (
        .din(new_Jinkela_wire_169),
        .dout(new_Jinkela_wire_170)
    );

    bfr new_Jinkela_buffer_2711 (
        .din(N303),
        .dout(new_Jinkela_wire_3121)
    );

    bfr new_Jinkela_buffer_7732 (
        .din(new_Jinkela_wire_9728),
        .dout(new_Jinkela_wire_9729)
    );

    bfr new_Jinkela_buffer_2473 (
        .din(new_Jinkela_wire_2874),
        .dout(new_Jinkela_wire_2875)
    );

    bfr new_Jinkela_buffer_201 (
        .din(new_Jinkela_wire_220),
        .dout(new_Jinkela_wire_221)
    );

    bfr new_Jinkela_buffer_7707 (
        .din(new_Jinkela_wire_9693),
        .dout(new_Jinkela_wire_9694)
    );

    bfr new_Jinkela_buffer_2520 (
        .din(new_Jinkela_wire_2921),
        .dout(new_Jinkela_wire_2922)
    );

    bfr new_Jinkela_buffer_159 (
        .din(new_Jinkela_wire_170),
        .dout(new_Jinkela_wire_171)
    );

    bfr new_Jinkela_buffer_2474 (
        .din(new_Jinkela_wire_2875),
        .dout(new_Jinkela_wire_2876)
    );

    bfr new_Jinkela_buffer_322 (
        .din(new_Jinkela_wire_346),
        .dout(new_Jinkela_wire_347)
    );

    bfr new_Jinkela_buffer_7741 (
        .din(new_Jinkela_wire_9743),
        .dout(new_Jinkela_wire_9744)
    );

    bfr new_Jinkela_buffer_7708 (
        .din(new_Jinkela_wire_9694),
        .dout(new_Jinkela_wire_9695)
    );

    bfr new_Jinkela_buffer_2642 (
        .din(new_Jinkela_wire_3047),
        .dout(new_Jinkela_wire_3048)
    );

    bfr new_Jinkela_buffer_160 (
        .din(new_Jinkela_wire_171),
        .dout(new_Jinkela_wire_172)
    );

    bfr new_Jinkela_buffer_2579 (
        .din(new_Jinkela_wire_2984),
        .dout(new_Jinkela_wire_2985)
    );

    bfr new_Jinkela_buffer_7733 (
        .din(new_Jinkela_wire_9729),
        .dout(new_Jinkela_wire_9730)
    );

    bfr new_Jinkela_buffer_2475 (
        .din(new_Jinkela_wire_2876),
        .dout(new_Jinkela_wire_2877)
    );

    bfr new_Jinkela_buffer_202 (
        .din(new_Jinkela_wire_221),
        .dout(new_Jinkela_wire_222)
    );

    bfr new_Jinkela_buffer_7709 (
        .din(new_Jinkela_wire_9695),
        .dout(new_Jinkela_wire_9696)
    );

    bfr new_Jinkela_buffer_2521 (
        .din(new_Jinkela_wire_2922),
        .dout(new_Jinkela_wire_2923)
    );

    bfr new_Jinkela_buffer_258 (
        .din(new_Jinkela_wire_282),
        .dout(new_Jinkela_wire_283)
    );

    bfr new_Jinkela_buffer_2476 (
        .din(new_Jinkela_wire_2877),
        .dout(new_Jinkela_wire_2878)
    );

    bfr new_Jinkela_buffer_203 (
        .din(new_Jinkela_wire_222),
        .dout(new_Jinkela_wire_223)
    );

    spl2 new_Jinkela_splitter_811 (
        .a(n_0854_),
        .b(new_Jinkela_wire_9770),
        .c(new_Jinkela_wire_9771)
    );

    bfr new_Jinkela_buffer_7710 (
        .din(new_Jinkela_wire_9696),
        .dout(new_Jinkela_wire_9697)
    );

    bfr new_Jinkela_buffer_395 (
        .din(N87),
        .dout(new_Jinkela_wire_427)
    );

    bfr new_Jinkela_buffer_7734 (
        .din(new_Jinkela_wire_9730),
        .dout(new_Jinkela_wire_9731)
    );

    bfr new_Jinkela_buffer_2477 (
        .din(new_Jinkela_wire_2878),
        .dout(new_Jinkela_wire_2879)
    );

    bfr new_Jinkela_buffer_204 (
        .din(new_Jinkela_wire_223),
        .dout(new_Jinkela_wire_224)
    );

    spl2 new_Jinkela_splitter_796 (
        .a(new_Jinkela_wire_9697),
        .b(new_Jinkela_wire_9698),
        .c(new_Jinkela_wire_9699)
    );

    bfr new_Jinkela_buffer_2522 (
        .din(new_Jinkela_wire_2923),
        .dout(new_Jinkela_wire_2924)
    );

    bfr new_Jinkela_buffer_259 (
        .din(new_Jinkela_wire_283),
        .dout(new_Jinkela_wire_284)
    );

    bfr new_Jinkela_buffer_7711 (
        .din(new_Jinkela_wire_9699),
        .dout(new_Jinkela_wire_9700)
    );

    bfr new_Jinkela_buffer_2478 (
        .din(new_Jinkela_wire_2879),
        .dout(new_Jinkela_wire_2880)
    );

    bfr new_Jinkela_buffer_205 (
        .din(new_Jinkela_wire_224),
        .dout(new_Jinkela_wire_225)
    );

    spl2 new_Jinkela_splitter_810 (
        .a(n_0593_),
        .b(new_Jinkela_wire_9768),
        .c(new_Jinkela_wire_9769)
    );

    bfr new_Jinkela_buffer_323 (
        .din(new_Jinkela_wire_347),
        .dout(new_Jinkela_wire_348)
    );

    bfr new_Jinkela_buffer_2580 (
        .din(new_Jinkela_wire_2985),
        .dout(new_Jinkela_wire_2986)
    );

    bfr new_Jinkela_buffer_2479 (
        .din(new_Jinkela_wire_2880),
        .dout(new_Jinkela_wire_2881)
    );

    bfr new_Jinkela_buffer_206 (
        .din(new_Jinkela_wire_225),
        .dout(new_Jinkela_wire_226)
    );

    spl3L new_Jinkela_splitter_812 (
        .a(n_1315_),
        .d(new_Jinkela_wire_9772),
        .b(new_Jinkela_wire_9773),
        .c(new_Jinkela_wire_9774)
    );

    spl2 new_Jinkela_splitter_797 (
        .a(new_Jinkela_wire_9700),
        .b(new_Jinkela_wire_9701),
        .c(new_Jinkela_wire_9702)
    );

    bfr new_Jinkela_buffer_2523 (
        .din(new_Jinkela_wire_2924),
        .dout(new_Jinkela_wire_2925)
    );

    bfr new_Jinkela_buffer_260 (
        .din(new_Jinkela_wire_284),
        .dout(new_Jinkela_wire_285)
    );

    bfr new_Jinkela_buffer_7772 (
        .din(new_Jinkela_wire_9804),
        .dout(new_Jinkela_wire_9805)
    );

    bfr new_Jinkela_buffer_2480 (
        .din(new_Jinkela_wire_2881),
        .dout(new_Jinkela_wire_2882)
    );

    bfr new_Jinkela_buffer_207 (
        .din(new_Jinkela_wire_226),
        .dout(new_Jinkela_wire_227)
    );

    bfr new_Jinkela_buffer_7771 (
        .din(n_0509_),
        .dout(new_Jinkela_wire_9804)
    );

    bfr new_Jinkela_buffer_324 (
        .din(new_Jinkela_wire_351),
        .dout(new_Jinkela_wire_352)
    );

    bfr new_Jinkela_buffer_7801 (
        .din(n_1304_),
        .dout(new_Jinkela_wire_9836)
    );

    bfr new_Jinkela_buffer_2481 (
        .din(new_Jinkela_wire_2882),
        .dout(new_Jinkela_wire_2883)
    );

    bfr new_Jinkela_buffer_208 (
        .din(new_Jinkela_wire_227),
        .dout(new_Jinkela_wire_228)
    );

    bfr new_Jinkela_buffer_7799 (
        .din(n_0613_),
        .dout(new_Jinkela_wire_9832)
    );

    bfr new_Jinkela_buffer_7746 (
        .din(new_Jinkela_wire_9774),
        .dout(new_Jinkela_wire_9775)
    );

    bfr new_Jinkela_buffer_2524 (
        .din(new_Jinkela_wire_2925),
        .dout(new_Jinkela_wire_2926)
    );

    bfr new_Jinkela_buffer_261 (
        .din(new_Jinkela_wire_285),
        .dout(new_Jinkela_wire_286)
    );

    bfr new_Jinkela_buffer_2482 (
        .din(new_Jinkela_wire_2883),
        .dout(new_Jinkela_wire_2884)
    );

    bfr new_Jinkela_buffer_209 (
        .din(new_Jinkela_wire_228),
        .dout(new_Jinkela_wire_229)
    );

    spl2 new_Jinkela_splitter_813 (
        .a(new_Jinkela_wire_9775),
        .b(new_Jinkela_wire_9776),
        .c(new_Jinkela_wire_9777)
    );

    bfr new_Jinkela_buffer_2708 (
        .din(new_Jinkela_wire_3117),
        .dout(new_Jinkela_wire_3118)
    );

    bfr new_Jinkela_buffer_327 (
        .din(new_Jinkela_wire_356),
        .dout(new_Jinkela_wire_357)
    );

    bfr new_Jinkela_buffer_325 (
        .din(new_Jinkela_wire_352),
        .dout(new_Jinkela_wire_353)
    );

    bfr new_Jinkela_buffer_2581 (
        .din(new_Jinkela_wire_2986),
        .dout(new_Jinkela_wire_2987)
    );

    bfr new_Jinkela_buffer_7747 (
        .din(new_Jinkela_wire_9777),
        .dout(new_Jinkela_wire_9778)
    );

    bfr new_Jinkela_buffer_2483 (
        .din(new_Jinkela_wire_2884),
        .dout(new_Jinkela_wire_2885)
    );

    bfr new_Jinkela_buffer_210 (
        .din(new_Jinkela_wire_229),
        .dout(new_Jinkela_wire_230)
    );

    bfr new_Jinkela_buffer_7800 (
        .din(new_Jinkela_wire_9832),
        .dout(new_Jinkela_wire_9833)
    );

    bfr new_Jinkela_buffer_2525 (
        .din(new_Jinkela_wire_2926),
        .dout(new_Jinkela_wire_2927)
    );

    bfr new_Jinkela_buffer_262 (
        .din(new_Jinkela_wire_286),
        .dout(new_Jinkela_wire_287)
    );

    bfr new_Jinkela_buffer_7773 (
        .din(new_Jinkela_wire_9805),
        .dout(new_Jinkela_wire_9806)
    );

    bfr new_Jinkela_buffer_211 (
        .din(new_Jinkela_wire_230),
        .dout(new_Jinkela_wire_231)
    );

    spl2 new_Jinkela_splitter_817 (
        .a(n_0780_),
        .b(new_Jinkela_wire_9843),
        .c(new_Jinkela_wire_9844)
    );

    bfr new_Jinkela_buffer_2526 (
        .din(new_Jinkela_wire_2927),
        .dout(new_Jinkela_wire_2928)
    );

    bfr new_Jinkela_buffer_330 (
        .din(N337),
        .dout(new_Jinkela_wire_360)
    );

    spl2 new_Jinkela_splitter_814 (
        .a(new_Jinkela_wire_9778),
        .b(new_Jinkela_wire_9779),
        .c(new_Jinkela_wire_9780)
    );

    bfr new_Jinkela_buffer_2644 (
        .din(new_Jinkela_wire_3051),
        .dout(new_Jinkela_wire_3052)
    );

    bfr new_Jinkela_buffer_212 (
        .din(new_Jinkela_wire_231),
        .dout(new_Jinkela_wire_232)
    );

    bfr new_Jinkela_buffer_7748 (
        .din(new_Jinkela_wire_9780),
        .dout(new_Jinkela_wire_9781)
    );

    bfr new_Jinkela_buffer_2582 (
        .din(new_Jinkela_wire_2987),
        .dout(new_Jinkela_wire_2988)
    );

    bfr new_Jinkela_buffer_2527 (
        .din(new_Jinkela_wire_2928),
        .dout(new_Jinkela_wire_2929)
    );

    bfr new_Jinkela_buffer_263 (
        .din(new_Jinkela_wire_287),
        .dout(new_Jinkela_wire_288)
    );

    bfr new_Jinkela_buffer_7774 (
        .din(new_Jinkela_wire_9806),
        .dout(new_Jinkela_wire_9807)
    );

    bfr new_Jinkela_buffer_213 (
        .din(new_Jinkela_wire_232),
        .dout(new_Jinkela_wire_233)
    );

    bfr new_Jinkela_buffer_7749 (
        .din(new_Jinkela_wire_9781),
        .dout(new_Jinkela_wire_9782)
    );

    bfr new_Jinkela_buffer_2528 (
        .din(new_Jinkela_wire_2929),
        .dout(new_Jinkela_wire_2930)
    );

    bfr new_Jinkela_buffer_214 (
        .din(new_Jinkela_wire_233),
        .dout(new_Jinkela_wire_234)
    );

    bfr new_Jinkela_buffer_2583 (
        .din(new_Jinkela_wire_2988),
        .dout(new_Jinkela_wire_2989)
    );

    bfr new_Jinkela_buffer_7775 (
        .din(new_Jinkela_wire_9807),
        .dout(new_Jinkela_wire_9808)
    );

    bfr new_Jinkela_buffer_2529 (
        .din(new_Jinkela_wire_2930),
        .dout(new_Jinkela_wire_2931)
    );

    bfr new_Jinkela_buffer_264 (
        .din(new_Jinkela_wire_288),
        .dout(new_Jinkela_wire_289)
    );

    bfr new_Jinkela_buffer_7750 (
        .din(new_Jinkela_wire_9782),
        .dout(new_Jinkela_wire_9783)
    );

    bfr new_Jinkela_buffer_215 (
        .din(new_Jinkela_wire_234),
        .dout(new_Jinkela_wire_235)
    );

    bfr new_Jinkela_buffer_2775 (
        .din(N61),
        .dout(new_Jinkela_wire_3190)
    );

    spl2 new_Jinkela_splitter_818 (
        .a(n_0445_),
        .b(new_Jinkela_wire_9845),
        .c(new_Jinkela_wire_9846)
    );

    bfr new_Jinkela_buffer_2530 (
        .din(new_Jinkela_wire_2931),
        .dout(new_Jinkela_wire_2932)
    );

    spl2 new_Jinkela_splitter_12 (
        .a(new_Jinkela_wire_353),
        .b(new_Jinkela_wire_354),
        .c(new_Jinkela_wire_355)
    );

    bfr new_Jinkela_buffer_7751 (
        .din(new_Jinkela_wire_9783),
        .dout(new_Jinkela_wire_9784)
    );

    spl2 new_Jinkela_splitter_137 (
        .a(new_Jinkela_wire_3052),
        .b(new_Jinkela_wire_3053),
        .c(new_Jinkela_wire_3054)
    );

    bfr new_Jinkela_buffer_216 (
        .din(new_Jinkela_wire_235),
        .dout(new_Jinkela_wire_236)
    );

    spl2 new_Jinkela_splitter_815 (
        .a(new_Jinkela_wire_9833),
        .b(new_Jinkela_wire_9834),
        .c(new_Jinkela_wire_9835)
    );

    bfr new_Jinkela_buffer_2584 (
        .din(new_Jinkela_wire_2989),
        .dout(new_Jinkela_wire_2990)
    );

    bfr new_Jinkela_buffer_7776 (
        .din(new_Jinkela_wire_9808),
        .dout(new_Jinkela_wire_9809)
    );

    bfr new_Jinkela_buffer_2531 (
        .din(new_Jinkela_wire_2932),
        .dout(new_Jinkela_wire_2933)
    );

    bfr new_Jinkela_buffer_265 (
        .din(new_Jinkela_wire_289),
        .dout(new_Jinkela_wire_290)
    );

    bfr new_Jinkela_buffer_7752 (
        .din(new_Jinkela_wire_9784),
        .dout(new_Jinkela_wire_9785)
    );

    bfr new_Jinkela_buffer_217 (
        .din(new_Jinkela_wire_236),
        .dout(new_Jinkela_wire_237)
    );

    bfr new_Jinkela_buffer_2532 (
        .din(new_Jinkela_wire_2933),
        .dout(new_Jinkela_wire_2934)
    );

    bfr new_Jinkela_buffer_399 (
        .din(N219),
        .dout(new_Jinkela_wire_431)
    );

    bfr new_Jinkela_buffer_7753 (
        .din(new_Jinkela_wire_9785),
        .dout(new_Jinkela_wire_9786)
    );

    bfr new_Jinkela_buffer_331 (
        .din(new_Jinkela_wire_360),
        .dout(new_Jinkela_wire_361)
    );

    bfr new_Jinkela_buffer_2645 (
        .din(new_Jinkela_wire_3054),
        .dout(new_Jinkela_wire_3055)
    );

    bfr new_Jinkela_buffer_218 (
        .din(new_Jinkela_wire_237),
        .dout(new_Jinkela_wire_238)
    );

    bfr new_Jinkela_buffer_2585 (
        .din(new_Jinkela_wire_2990),
        .dout(new_Jinkela_wire_2991)
    );

    bfr new_Jinkela_buffer_7777 (
        .din(new_Jinkela_wire_9809),
        .dout(new_Jinkela_wire_9810)
    );

    bfr new_Jinkela_buffer_2533 (
        .din(new_Jinkela_wire_2934),
        .dout(new_Jinkela_wire_2935)
    );

    bfr new_Jinkela_buffer_266 (
        .din(new_Jinkela_wire_290),
        .dout(new_Jinkela_wire_291)
    );

    bfr new_Jinkela_buffer_7754 (
        .din(new_Jinkela_wire_9786),
        .dout(new_Jinkela_wire_9787)
    );

    bfr new_Jinkela_buffer_219 (
        .din(new_Jinkela_wire_238),
        .dout(new_Jinkela_wire_239)
    );

    spl2 new_Jinkela_splitter_819 (
        .a(n_0041_),
        .b(new_Jinkela_wire_9847),
        .c(new_Jinkela_wire_9848)
    );

    bfr new_Jinkela_buffer_2534 (
        .din(new_Jinkela_wire_2935),
        .dout(new_Jinkela_wire_2936)
    );

    bfr new_Jinkela_buffer_328 (
        .din(new_Jinkela_wire_357),
        .dout(new_Jinkela_wire_358)
    );

    bfr new_Jinkela_buffer_7755 (
        .din(new_Jinkela_wire_9787),
        .dout(new_Jinkela_wire_9788)
    );

    bfr new_Jinkela_buffer_2709 (
        .din(new_Jinkela_wire_3118),
        .dout(new_Jinkela_wire_3119)
    );

    bfr new_Jinkela_buffer_220 (
        .din(new_Jinkela_wire_239),
        .dout(new_Jinkela_wire_240)
    );

    bfr new_Jinkela_buffer_7802 (
        .din(new_Jinkela_wire_9836),
        .dout(new_Jinkela_wire_9837)
    );

    bfr new_Jinkela_buffer_2586 (
        .din(new_Jinkela_wire_2991),
        .dout(new_Jinkela_wire_2992)
    );

    bfr new_Jinkela_buffer_7778 (
        .din(new_Jinkela_wire_9810),
        .dout(new_Jinkela_wire_9811)
    );

    bfr new_Jinkela_buffer_1750 (
        .din(new_Jinkela_wire_2100),
        .dout(new_Jinkela_wire_2101)
    );

    bfr new_Jinkela_buffer_3371 (
        .din(new_Jinkela_wire_3905),
        .dout(new_Jinkela_wire_3906)
    );

    bfr new_Jinkela_buffer_1704 (
        .din(new_Jinkela_wire_2049),
        .dout(new_Jinkela_wire_2050)
    );

    bfr new_Jinkela_buffer_6699 (
        .din(new_Jinkela_wire_8220),
        .dout(new_Jinkela_wire_8221)
    );

    spl2 new_Jinkela_splitter_204 (
        .a(n_0721_),
        .b(new_Jinkela_wire_4045),
        .c(new_Jinkela_wire_4046)
    );

    bfr new_Jinkela_buffer_1882 (
        .din(N310),
        .dout(new_Jinkela_wire_2237)
    );

    bfr new_Jinkela_buffer_3372 (
        .din(new_Jinkela_wire_3906),
        .dout(new_Jinkela_wire_3907)
    );

    bfr new_Jinkela_buffer_6747 (
        .din(new_Jinkela_wire_8304),
        .dout(new_Jinkela_wire_8305)
    );

    bfr new_Jinkela_buffer_1705 (
        .din(new_Jinkela_wire_2050),
        .dout(new_Jinkela_wire_2051)
    );

    bfr new_Jinkela_buffer_6700 (
        .din(new_Jinkela_wire_8221),
        .dout(new_Jinkela_wire_8222)
    );

    bfr new_Jinkela_buffer_3393 (
        .din(new_Jinkela_wire_3954),
        .dout(new_Jinkela_wire_3955)
    );

    bfr new_Jinkela_buffer_1945 (
        .din(new_Jinkela_wire_2307),
        .dout(new_Jinkela_wire_2308)
    );

    spl2 new_Jinkela_splitter_202 (
        .a(n_0294_),
        .b(new_Jinkela_wire_4014),
        .c(new_Jinkela_wire_4015)
    );

    bfr new_Jinkela_buffer_1751 (
        .din(new_Jinkela_wire_2101),
        .dout(new_Jinkela_wire_2102)
    );

    bfr new_Jinkela_buffer_3373 (
        .din(new_Jinkela_wire_3907),
        .dout(new_Jinkela_wire_3908)
    );

    bfr new_Jinkela_buffer_6755 (
        .din(n_0330_),
        .dout(new_Jinkela_wire_8322)
    );

    bfr new_Jinkela_buffer_1706 (
        .din(new_Jinkela_wire_2051),
        .dout(new_Jinkela_wire_2052)
    );

    bfr new_Jinkela_buffer_6701 (
        .din(new_Jinkela_wire_8222),
        .dout(new_Jinkela_wire_8223)
    );

    bfr new_Jinkela_buffer_1879 (
        .din(new_Jinkela_wire_2233),
        .dout(new_Jinkela_wire_2234)
    );

    bfr new_Jinkela_buffer_3374 (
        .din(new_Jinkela_wire_3908),
        .dout(new_Jinkela_wire_3909)
    );

    bfr new_Jinkela_buffer_6748 (
        .din(new_Jinkela_wire_8305),
        .dout(new_Jinkela_wire_8306)
    );

    bfr new_Jinkela_buffer_1707 (
        .din(new_Jinkela_wire_2052),
        .dout(new_Jinkela_wire_2053)
    );

    bfr new_Jinkela_buffer_6702 (
        .din(new_Jinkela_wire_8223),
        .dout(new_Jinkela_wire_8224)
    );

    bfr new_Jinkela_buffer_3394 (
        .din(new_Jinkela_wire_3955),
        .dout(new_Jinkela_wire_3956)
    );

    bfr new_Jinkela_buffer_1752 (
        .din(new_Jinkela_wire_2102),
        .dout(new_Jinkela_wire_2103)
    );

    bfr new_Jinkela_buffer_3375 (
        .din(new_Jinkela_wire_3909),
        .dout(new_Jinkela_wire_3910)
    );

    bfr new_Jinkela_buffer_6753 (
        .din(n_1096_),
        .dout(new_Jinkela_wire_8315)
    );

    bfr new_Jinkela_buffer_1708 (
        .din(new_Jinkela_wire_2053),
        .dout(new_Jinkela_wire_2054)
    );

    bfr new_Jinkela_buffer_6703 (
        .din(new_Jinkela_wire_8224),
        .dout(new_Jinkela_wire_8225)
    );

    bfr new_Jinkela_buffer_3445 (
        .din(n_0082_),
        .dout(new_Jinkela_wire_4016)
    );

    bfr new_Jinkela_buffer_6750 (
        .din(new_Jinkela_wire_8309),
        .dout(new_Jinkela_wire_8310)
    );

    bfr new_Jinkela_buffer_1815 (
        .din(new_Jinkela_wire_2167),
        .dout(new_Jinkela_wire_2168)
    );

    bfr new_Jinkela_buffer_3395 (
        .din(new_Jinkela_wire_3956),
        .dout(new_Jinkela_wire_3957)
    );

    bfr new_Jinkela_buffer_1709 (
        .din(new_Jinkela_wire_2054),
        .dout(new_Jinkela_wire_2055)
    );

    bfr new_Jinkela_buffer_6704 (
        .din(new_Jinkela_wire_8225),
        .dout(new_Jinkela_wire_8226)
    );

    bfr new_Jinkela_buffer_3472 (
        .din(new_Jinkela_wire_4046),
        .dout(new_Jinkela_wire_4047)
    );

    spl2 new_Jinkela_splitter_625 (
        .a(n_0523_),
        .b(new_Jinkela_wire_8325),
        .c(new_Jinkela_wire_8326)
    );

    bfr new_Jinkela_buffer_1753 (
        .din(new_Jinkela_wire_2103),
        .dout(new_Jinkela_wire_2104)
    );

    bfr new_Jinkela_buffer_3396 (
        .din(new_Jinkela_wire_3957),
        .dout(new_Jinkela_wire_3958)
    );

    bfr new_Jinkela_buffer_6751 (
        .din(new_Jinkela_wire_8310),
        .dout(new_Jinkela_wire_8311)
    );

    bfr new_Jinkela_buffer_1710 (
        .din(new_Jinkela_wire_2055),
        .dout(new_Jinkela_wire_2056)
    );

    bfr new_Jinkela_buffer_6705 (
        .din(new_Jinkela_wire_8226),
        .dout(new_Jinkela_wire_8227)
    );

    spl2 new_Jinkela_splitter_200 (
        .a(new_Jinkela_wire_4009),
        .b(new_Jinkela_wire_4010),
        .c(new_Jinkela_wire_4011)
    );

    bfr new_Jinkela_buffer_3474 (
        .din(n_0343_),
        .dout(new_Jinkela_wire_4049)
    );

    spl2 new_Jinkela_splitter_117 (
        .a(N355),
        .b(new_Jinkela_wire_2306),
        .c(new_Jinkela_wire_2307)
    );

    bfr new_Jinkela_buffer_3397 (
        .din(new_Jinkela_wire_3958),
        .dout(new_Jinkela_wire_3959)
    );

    bfr new_Jinkela_buffer_1711 (
        .din(new_Jinkela_wire_2056),
        .dout(new_Jinkela_wire_2057)
    );

    bfr new_Jinkela_buffer_6706 (
        .din(new_Jinkela_wire_8227),
        .dout(new_Jinkela_wire_8228)
    );

    bfr new_Jinkela_buffer_1754 (
        .din(new_Jinkela_wire_2104),
        .dout(new_Jinkela_wire_2105)
    );

    bfr new_Jinkela_buffer_3398 (
        .din(new_Jinkela_wire_3959),
        .dout(new_Jinkela_wire_3960)
    );

    bfr new_Jinkela_buffer_1712 (
        .din(new_Jinkela_wire_2057),
        .dout(new_Jinkela_wire_2058)
    );

    bfr new_Jinkela_buffer_6707 (
        .din(new_Jinkela_wire_8228),
        .dout(new_Jinkela_wire_8229)
    );

    bfr new_Jinkela_buffer_3446 (
        .din(new_Jinkela_wire_4016),
        .dout(new_Jinkela_wire_4017)
    );

    bfr new_Jinkela_buffer_6752 (
        .din(new_Jinkela_wire_8311),
        .dout(new_Jinkela_wire_8312)
    );

    spl2 new_Jinkela_splitter_113 (
        .a(new_Jinkela_wire_2168),
        .b(new_Jinkela_wire_2169),
        .c(new_Jinkela_wire_2170)
    );

    bfr new_Jinkela_buffer_3399 (
        .din(new_Jinkela_wire_3960),
        .dout(new_Jinkela_wire_3961)
    );

    bfr new_Jinkela_buffer_1713 (
        .din(new_Jinkela_wire_2058),
        .dout(new_Jinkela_wire_2059)
    );

    bfr new_Jinkela_buffer_6708 (
        .din(new_Jinkela_wire_8229),
        .dout(new_Jinkela_wire_8230)
    );

    spl3L new_Jinkela_splitter_622 (
        .a(new_Jinkela_wire_8315),
        .d(new_Jinkela_wire_8316),
        .b(new_Jinkela_wire_8317),
        .c(new_Jinkela_wire_8318)
    );

    bfr new_Jinkela_buffer_1755 (
        .din(new_Jinkela_wire_2105),
        .dout(new_Jinkela_wire_2106)
    );

    bfr new_Jinkela_buffer_3400 (
        .din(new_Jinkela_wire_3961),
        .dout(new_Jinkela_wire_3962)
    );

    bfr new_Jinkela_buffer_1714 (
        .din(new_Jinkela_wire_2059),
        .dout(new_Jinkela_wire_2060)
    );

    bfr new_Jinkela_buffer_6709 (
        .din(new_Jinkela_wire_8230),
        .dout(new_Jinkela_wire_8231)
    );

    spl2 new_Jinkela_splitter_203 (
        .a(new_Jinkela_wire_4017),
        .b(new_Jinkela_wire_4018),
        .c(new_Jinkela_wire_4019)
    );

    spl2 new_Jinkela_splitter_621 (
        .a(new_Jinkela_wire_8312),
        .b(new_Jinkela_wire_8313),
        .c(new_Jinkela_wire_8314)
    );

    bfr new_Jinkela_buffer_1816 (
        .din(new_Jinkela_wire_2170),
        .dout(new_Jinkela_wire_2171)
    );

    bfr new_Jinkela_buffer_3401 (
        .din(new_Jinkela_wire_3962),
        .dout(new_Jinkela_wire_3963)
    );

    bfr new_Jinkela_buffer_1715 (
        .din(new_Jinkela_wire_2060),
        .dout(new_Jinkela_wire_2061)
    );

    bfr new_Jinkela_buffer_6710 (
        .din(new_Jinkela_wire_8231),
        .dout(new_Jinkela_wire_8232)
    );

    bfr new_Jinkela_buffer_3447 (
        .din(new_Jinkela_wire_4019),
        .dout(new_Jinkela_wire_4020)
    );

    spl2 new_Jinkela_splitter_624 (
        .a(n_1271_),
        .b(new_Jinkela_wire_8323),
        .c(new_Jinkela_wire_8324)
    );

    bfr new_Jinkela_buffer_1756 (
        .din(new_Jinkela_wire_2106),
        .dout(new_Jinkela_wire_2107)
    );

    bfr new_Jinkela_buffer_3402 (
        .din(new_Jinkela_wire_3963),
        .dout(new_Jinkela_wire_3964)
    );

    bfr new_Jinkela_buffer_1716 (
        .din(new_Jinkela_wire_2061),
        .dout(new_Jinkela_wire_2062)
    );

    bfr new_Jinkela_buffer_6711 (
        .din(new_Jinkela_wire_8232),
        .dout(new_Jinkela_wire_8233)
    );

    bfr new_Jinkela_buffer_3491 (
        .din(n_0454_),
        .dout(new_Jinkela_wire_4070)
    );

    bfr new_Jinkela_buffer_6754 (
        .din(new_Jinkela_wire_8318),
        .dout(new_Jinkela_wire_8319)
    );

    bfr new_Jinkela_buffer_1880 (
        .din(new_Jinkela_wire_2234),
        .dout(new_Jinkela_wire_2235)
    );

    bfr new_Jinkela_buffer_3403 (
        .din(new_Jinkela_wire_3964),
        .dout(new_Jinkela_wire_3965)
    );

    bfr new_Jinkela_buffer_1717 (
        .din(new_Jinkela_wire_2062),
        .dout(new_Jinkela_wire_2063)
    );

    bfr new_Jinkela_buffer_6712 (
        .din(new_Jinkela_wire_8233),
        .dout(new_Jinkela_wire_8234)
    );

    spl2 new_Jinkela_splitter_208 (
        .a(n_0650_),
        .b(new_Jinkela_wire_4078),
        .c(new_Jinkela_wire_4079)
    );

    spl2 new_Jinkela_splitter_626 (
        .a(n_0859_),
        .b(new_Jinkela_wire_8327),
        .c(new_Jinkela_wire_8328)
    );

    bfr new_Jinkela_buffer_1757 (
        .din(new_Jinkela_wire_2107),
        .dout(new_Jinkela_wire_2108)
    );

    bfr new_Jinkela_buffer_3404 (
        .din(new_Jinkela_wire_3965),
        .dout(new_Jinkela_wire_3966)
    );

    spl2 new_Jinkela_splitter_623 (
        .a(new_Jinkela_wire_8319),
        .b(new_Jinkela_wire_8320),
        .c(new_Jinkela_wire_8321)
    );

    bfr new_Jinkela_buffer_1718 (
        .din(new_Jinkela_wire_2063),
        .dout(new_Jinkela_wire_2064)
    );

    bfr new_Jinkela_buffer_6713 (
        .din(new_Jinkela_wire_8234),
        .dout(new_Jinkela_wire_8235)
    );

    spl2 new_Jinkela_splitter_205 (
        .a(new_Jinkela_wire_4049),
        .b(new_Jinkela_wire_4050),
        .c(new_Jinkela_wire_4051)
    );

    bfr new_Jinkela_buffer_3448 (
        .din(new_Jinkela_wire_4020),
        .dout(new_Jinkela_wire_4021)
    );

    bfr new_Jinkela_buffer_2009 (
        .din(N173),
        .dout(new_Jinkela_wire_2374)
    );

    bfr new_Jinkela_buffer_3405 (
        .din(new_Jinkela_wire_3966),
        .dout(new_Jinkela_wire_3967)
    );

    bfr new_Jinkela_buffer_6714 (
        .din(new_Jinkela_wire_8235),
        .dout(new_Jinkela_wire_8236)
    );

    bfr new_Jinkela_buffer_1758 (
        .din(new_Jinkela_wire_2108),
        .dout(new_Jinkela_wire_2109)
    );

    bfr new_Jinkela_buffer_3473 (
        .din(new_Jinkela_wire_4047),
        .dout(new_Jinkela_wire_4048)
    );

    bfr new_Jinkela_buffer_1817 (
        .din(new_Jinkela_wire_2171),
        .dout(new_Jinkela_wire_2172)
    );

    bfr new_Jinkela_buffer_3406 (
        .din(new_Jinkela_wire_3967),
        .dout(new_Jinkela_wire_3968)
    );

    bfr new_Jinkela_buffer_6782 (
        .din(n_0240_),
        .dout(new_Jinkela_wire_8358)
    );

    bfr new_Jinkela_buffer_6715 (
        .din(new_Jinkela_wire_8236),
        .dout(new_Jinkela_wire_8237)
    );

    bfr new_Jinkela_buffer_1759 (
        .din(new_Jinkela_wire_2109),
        .dout(new_Jinkela_wire_2110)
    );

    bfr new_Jinkela_buffer_3449 (
        .din(new_Jinkela_wire_4021),
        .dout(new_Jinkela_wire_4022)
    );

    bfr new_Jinkela_buffer_6756 (
        .din(n_0390_),
        .dout(new_Jinkela_wire_8329)
    );

    bfr new_Jinkela_buffer_1881 (
        .din(new_Jinkela_wire_2235),
        .dout(new_Jinkela_wire_2236)
    );

    bfr new_Jinkela_buffer_3407 (
        .din(new_Jinkela_wire_3968),
        .dout(new_Jinkela_wire_3969)
    );

    bfr new_Jinkela_buffer_6781 (
        .din(n_0077_),
        .dout(new_Jinkela_wire_8357)
    );

    bfr new_Jinkela_buffer_6716 (
        .din(new_Jinkela_wire_8237),
        .dout(new_Jinkela_wire_8238)
    );

    bfr new_Jinkela_buffer_1760 (
        .din(new_Jinkela_wire_2110),
        .dout(new_Jinkela_wire_2111)
    );

    spl2 new_Jinkela_splitter_209 (
        .a(n_1322_),
        .b(new_Jinkela_wire_4080),
        .c(new_Jinkela_wire_4081)
    );

    bfr new_Jinkela_buffer_1818 (
        .din(new_Jinkela_wire_2172),
        .dout(new_Jinkela_wire_2173)
    );

    bfr new_Jinkela_buffer_3408 (
        .din(new_Jinkela_wire_3969),
        .dout(new_Jinkela_wire_3970)
    );

    bfr new_Jinkela_buffer_6757 (
        .din(new_Jinkela_wire_8329),
        .dout(new_Jinkela_wire_8330)
    );

    bfr new_Jinkela_buffer_6717 (
        .din(new_Jinkela_wire_8238),
        .dout(new_Jinkela_wire_8239)
    );

    bfr new_Jinkela_buffer_1761 (
        .din(new_Jinkela_wire_2111),
        .dout(new_Jinkela_wire_2112)
    );

    bfr new_Jinkela_buffer_3450 (
        .din(new_Jinkela_wire_4022),
        .dout(new_Jinkela_wire_4023)
    );

    bfr new_Jinkela_buffer_6758 (
        .din(new_Jinkela_wire_8330),
        .dout(new_Jinkela_wire_8331)
    );

    bfr new_Jinkela_buffer_3409 (
        .din(new_Jinkela_wire_3970),
        .dout(new_Jinkela_wire_3971)
    );

    bfr new_Jinkela_buffer_1883 (
        .din(new_Jinkela_wire_2237),
        .dout(new_Jinkela_wire_2238)
    );

    bfr new_Jinkela_buffer_6718 (
        .din(new_Jinkela_wire_8239),
        .dout(new_Jinkela_wire_8240)
    );

    bfr new_Jinkela_buffer_1762 (
        .din(new_Jinkela_wire_2112),
        .dout(new_Jinkela_wire_2113)
    );

    bfr new_Jinkela_buffer_1819 (
        .din(new_Jinkela_wire_2173),
        .dout(new_Jinkela_wire_2174)
    );

    bfr new_Jinkela_buffer_3410 (
        .din(new_Jinkela_wire_3971),
        .dout(new_Jinkela_wire_3972)
    );

    bfr new_Jinkela_buffer_6719 (
        .din(new_Jinkela_wire_8240),
        .dout(new_Jinkela_wire_8241)
    );

    bfr new_Jinkela_buffer_1763 (
        .din(new_Jinkela_wire_2113),
        .dout(new_Jinkela_wire_2114)
    );

    bfr new_Jinkela_buffer_3475 (
        .din(new_Jinkela_wire_4051),
        .dout(new_Jinkela_wire_4052)
    );

    bfr new_Jinkela_buffer_3451 (
        .din(new_Jinkela_wire_4023),
        .dout(new_Jinkela_wire_4024)
    );

    bfr new_Jinkela_buffer_6785 (
        .din(n_0737_),
        .dout(new_Jinkela_wire_8361)
    );

    bfr new_Jinkela_buffer_5899 (
        .din(new_Jinkela_wire_7138),
        .dout(new_Jinkela_wire_7139)
    );

    bfr new_Jinkela_buffer_5969 (
        .din(new_Jinkela_wire_7217),
        .dout(new_Jinkela_wire_7218)
    );

    bfr new_Jinkela_buffer_5900 (
        .din(new_Jinkela_wire_7139),
        .dout(new_Jinkela_wire_7140)
    );

    bfr new_Jinkela_buffer_5955 (
        .din(new_Jinkela_wire_7196),
        .dout(new_Jinkela_wire_7197)
    );

    bfr new_Jinkela_buffer_5901 (
        .din(new_Jinkela_wire_7140),
        .dout(new_Jinkela_wire_7141)
    );

    bfr new_Jinkela_buffer_5960 (
        .din(new_Jinkela_wire_7208),
        .dout(new_Jinkela_wire_7209)
    );

    bfr new_Jinkela_buffer_5902 (
        .din(new_Jinkela_wire_7141),
        .dout(new_Jinkela_wire_7142)
    );

    bfr new_Jinkela_buffer_5956 (
        .din(new_Jinkela_wire_7197),
        .dout(new_Jinkela_wire_7198)
    );

    bfr new_Jinkela_buffer_5903 (
        .din(new_Jinkela_wire_7142),
        .dout(new_Jinkela_wire_7143)
    );

    spl2 new_Jinkela_splitter_491 (
        .a(n_0054_),
        .b(new_Jinkela_wire_7234),
        .c(new_Jinkela_wire_7235)
    );

    bfr new_Jinkela_buffer_5904 (
        .din(new_Jinkela_wire_7143),
        .dout(new_Jinkela_wire_7144)
    );

    bfr new_Jinkela_buffer_5957 (
        .din(new_Jinkela_wire_7198),
        .dout(new_Jinkela_wire_7199)
    );

    bfr new_Jinkela_buffer_5905 (
        .din(new_Jinkela_wire_7144),
        .dout(new_Jinkela_wire_7145)
    );

    bfr new_Jinkela_buffer_5961 (
        .din(new_Jinkela_wire_7209),
        .dout(new_Jinkela_wire_7210)
    );

    bfr new_Jinkela_buffer_5906 (
        .din(new_Jinkela_wire_7145),
        .dout(new_Jinkela_wire_7146)
    );

    bfr new_Jinkela_buffer_5970 (
        .din(new_Jinkela_wire_7218),
        .dout(new_Jinkela_wire_7219)
    );

    bfr new_Jinkela_buffer_5907 (
        .din(new_Jinkela_wire_7146),
        .dout(new_Jinkela_wire_7147)
    );

    bfr new_Jinkela_buffer_5962 (
        .din(new_Jinkela_wire_7210),
        .dout(new_Jinkela_wire_7211)
    );

    bfr new_Jinkela_buffer_5908 (
        .din(new_Jinkela_wire_7147),
        .dout(new_Jinkela_wire_7148)
    );

    spl2 new_Jinkela_splitter_489 (
        .a(new_Jinkela_wire_7224),
        .b(new_Jinkela_wire_7225),
        .c(new_Jinkela_wire_7226)
    );

    bfr new_Jinkela_buffer_5909 (
        .din(new_Jinkela_wire_7148),
        .dout(new_Jinkela_wire_7149)
    );

    bfr new_Jinkela_buffer_5963 (
        .din(new_Jinkela_wire_7211),
        .dout(new_Jinkela_wire_7212)
    );

    bfr new_Jinkela_buffer_5910 (
        .din(new_Jinkela_wire_7149),
        .dout(new_Jinkela_wire_7150)
    );

    bfr new_Jinkela_buffer_5971 (
        .din(new_Jinkela_wire_7219),
        .dout(new_Jinkela_wire_7220)
    );

    bfr new_Jinkela_buffer_5911 (
        .din(new_Jinkela_wire_7150),
        .dout(new_Jinkela_wire_7151)
    );

    bfr new_Jinkela_buffer_5964 (
        .din(new_Jinkela_wire_7212),
        .dout(new_Jinkela_wire_7213)
    );

    bfr new_Jinkela_buffer_5912 (
        .din(new_Jinkela_wire_7151),
        .dout(new_Jinkela_wire_7152)
    );

    bfr new_Jinkela_buffer_5975 (
        .din(new_Jinkela_wire_7227),
        .dout(new_Jinkela_wire_7228)
    );

    bfr new_Jinkela_buffer_5913 (
        .din(new_Jinkela_wire_7152),
        .dout(new_Jinkela_wire_7153)
    );

    bfr new_Jinkela_buffer_5965 (
        .din(new_Jinkela_wire_7213),
        .dout(new_Jinkela_wire_7214)
    );

    bfr new_Jinkela_buffer_5914 (
        .din(new_Jinkela_wire_7153),
        .dout(new_Jinkela_wire_7154)
    );

    bfr new_Jinkela_buffer_5972 (
        .din(new_Jinkela_wire_7220),
        .dout(new_Jinkela_wire_7221)
    );

    bfr new_Jinkela_buffer_5915 (
        .din(new_Jinkela_wire_7154),
        .dout(new_Jinkela_wire_7155)
    );

    bfr new_Jinkela_buffer_5966 (
        .din(new_Jinkela_wire_7214),
        .dout(new_Jinkela_wire_7215)
    );

    bfr new_Jinkela_buffer_5916 (
        .din(new_Jinkela_wire_7155),
        .dout(new_Jinkela_wire_7156)
    );

    bfr new_Jinkela_buffer_5979 (
        .din(n_0821_),
        .dout(new_Jinkela_wire_7236)
    );

    bfr new_Jinkela_buffer_5917 (
        .din(new_Jinkela_wire_7156),
        .dout(new_Jinkela_wire_7157)
    );

    bfr new_Jinkela_buffer_5982 (
        .din(n_0936_),
        .dout(new_Jinkela_wire_7241)
    );

    bfr new_Jinkela_buffer_5967 (
        .din(new_Jinkela_wire_7215),
        .dout(new_Jinkela_wire_7216)
    );

    bfr new_Jinkela_buffer_5918 (
        .din(new_Jinkela_wire_7157),
        .dout(new_Jinkela_wire_7158)
    );

    spl2 new_Jinkela_splitter_488 (
        .a(new_Jinkela_wire_7221),
        .b(new_Jinkela_wire_7222),
        .c(new_Jinkela_wire_7223)
    );

    bfr new_Jinkela_buffer_5919 (
        .din(new_Jinkela_wire_7158),
        .dout(new_Jinkela_wire_7159)
    );

    and_bi n_2664_ (
        .a(new_Jinkela_wire_4088),
        .b(new_Jinkela_wire_5166),
        .c(n_0521_)
    );

    bfr new_Jinkela_buffer_5098 (
        .din(new_Jinkela_wire_6075),
        .dout(new_Jinkela_wire_6076)
    );

    and_ii n_1947_ (
        .a(new_Jinkela_wire_7330),
        .b(new_Jinkela_wire_9447),
        .c(n_1213_)
    );

    bfr new_Jinkela_buffer_5072 (
        .din(new_Jinkela_wire_6047),
        .dout(new_Jinkela_wire_6048)
    );

    bfr new_Jinkela_buffer_6720 (
        .din(new_Jinkela_wire_8241),
        .dout(new_Jinkela_wire_8242)
    );

    and_bi n_2665_ (
        .a(new_Jinkela_wire_5167),
        .b(new_Jinkela_wire_4089),
        .c(n_0522_)
    );

    bfr new_Jinkela_buffer_6783 (
        .din(new_Jinkela_wire_8358),
        .dout(new_Jinkela_wire_8359)
    );

    and_bi n_1948_ (
        .a(new_Jinkela_wire_1358),
        .b(new_Jinkela_wire_191),
        .c(n_1214_)
    );

    spl3L new_Jinkela_splitter_627 (
        .a(new_Jinkela_wire_8331),
        .d(new_Jinkela_wire_8332),
        .b(new_Jinkela_wire_8333),
        .c(new_Jinkela_wire_8334)
    );

    and_ii n_2666_ (
        .a(n_0522_),
        .b(n_0521_),
        .c(n_0523_)
    );

    and_bb n_1949_ (
        .a(new_Jinkela_wire_5105),
        .b(new_Jinkela_wire_10563),
        .c(n_1215_)
    );

    bfr new_Jinkela_buffer_5073 (
        .din(new_Jinkela_wire_6048),
        .dout(new_Jinkela_wire_6049)
    );

    bfr new_Jinkela_buffer_6721 (
        .din(new_Jinkela_wire_8242),
        .dout(new_Jinkela_wire_8243)
    );

    and_bb n_2667_ (
        .a(new_Jinkela_wire_8326),
        .b(new_Jinkela_wire_7413),
        .c(n_0524_)
    );

    and_ii n_1950_ (
        .a(new_Jinkela_wire_5102),
        .b(new_Jinkela_wire_9459),
        .c(n_1216_)
    );

    and_ii n_2668_ (
        .a(new_Jinkela_wire_8325),
        .b(new_Jinkela_wire_7412),
        .c(n_0525_)
    );

    bfr new_Jinkela_buffer_5099 (
        .din(new_Jinkela_wire_6076),
        .dout(new_Jinkela_wire_6077)
    );

    and_bb n_1951_ (
        .a(new_Jinkela_wire_4087),
        .b(new_Jinkela_wire_7333),
        .c(n_1217_)
    );

    bfr new_Jinkela_buffer_5074 (
        .din(new_Jinkela_wire_6049),
        .dout(new_Jinkela_wire_6050)
    );

    bfr new_Jinkela_buffer_6722 (
        .din(new_Jinkela_wire_8243),
        .dout(new_Jinkela_wire_8244)
    );

    and_ii n_2669_ (
        .a(n_0525_),
        .b(n_0524_),
        .c(n_0526_)
    );

    spl4L new_Jinkela_splitter_628 (
        .a(n_0662_),
        .d(new_Jinkela_wire_8362),
        .b(new_Jinkela_wire_8363),
        .e(new_Jinkela_wire_8364),
        .c(new_Jinkela_wire_8365)
    );

    and_ii n_1952_ (
        .a(n_1217_),
        .b(n_1215_),
        .c(n_1218_)
    );

    bfr new_Jinkela_buffer_6759 (
        .din(new_Jinkela_wire_8334),
        .dout(new_Jinkela_wire_8335)
    );

    or_bb n_2670_ (
        .a(new_Jinkela_wire_7013),
        .b(new_Jinkela_wire_9893),
        .c(n_0527_)
    );

    and_bb n_1953_ (
        .a(new_Jinkela_wire_8103),
        .b(new_Jinkela_wire_4507),
        .c(n_1219_)
    );

    bfr new_Jinkela_buffer_5075 (
        .din(new_Jinkela_wire_6050),
        .dout(new_Jinkela_wire_6051)
    );

    bfr new_Jinkela_buffer_6723 (
        .din(new_Jinkela_wire_8244),
        .dout(new_Jinkela_wire_8245)
    );

    and_bb n_2671_ (
        .a(new_Jinkela_wire_7012),
        .b(new_Jinkela_wire_9894),
        .c(n_0528_)
    );

    and_ii n_1954_ (
        .a(new_Jinkela_wire_8102),
        .b(new_Jinkela_wire_4506),
        .c(n_1220_)
    );

    bfr new_Jinkela_buffer_5116 (
        .din(new_Jinkela_wire_6095),
        .dout(new_Jinkela_wire_6096)
    );

    spl2 new_Jinkela_splitter_629 (
        .a(n_0327_),
        .b(new_Jinkela_wire_8366),
        .c(new_Jinkela_wire_8367)
    );

    and_bi n_2672_ (
        .a(n_0527_),
        .b(n_0528_),
        .c(n_0529_)
    );

    bfr new_Jinkela_buffer_5100 (
        .din(new_Jinkela_wire_6077),
        .dout(new_Jinkela_wire_6078)
    );

    or_bb n_1955_ (
        .a(n_1220_),
        .b(n_1219_),
        .c(n_1221_)
    );

    bfr new_Jinkela_buffer_5076 (
        .din(new_Jinkela_wire_6051),
        .dout(new_Jinkela_wire_6052)
    );

    bfr new_Jinkela_buffer_6724 (
        .din(new_Jinkela_wire_8245),
        .dout(new_Jinkela_wire_8246)
    );

    and_bi n_2673_ (
        .a(new_Jinkela_wire_9418),
        .b(new_Jinkela_wire_8867),
        .c(n_0530_)
    );

    and_ii n_1956_ (
        .a(new_Jinkela_wire_8438),
        .b(new_Jinkela_wire_3948),
        .c(n_1222_)
    );

    bfr new_Jinkela_buffer_6760 (
        .din(new_Jinkela_wire_8335),
        .dout(new_Jinkela_wire_8336)
    );

    and_bi n_2674_ (
        .a(new_Jinkela_wire_6532),
        .b(new_Jinkela_wire_10527),
        .c(n_0531_)
    );

    and_bb n_1957_ (
        .a(new_Jinkela_wire_8437),
        .b(new_Jinkela_wire_3947),
        .c(n_1223_)
    );

    bfr new_Jinkela_buffer_5077 (
        .din(new_Jinkela_wire_6052),
        .dout(new_Jinkela_wire_6053)
    );

    bfr new_Jinkela_buffer_6725 (
        .din(new_Jinkela_wire_8246),
        .dout(new_Jinkela_wire_8247)
    );

    and_bi n_2675_ (
        .a(new_Jinkela_wire_3877),
        .b(n_0531_),
        .c(n_0532_)
    );

    and_ii n_1958_ (
        .a(n_1223_),
        .b(n_1222_),
        .c(n_1224_)
    );

    spl2 new_Jinkela_splitter_383 (
        .a(n_0560_),
        .b(new_Jinkela_wire_6132),
        .c(new_Jinkela_wire_6133)
    );

    and_bi n_2676_ (
        .a(new_Jinkela_wire_8332),
        .b(new_Jinkela_wire_4644),
        .c(n_0533_)
    );

    bfr new_Jinkela_buffer_5101 (
        .din(new_Jinkela_wire_6078),
        .dout(new_Jinkela_wire_6079)
    );

    and_bb n_1959_ (
        .a(new_Jinkela_wire_2470),
        .b(new_Jinkela_wire_1289),
        .c(n_1225_)
    );

    bfr new_Jinkela_buffer_5078 (
        .din(new_Jinkela_wire_6053),
        .dout(new_Jinkela_wire_6054)
    );

    bfr new_Jinkela_buffer_6726 (
        .din(new_Jinkela_wire_8247),
        .dout(new_Jinkela_wire_8248)
    );

    and_bi n_2677_ (
        .a(new_Jinkela_wire_4643),
        .b(new_Jinkela_wire_8333),
        .c(n_0534_)
    );

    and_ii n_1960_ (
        .a(new_Jinkela_wire_9955),
        .b(new_Jinkela_wire_8279),
        .c(n_1226_)
    );

    bfr new_Jinkela_buffer_6761 (
        .din(new_Jinkela_wire_8336),
        .dout(new_Jinkela_wire_8337)
    );

    or_bb n_2678_ (
        .a(n_0534_),
        .b(n_0533_),
        .c(n_0535_)
    );

    and_bi n_1961_ (
        .a(new_Jinkela_wire_1218),
        .b(new_Jinkela_wire_2816),
        .c(n_1227_)
    );

    bfr new_Jinkela_buffer_5079 (
        .din(new_Jinkela_wire_6054),
        .dout(new_Jinkela_wire_6055)
    );

    bfr new_Jinkela_buffer_6727 (
        .din(new_Jinkela_wire_8248),
        .dout(new_Jinkela_wire_8249)
    );

    and_bi n_2679_ (
        .a(new_Jinkela_wire_10529),
        .b(new_Jinkela_wire_9779),
        .c(n_0536_)
    );

    and_ii n_1962_ (
        .a(n_1227_),
        .b(new_Jinkela_wire_9438),
        .c(n_1228_)
    );

    bfr new_Jinkela_buffer_5119 (
        .din(new_Jinkela_wire_6110),
        .dout(new_Jinkela_wire_6111)
    );

    spl2 new_Jinkela_splitter_630 (
        .a(n_0429_),
        .b(new_Jinkela_wire_8369),
        .c(new_Jinkela_wire_8370)
    );

    and_bi n_2680_ (
        .a(new_Jinkela_wire_9772),
        .b(new_Jinkela_wire_3780),
        .c(n_0537_)
    );

    bfr new_Jinkela_buffer_5102 (
        .din(new_Jinkela_wire_6079),
        .dout(new_Jinkela_wire_6080)
    );

    and_ii n_1963_ (
        .a(new_Jinkela_wire_6109),
        .b(new_Jinkela_wire_7328),
        .c(n_1229_)
    );

    bfr new_Jinkela_buffer_5080 (
        .din(new_Jinkela_wire_6055),
        .dout(new_Jinkela_wire_6056)
    );

    bfr new_Jinkela_buffer_6728 (
        .din(new_Jinkela_wire_8249),
        .dout(new_Jinkela_wire_8250)
    );

    and_ii n_2681_ (
        .a(new_Jinkela_wire_9479),
        .b(n_0536_),
        .c(n_0538_)
    );

    bfr new_Jinkela_buffer_6787 (
        .din(n_0421_),
        .dout(new_Jinkela_wire_8371)
    );

    and_bb n_1964_ (
        .a(new_Jinkela_wire_6108),
        .b(new_Jinkela_wire_7326),
        .c(n_1230_)
    );

    bfr new_Jinkela_buffer_6762 (
        .din(new_Jinkela_wire_8337),
        .dout(new_Jinkela_wire_8338)
    );

    and_bi n_2682_ (
        .a(new_Jinkela_wire_8164),
        .b(new_Jinkela_wire_4096),
        .c(n_0539_)
    );

    spl2 new_Jinkela_splitter_384 (
        .a(n_1355_),
        .b(new_Jinkela_wire_6134),
        .c(new_Jinkela_wire_6136)
    );

    and_ii n_1965_ (
        .a(n_1230_),
        .b(n_1229_),
        .c(n_1231_)
    );

    bfr new_Jinkela_buffer_5081 (
        .din(new_Jinkela_wire_6056),
        .dout(new_Jinkela_wire_6057)
    );

    bfr new_Jinkela_buffer_6729 (
        .din(new_Jinkela_wire_8250),
        .dout(new_Jinkela_wire_8251)
    );

    and_bi n_2683_ (
        .a(new_Jinkela_wire_4095),
        .b(new_Jinkela_wire_8163),
        .c(n_0540_)
    );

    and_bb n_1966_ (
        .a(new_Jinkela_wire_91),
        .b(new_Jinkela_wire_1235),
        .c(n_1232_)
    );

    bfr new_Jinkela_buffer_5120 (
        .din(new_Jinkela_wire_6111),
        .dout(new_Jinkela_wire_6112)
    );

    and_ii n_2684_ (
        .a(n_0540_),
        .b(n_0539_),
        .c(n_0541_)
    );

    bfr new_Jinkela_buffer_5103 (
        .din(new_Jinkela_wire_6080),
        .dout(new_Jinkela_wire_6081)
    );

    and_ii n_1967_ (
        .a(new_Jinkela_wire_8874),
        .b(new_Jinkela_wire_9549),
        .c(n_1233_)
    );

    bfr new_Jinkela_buffer_5082 (
        .din(new_Jinkela_wire_6057),
        .dout(new_Jinkela_wire_6058)
    );

    bfr new_Jinkela_buffer_6730 (
        .din(new_Jinkela_wire_8251),
        .dout(new_Jinkela_wire_8252)
    );

    or_bi n_2685_ (
        .a(new_Jinkela_wire_8308),
        .b(new_Jinkela_wire_8189),
        .c(n_0542_)
    );

    and_bb n_1968_ (
        .a(new_Jinkela_wire_1398),
        .b(new_Jinkela_wire_1208),
        .c(n_1234_)
    );

    bfr new_Jinkela_buffer_6763 (
        .din(new_Jinkela_wire_8338),
        .dout(new_Jinkela_wire_8339)
    );

    and_bi n_2686_ (
        .a(new_Jinkela_wire_8307),
        .b(new_Jinkela_wire_8188),
        .c(n_0543_)
    );

    and_ii n_1969_ (
        .a(new_Jinkela_wire_5882),
        .b(new_Jinkela_wire_4337),
        .c(n_1235_)
    );

    bfr new_Jinkela_buffer_6731 (
        .din(new_Jinkela_wire_8252),
        .dout(new_Jinkela_wire_8253)
    );

    or_bi n_2687_ (
        .a(n_0543_),
        .b(n_0542_),
        .c(n_0544_)
    );

    bfr new_Jinkela_buffer_5104 (
        .din(new_Jinkela_wire_6081),
        .dout(new_Jinkela_wire_6082)
    );

    and_ii n_1970_ (
        .a(new_Jinkela_wire_9383),
        .b(new_Jinkela_wire_4973),
        .c(n_1236_)
    );

    bfr new_Jinkela_buffer_6786 (
        .din(new_Jinkela_wire_8367),
        .dout(new_Jinkela_wire_8368)
    );

    and_bi n_2688_ (
        .a(new_Jinkela_wire_4679),
        .b(new_Jinkela_wire_9424),
        .c(n_0545_)
    );

    and_bb n_1971_ (
        .a(new_Jinkela_wire_9384),
        .b(new_Jinkela_wire_4974),
        .c(n_1237_)
    );

    bfr new_Jinkela_buffer_5121 (
        .din(new_Jinkela_wire_6112),
        .dout(new_Jinkela_wire_6113)
    );

    bfr new_Jinkela_buffer_6732 (
        .din(new_Jinkela_wire_8253),
        .dout(new_Jinkela_wire_8254)
    );

    and_ii n_2689_ (
        .a(n_0545_),
        .b(n_0530_),
        .c(n_0546_)
    );

    bfr new_Jinkela_buffer_5105 (
        .din(new_Jinkela_wire_6082),
        .dout(new_Jinkela_wire_6083)
    );

    and_ii n_1972_ (
        .a(n_1237_),
        .b(n_1236_),
        .c(n_1238_)
    );

    bfr new_Jinkela_buffer_6764 (
        .din(new_Jinkela_wire_8339),
        .dout(new_Jinkela_wire_8340)
    );

    and_bi n_2690_ (
        .a(new_Jinkela_wire_5369),
        .b(new_Jinkela_wire_5923),
        .c(n_0547_)
    );

    and_bi n_1973_ (
        .a(new_Jinkela_wire_6265),
        .b(new_Jinkela_wire_9008),
        .c(n_1239_)
    );

    spl2 new_Jinkela_splitter_387 (
        .a(n_0678_),
        .b(new_Jinkela_wire_6152),
        .c(new_Jinkela_wire_6153)
    );

    bfr new_Jinkela_buffer_6733 (
        .din(new_Jinkela_wire_8254),
        .dout(new_Jinkela_wire_8255)
    );

    and_ii n_2691_ (
        .a(new_Jinkela_wire_5977),
        .b(new_Jinkela_wire_5645),
        .c(n_0548_)
    );

    bfr new_Jinkela_buffer_5106 (
        .din(new_Jinkela_wire_6083),
        .dout(new_Jinkela_wire_6084)
    );

    and_bi n_1974_ (
        .a(new_Jinkela_wire_9007),
        .b(new_Jinkela_wire_6264),
        .c(n_1240_)
    );

    spl2 new_Jinkela_splitter_631 (
        .a(new_Jinkela_wire_8371),
        .b(new_Jinkela_wire_8372),
        .c(new_Jinkela_wire_8373)
    );

    and_bi n_2692_ (
        .a(new_Jinkela_wire_8942),
        .b(new_Jinkela_wire_9400),
        .c(n_0549_)
    );

    bfr new_Jinkela_buffer_5136 (
        .din(new_Jinkela_wire_6134),
        .dout(new_Jinkela_wire_6135)
    );

    and_ii n_1975_ (
        .a(n_1240_),
        .b(n_1239_),
        .c(n_1241_)
    );

    bfr new_Jinkela_buffer_5122 (
        .din(new_Jinkela_wire_6113),
        .dout(new_Jinkela_wire_6114)
    );

    bfr new_Jinkela_buffer_6734 (
        .din(new_Jinkela_wire_8255),
        .dout(new_Jinkela_wire_8256)
    );

    and_bi n_2693_ (
        .a(new_Jinkela_wire_9399),
        .b(new_Jinkela_wire_8943),
        .c(n_0550_)
    );

    spl2 new_Jinkela_splitter_632 (
        .a(n_0019_),
        .b(new_Jinkela_wire_8374),
        .c(new_Jinkela_wire_8378)
    );

    bfr new_Jinkela_buffer_5107 (
        .din(new_Jinkela_wire_6084),
        .dout(new_Jinkela_wire_6085)
    );

    and_bi n_1976_ (
        .a(new_Jinkela_wire_8947),
        .b(new_Jinkela_wire_9013),
        .c(n_1242_)
    );

    bfr new_Jinkela_buffer_6765 (
        .din(new_Jinkela_wire_8340),
        .dout(new_Jinkela_wire_8341)
    );

    and_ii n_2694_ (
        .a(n_0550_),
        .b(n_0549_),
        .c(n_0551_)
    );

    and_bi n_1977_ (
        .a(new_Jinkela_wire_9012),
        .b(new_Jinkela_wire_8946),
        .c(n_1243_)
    );

    bfr new_Jinkela_buffer_6735 (
        .din(new_Jinkela_wire_8256),
        .dout(new_Jinkela_wire_8257)
    );

    and_bb n_2695_ (
        .a(new_Jinkela_wire_5006),
        .b(new_Jinkela_wire_6540),
        .c(n_0552_)
    );

    bfr new_Jinkela_buffer_5108 (
        .din(new_Jinkela_wire_6085),
        .dout(new_Jinkela_wire_6086)
    );

    or_bb n_1978_ (
        .a(n_1243_),
        .b(n_1242_),
        .c(n_1244_)
    );

    and_ii n_2696_ (
        .a(new_Jinkela_wire_5005),
        .b(new_Jinkela_wire_6539),
        .c(n_0553_)
    );

    and_bb n_1979_ (
        .a(new_Jinkela_wire_791),
        .b(new_Jinkela_wire_1357),
        .c(n_1245_)
    );

    bfr new_Jinkela_buffer_5123 (
        .din(new_Jinkela_wire_6114),
        .dout(new_Jinkela_wire_6115)
    );

    bfr new_Jinkela_buffer_6736 (
        .din(new_Jinkela_wire_8257),
        .dout(new_Jinkela_wire_8258)
    );

    and_ii n_2697_ (
        .a(n_0553_),
        .b(n_0552_),
        .c(n_0554_)
    );

    and_ii n_1980_ (
        .a(new_Jinkela_wire_8823),
        .b(new_Jinkela_wire_5067),
        .c(n_1246_)
    );

    bfr new_Jinkela_buffer_5146 (
        .din(new_Jinkela_wire_6155),
        .dout(new_Jinkela_wire_6156)
    );

    bfr new_Jinkela_buffer_6766 (
        .din(new_Jinkela_wire_8341),
        .dout(new_Jinkela_wire_8342)
    );

    and_bi n_2698_ (
        .a(new_Jinkela_wire_6556),
        .b(new_Jinkela_wire_8388),
        .c(n_0555_)
    );

    spl4L new_Jinkela_splitter_385 (
        .a(new_Jinkela_wire_6136),
        .d(new_Jinkela_wire_6137),
        .b(new_Jinkela_wire_6138),
        .e(new_Jinkela_wire_6139),
        .c(new_Jinkela_wire_6140)
    );

    and_bb n_1981_ (
        .a(new_Jinkela_wire_690),
        .b(new_Jinkela_wire_1258),
        .c(n_1247_)
    );

    bfr new_Jinkela_buffer_5124 (
        .din(new_Jinkela_wire_6115),
        .dout(new_Jinkela_wire_6116)
    );

    bfr new_Jinkela_buffer_6737 (
        .din(new_Jinkela_wire_8258),
        .dout(new_Jinkela_wire_8259)
    );

    and_bi n_2699_ (
        .a(new_Jinkela_wire_8387),
        .b(new_Jinkela_wire_6555),
        .c(n_0556_)
    );

    and_bi n_1982_ (
        .a(new_Jinkela_wire_8363),
        .b(new_Jinkela_wire_7997),
        .c(n_1248_)
    );

    and_ii n_2700_ (
        .a(n_0556_),
        .b(n_0555_),
        .c(n_0557_)
    );

    spl2 new_Jinkela_splitter_388 (
        .a(n_1338_),
        .b(new_Jinkela_wire_6154),
        .c(new_Jinkela_wire_6155)
    );

    and_bb n_1983_ (
        .a(new_Jinkela_wire_4857),
        .b(new_Jinkela_wire_9497),
        .c(n_1249_)
    );

    bfr new_Jinkela_buffer_5125 (
        .din(new_Jinkela_wire_6116),
        .dout(new_Jinkela_wire_6117)
    );

    bfr new_Jinkela_buffer_6738 (
        .din(new_Jinkela_wire_8259),
        .dout(new_Jinkela_wire_8260)
    );

    and_bi n_2701_ (
        .a(new_Jinkela_wire_9431),
        .b(new_Jinkela_wire_8891),
        .c(n_0558_)
    );

    and_ii n_1984_ (
        .a(new_Jinkela_wire_4856),
        .b(new_Jinkela_wire_9496),
        .c(n_1250_)
    );

    spl2 new_Jinkela_splitter_386 (
        .a(new_Jinkela_wire_6140),
        .b(new_Jinkela_wire_6141),
        .c(new_Jinkela_wire_6142)
    );

    bfr new_Jinkela_buffer_6767 (
        .din(new_Jinkela_wire_8342),
        .dout(new_Jinkela_wire_8343)
    );

    and_bi n_2702_ (
        .a(new_Jinkela_wire_3685),
        .b(new_Jinkela_wire_6557),
        .c(n_0559_)
    );

    and_ii n_1985_ (
        .a(n_1250_),
        .b(n_1249_),
        .c(n_1251_)
    );

    bfr new_Jinkela_buffer_5126 (
        .din(new_Jinkela_wire_6117),
        .dout(new_Jinkela_wire_6118)
    );

    bfr new_Jinkela_buffer_6739 (
        .din(new_Jinkela_wire_8260),
        .dout(new_Jinkela_wire_8261)
    );

    or_bb n_2703_ (
        .a(n_0559_),
        .b(new_Jinkela_wire_7812),
        .c(n_0560_)
    );

    and_bb n_1986_ (
        .a(new_Jinkela_wire_195),
        .b(new_Jinkela_wire_1330),
        .c(n_1252_)
    );

    bfr new_Jinkela_buffer_6789 (
        .din(n_0554_),
        .dout(new_Jinkela_wire_8384)
    );

    and_bi n_2704_ (
        .a(new_Jinkela_wire_3593),
        .b(new_Jinkela_wire_4487),
        .c(n_0561_)
    );

    bfr new_Jinkela_buffer_5157 (
        .din(new_net_2564),
        .dout(new_Jinkela_wire_6167)
    );

    and_ii n_1987_ (
        .a(new_Jinkela_wire_9548),
        .b(new_Jinkela_wire_7849),
        .c(n_1253_)
    );

    bfr new_Jinkela_buffer_5127 (
        .din(new_Jinkela_wire_6118),
        .dout(new_Jinkela_wire_6119)
    );

    bfr new_Jinkela_buffer_6740 (
        .din(new_Jinkela_wire_8261),
        .dout(new_Jinkela_wire_8262)
    );

    and_ii n_2705_ (
        .a(new_Jinkela_wire_8762),
        .b(new_Jinkela_wire_9929),
        .c(n_0562_)
    );

    and_bb n_1988_ (
        .a(new_Jinkela_wire_1985),
        .b(new_Jinkela_wire_1240),
        .c(n_1254_)
    );

    bfr new_Jinkela_buffer_5137 (
        .din(new_Jinkela_wire_6142),
        .dout(new_Jinkela_wire_6143)
    );

    bfr new_Jinkela_buffer_6768 (
        .din(new_Jinkela_wire_8343),
        .dout(new_Jinkela_wire_8344)
    );

    bfr new_Jinkela_buffer_267 (
        .din(new_Jinkela_wire_291),
        .dout(new_Jinkela_wire_292)
    );

    bfr new_Jinkela_buffer_221 (
        .din(new_Jinkela_wire_240),
        .dout(new_Jinkela_wire_241)
    );

    bfr new_Jinkela_buffer_1764 (
        .din(new_Jinkela_wire_2114),
        .dout(new_Jinkela_wire_2115)
    );

    bfr new_Jinkela_buffer_329 (
        .din(new_Jinkela_wire_358),
        .dout(new_Jinkela_wire_359)
    );

    bfr new_Jinkela_buffer_1820 (
        .din(new_Jinkela_wire_2174),
        .dout(new_Jinkela_wire_2175)
    );

    bfr new_Jinkela_buffer_222 (
        .din(new_Jinkela_wire_241),
        .dout(new_Jinkela_wire_242)
    );

    bfr new_Jinkela_buffer_1765 (
        .din(new_Jinkela_wire_2115),
        .dout(new_Jinkela_wire_2116)
    );

    bfr new_Jinkela_buffer_268 (
        .din(new_Jinkela_wire_292),
        .dout(new_Jinkela_wire_293)
    );

    bfr new_Jinkela_buffer_223 (
        .din(new_Jinkela_wire_242),
        .dout(new_Jinkela_wire_243)
    );

    bfr new_Jinkela_buffer_1766 (
        .din(new_Jinkela_wire_2116),
        .dout(new_Jinkela_wire_2117)
    );

    bfr new_Jinkela_buffer_1821 (
        .din(new_Jinkela_wire_2175),
        .dout(new_Jinkela_wire_2176)
    );

    bfr new_Jinkela_buffer_224 (
        .din(new_Jinkela_wire_243),
        .dout(new_Jinkela_wire_244)
    );

    bfr new_Jinkela_buffer_1767 (
        .din(new_Jinkela_wire_2117),
        .dout(new_Jinkela_wire_2118)
    );

    bfr new_Jinkela_buffer_269 (
        .din(new_Jinkela_wire_293),
        .dout(new_Jinkela_wire_294)
    );

    bfr new_Jinkela_buffer_1884 (
        .din(new_Jinkela_wire_2238),
        .dout(new_Jinkela_wire_2239)
    );

    bfr new_Jinkela_buffer_225 (
        .din(new_Jinkela_wire_244),
        .dout(new_Jinkela_wire_245)
    );

    bfr new_Jinkela_buffer_1768 (
        .din(new_Jinkela_wire_2118),
        .dout(new_Jinkela_wire_2119)
    );

    bfr new_Jinkela_buffer_396 (
        .din(new_Jinkela_wire_427),
        .dout(new_Jinkela_wire_428)
    );

    bfr new_Jinkela_buffer_1822 (
        .din(new_Jinkela_wire_2176),
        .dout(new_Jinkela_wire_2177)
    );

    bfr new_Jinkela_buffer_332 (
        .din(new_Jinkela_wire_361),
        .dout(new_Jinkela_wire_362)
    );

    bfr new_Jinkela_buffer_226 (
        .din(new_Jinkela_wire_245),
        .dout(new_Jinkela_wire_246)
    );

    bfr new_Jinkela_buffer_1769 (
        .din(new_Jinkela_wire_2119),
        .dout(new_Jinkela_wire_2120)
    );

    bfr new_Jinkela_buffer_270 (
        .din(new_Jinkela_wire_294),
        .dout(new_Jinkela_wire_295)
    );

    spl2 new_Jinkela_splitter_114 (
        .a(new_Jinkela_wire_2239),
        .b(new_Jinkela_wire_2240),
        .c(new_Jinkela_wire_2241)
    );

    bfr new_Jinkela_buffer_227 (
        .din(new_Jinkela_wire_246),
        .dout(new_Jinkela_wire_247)
    );

    bfr new_Jinkela_buffer_1770 (
        .din(new_Jinkela_wire_2120),
        .dout(new_Jinkela_wire_2121)
    );

    bfr new_Jinkela_buffer_1823 (
        .din(new_Jinkela_wire_2177),
        .dout(new_Jinkela_wire_2178)
    );

    bfr new_Jinkela_buffer_228 (
        .din(new_Jinkela_wire_247),
        .dout(new_Jinkela_wire_248)
    );

    bfr new_Jinkela_buffer_1771 (
        .din(new_Jinkela_wire_2121),
        .dout(new_Jinkela_wire_2122)
    );

    bfr new_Jinkela_buffer_271 (
        .din(new_Jinkela_wire_295),
        .dout(new_Jinkela_wire_296)
    );

    spl2 new_Jinkela_splitter_115 (
        .a(new_Jinkela_wire_2241),
        .b(new_Jinkela_wire_2242),
        .c(new_Jinkela_wire_2243)
    );

    bfr new_Jinkela_buffer_229 (
        .din(new_Jinkela_wire_248),
        .dout(new_Jinkela_wire_249)
    );

    bfr new_Jinkela_buffer_1772 (
        .din(new_Jinkela_wire_2122),
        .dout(new_Jinkela_wire_2123)
    );

    bfr new_Jinkela_buffer_403 (
        .din(N229),
        .dout(new_Jinkela_wire_435)
    );

    bfr new_Jinkela_buffer_1824 (
        .din(new_Jinkela_wire_2178),
        .dout(new_Jinkela_wire_2179)
    );

    spl2 new_Jinkela_splitter_13 (
        .a(new_Jinkela_wire_362),
        .b(new_Jinkela_wire_363),
        .c(new_Jinkela_wire_364)
    );

    bfr new_Jinkela_buffer_230 (
        .din(new_Jinkela_wire_249),
        .dout(new_Jinkela_wire_250)
    );

    bfr new_Jinkela_buffer_1773 (
        .din(new_Jinkela_wire_2123),
        .dout(new_Jinkela_wire_2124)
    );

    bfr new_Jinkela_buffer_272 (
        .din(new_Jinkela_wire_296),
        .dout(new_Jinkela_wire_297)
    );

    bfr new_Jinkela_buffer_2081 (
        .din(N235),
        .dout(new_Jinkela_wire_2451)
    );

    bfr new_Jinkela_buffer_231 (
        .din(new_Jinkela_wire_250),
        .dout(new_Jinkela_wire_251)
    );

    bfr new_Jinkela_buffer_1774 (
        .din(new_Jinkela_wire_2124),
        .dout(new_Jinkela_wire_2125)
    );

    bfr new_Jinkela_buffer_1825 (
        .din(new_Jinkela_wire_2179),
        .dout(new_Jinkela_wire_2180)
    );

    bfr new_Jinkela_buffer_333 (
        .din(new_Jinkela_wire_364),
        .dout(new_Jinkela_wire_365)
    );

    bfr new_Jinkela_buffer_232 (
        .din(new_Jinkela_wire_251),
        .dout(new_Jinkela_wire_252)
    );

    bfr new_Jinkela_buffer_1775 (
        .din(new_Jinkela_wire_2125),
        .dout(new_Jinkela_wire_2126)
    );

    bfr new_Jinkela_buffer_273 (
        .din(new_Jinkela_wire_297),
        .dout(new_Jinkela_wire_298)
    );

    bfr new_Jinkela_buffer_1946 (
        .din(new_Jinkela_wire_2308),
        .dout(new_Jinkela_wire_2309)
    );

    spl2 new_Jinkela_splitter_116 (
        .a(new_Jinkela_wire_2243),
        .b(new_Jinkela_wire_2244),
        .c(new_Jinkela_wire_2245)
    );

    bfr new_Jinkela_buffer_233 (
        .din(new_Jinkela_wire_252),
        .dout(new_Jinkela_wire_253)
    );

    bfr new_Jinkela_buffer_1776 (
        .din(new_Jinkela_wire_2126),
        .dout(new_Jinkela_wire_2127)
    );

    bfr new_Jinkela_buffer_1826 (
        .din(new_Jinkela_wire_2180),
        .dout(new_Jinkela_wire_2181)
    );

    bfr new_Jinkela_buffer_234 (
        .din(new_Jinkela_wire_253),
        .dout(new_Jinkela_wire_254)
    );

    bfr new_Jinkela_buffer_1777 (
        .din(new_Jinkela_wire_2127),
        .dout(new_Jinkela_wire_2128)
    );

    bfr new_Jinkela_buffer_274 (
        .din(new_Jinkela_wire_298),
        .dout(new_Jinkela_wire_299)
    );

    bfr new_Jinkela_buffer_235 (
        .din(new_Jinkela_wire_254),
        .dout(new_Jinkela_wire_255)
    );

    bfr new_Jinkela_buffer_1778 (
        .din(new_Jinkela_wire_2128),
        .dout(new_Jinkela_wire_2129)
    );

    bfr new_Jinkela_buffer_397 (
        .din(new_Jinkela_wire_428),
        .dout(new_Jinkela_wire_429)
    );

    bfr new_Jinkela_buffer_1827 (
        .din(new_Jinkela_wire_2181),
        .dout(new_Jinkela_wire_2182)
    );

    bfr new_Jinkela_buffer_236 (
        .din(new_Jinkela_wire_255),
        .dout(new_Jinkela_wire_256)
    );

    bfr new_Jinkela_buffer_1779 (
        .din(new_Jinkela_wire_2129),
        .dout(new_Jinkela_wire_2130)
    );

    bfr new_Jinkela_buffer_275 (
        .din(new_Jinkela_wire_299),
        .dout(new_Jinkela_wire_300)
    );

    bfr new_Jinkela_buffer_2010 (
        .din(new_Jinkela_wire_2374),
        .dout(new_Jinkela_wire_2375)
    );

    bfr new_Jinkela_buffer_1885 (
        .din(new_Jinkela_wire_2245),
        .dout(new_Jinkela_wire_2246)
    );

    bfr new_Jinkela_buffer_237 (
        .din(new_Jinkela_wire_256),
        .dout(new_Jinkela_wire_257)
    );

    bfr new_Jinkela_buffer_1780 (
        .din(new_Jinkela_wire_2130),
        .dout(new_Jinkela_wire_2131)
    );

    bfr new_Jinkela_buffer_400 (
        .din(new_Jinkela_wire_431),
        .dout(new_Jinkela_wire_432)
    );

    bfr new_Jinkela_buffer_1828 (
        .din(new_Jinkela_wire_2182),
        .dout(new_Jinkela_wire_2183)
    );

    bfr new_Jinkela_buffer_334 (
        .din(new_Jinkela_wire_365),
        .dout(new_Jinkela_wire_366)
    );

    bfr new_Jinkela_buffer_238 (
        .din(new_Jinkela_wire_257),
        .dout(new_Jinkela_wire_258)
    );

    bfr new_Jinkela_buffer_1781 (
        .din(new_Jinkela_wire_2131),
        .dout(new_Jinkela_wire_2132)
    );

    bfr new_Jinkela_buffer_276 (
        .din(new_Jinkela_wire_300),
        .dout(new_Jinkela_wire_301)
    );

    bfr new_Jinkela_buffer_2014 (
        .din(new_Jinkela_wire_2378),
        .dout(new_Jinkela_wire_2379)
    );

    bfr new_Jinkela_buffer_239 (
        .din(new_Jinkela_wire_258),
        .dout(new_Jinkela_wire_259)
    );

    bfr new_Jinkela_buffer_1782 (
        .din(new_Jinkela_wire_2132),
        .dout(new_Jinkela_wire_2133)
    );

    bfr new_Jinkela_buffer_1829 (
        .din(new_Jinkela_wire_2183),
        .dout(new_Jinkela_wire_2184)
    );

    bfr new_Jinkela_buffer_240 (
        .din(new_Jinkela_wire_259),
        .dout(new_Jinkela_wire_260)
    );

    bfr new_Jinkela_buffer_1783 (
        .din(new_Jinkela_wire_2133),
        .dout(new_Jinkela_wire_2134)
    );

    bfr new_Jinkela_buffer_277 (
        .din(new_Jinkela_wire_301),
        .dout(new_Jinkela_wire_302)
    );

    spl2 new_Jinkela_splitter_118 (
        .a(new_Jinkela_wire_2309),
        .b(new_Jinkela_wire_2310),
        .c(new_Jinkela_wire_2311)
    );

    bfr new_Jinkela_buffer_241 (
        .din(new_Jinkela_wire_260),
        .dout(new_Jinkela_wire_261)
    );

    bfr new_Jinkela_buffer_1784 (
        .din(new_Jinkela_wire_2134),
        .dout(new_Jinkela_wire_2135)
    );

    bfr new_Jinkela_buffer_5920 (
        .din(new_Jinkela_wire_7159),
        .dout(new_Jinkela_wire_7160)
    );

    spl2 new_Jinkela_splitter_493 (
        .a(n_0896_),
        .b(new_Jinkela_wire_7244),
        .c(new_Jinkela_wire_7245)
    );

    bfr new_Jinkela_buffer_5921 (
        .din(new_Jinkela_wire_7160),
        .dout(new_Jinkela_wire_7161)
    );

    bfr new_Jinkela_buffer_5976 (
        .din(new_Jinkela_wire_7228),
        .dout(new_Jinkela_wire_7229)
    );

    bfr new_Jinkela_buffer_5922 (
        .din(new_Jinkela_wire_7161),
        .dout(new_Jinkela_wire_7162)
    );

    bfr new_Jinkela_buffer_5977 (
        .din(new_Jinkela_wire_7229),
        .dout(new_Jinkela_wire_7230)
    );

    bfr new_Jinkela_buffer_5923 (
        .din(new_Jinkela_wire_7162),
        .dout(new_Jinkela_wire_7163)
    );

    bfr new_Jinkela_buffer_5980 (
        .din(new_Jinkela_wire_7236),
        .dout(new_Jinkela_wire_7237)
    );

    bfr new_Jinkela_buffer_5924 (
        .din(new_Jinkela_wire_7163),
        .dout(new_Jinkela_wire_7164)
    );

    bfr new_Jinkela_buffer_5978 (
        .din(new_Jinkela_wire_7230),
        .dout(new_Jinkela_wire_7231)
    );

    bfr new_Jinkela_buffer_5925 (
        .din(new_Jinkela_wire_7164),
        .dout(new_Jinkela_wire_7165)
    );

    spl3L new_Jinkela_splitter_494 (
        .a(n_1102_),
        .d(new_Jinkela_wire_7246),
        .b(new_Jinkela_wire_7247),
        .c(new_Jinkela_wire_7248)
    );

    bfr new_Jinkela_buffer_5926 (
        .din(new_Jinkela_wire_7165),
        .dout(new_Jinkela_wire_7166)
    );

    bfr new_Jinkela_buffer_5983 (
        .din(new_Jinkela_wire_7241),
        .dout(new_Jinkela_wire_7242)
    );

    spl2 new_Jinkela_splitter_490 (
        .a(new_Jinkela_wire_7231),
        .b(new_Jinkela_wire_7232),
        .c(new_Jinkela_wire_7233)
    );

    bfr new_Jinkela_buffer_5927 (
        .din(new_Jinkela_wire_7166),
        .dout(new_Jinkela_wire_7167)
    );

    bfr new_Jinkela_buffer_5928 (
        .din(new_Jinkela_wire_7167),
        .dout(new_Jinkela_wire_7168)
    );

    bfr new_Jinkela_buffer_5981 (
        .din(new_Jinkela_wire_7237),
        .dout(new_Jinkela_wire_7238)
    );

    bfr new_Jinkela_buffer_5929 (
        .din(new_Jinkela_wire_7168),
        .dout(new_Jinkela_wire_7169)
    );

    spl2 new_Jinkela_splitter_492 (
        .a(new_Jinkela_wire_7238),
        .b(new_Jinkela_wire_7239),
        .c(new_Jinkela_wire_7240)
    );

    bfr new_Jinkela_buffer_5930 (
        .din(new_Jinkela_wire_7169),
        .dout(new_Jinkela_wire_7170)
    );

    bfr new_Jinkela_buffer_5931 (
        .din(new_Jinkela_wire_7170),
        .dout(new_Jinkela_wire_7171)
    );

    bfr new_Jinkela_buffer_5932 (
        .din(new_Jinkela_wire_7171),
        .dout(new_Jinkela_wire_7172)
    );

    bfr new_Jinkela_buffer_5984 (
        .din(new_Jinkela_wire_7242),
        .dout(new_Jinkela_wire_7243)
    );

    spl2 new_Jinkela_splitter_0 (
        .a(N1),
        .b(new_Jinkela_wire_0),
        .c(new_Jinkela_wire_1)
    );

    spl2 new_Jinkela_splitter_496 (
        .a(n_0546_),
        .b(new_Jinkela_wire_7251),
        .c(new_Jinkela_wire_7252)
    );

    bfr new_Jinkela_buffer_5933 (
        .din(new_Jinkela_wire_7172),
        .dout(new_Jinkela_wire_7173)
    );

    bfr new_Jinkela_buffer_64 (
        .din(N160),
        .dout(new_Jinkela_wire_72)
    );

    bfr new_Jinkela_buffer_5985 (
        .din(new_net_2545),
        .dout(new_Jinkela_wire_7253)
    );

    spl2 new_Jinkela_splitter_2 (
        .a(N164),
        .b(new_Jinkela_wire_70),
        .c(new_Jinkela_wire_71)
    );

    bfr new_Jinkela_buffer_5986 (
        .din(new_Jinkela_wire_7253),
        .dout(new_Jinkela_wire_7254)
    );

    bfr new_Jinkela_buffer_5934 (
        .din(new_Jinkela_wire_7173),
        .dout(new_Jinkela_wire_7174)
    );

    bfr new_Jinkela_buffer_68 (
        .din(N82),
        .dout(new_Jinkela_wire_76)
    );

    spl2 new_Jinkela_splitter_495 (
        .a(new_Jinkela_wire_7248),
        .b(new_Jinkela_wire_7249),
        .c(new_Jinkela_wire_7250)
    );

    bfr new_Jinkela_buffer_1 (
        .din(new_Jinkela_wire_2),
        .dout(new_Jinkela_wire_3)
    );

    spl4L new_Jinkela_splitter_498 (
        .a(n_0689_),
        .d(new_Jinkela_wire_7264),
        .b(new_Jinkela_wire_7265),
        .e(new_Jinkela_wire_7266),
        .c(new_Jinkela_wire_7267)
    );

    bfr new_Jinkela_buffer_5935 (
        .din(new_Jinkela_wire_7174),
        .dout(new_Jinkela_wire_7175)
    );

    bfr new_Jinkela_buffer_65 (
        .din(new_Jinkela_wire_72),
        .dout(new_Jinkela_wire_73)
    );

    bfr new_Jinkela_buffer_2 (
        .din(new_Jinkela_wire_3),
        .dout(new_Jinkela_wire_4)
    );

    bfr new_Jinkela_buffer_5936 (
        .din(new_Jinkela_wire_7175),
        .dout(new_Jinkela_wire_7176)
    );

    bfr new_Jinkela_buffer_72 (
        .din(N84),
        .dout(new_Jinkela_wire_80)
    );

    bfr new_Jinkela_buffer_3 (
        .din(new_Jinkela_wire_4),
        .dout(new_Jinkela_wire_5)
    );

    spl2 new_Jinkela_splitter_497 (
        .a(n_0377_),
        .b(new_Jinkela_wire_7262),
        .c(new_Jinkela_wire_7263)
    );

    bfr new_Jinkela_buffer_5937 (
        .din(new_Jinkela_wire_7176),
        .dout(new_Jinkela_wire_7177)
    );

    bfr new_Jinkela_buffer_66 (
        .din(new_Jinkela_wire_73),
        .dout(new_Jinkela_wire_74)
    );

    spl4L new_Jinkela_splitter_500 (
        .a(n_1255_),
        .d(new_Jinkela_wire_7270),
        .b(new_Jinkela_wire_7271),
        .e(new_Jinkela_wire_7272),
        .c(new_Jinkela_wire_7273)
    );

    bfr new_Jinkela_buffer_4 (
        .din(new_Jinkela_wire_5),
        .dout(new_Jinkela_wire_6)
    );

    bfr new_Jinkela_buffer_5938 (
        .din(new_Jinkela_wire_7177),
        .dout(new_Jinkela_wire_7178)
    );

    bfr new_Jinkela_buffer_69 (
        .din(new_Jinkela_wire_76),
        .dout(new_Jinkela_wire_77)
    );

    bfr new_Jinkela_buffer_5987 (
        .din(new_Jinkela_wire_7254),
        .dout(new_Jinkela_wire_7255)
    );

    bfr new_Jinkela_buffer_5 (
        .din(new_Jinkela_wire_6),
        .dout(new_Jinkela_wire_7)
    );

    bfr new_Jinkela_buffer_5939 (
        .din(new_Jinkela_wire_7178),
        .dout(new_Jinkela_wire_7179)
    );

    bfr new_Jinkela_buffer_67 (
        .din(new_Jinkela_wire_74),
        .dout(new_Jinkela_wire_75)
    );

    bfr new_Jinkela_buffer_6 (
        .din(new_Jinkela_wire_7),
        .dout(new_Jinkela_wire_8)
    );

    spl2 new_Jinkela_splitter_499 (
        .a(n_0402_),
        .b(new_Jinkela_wire_7268),
        .c(new_Jinkela_wire_7269)
    );

    bfr new_Jinkela_buffer_5940 (
        .din(new_Jinkela_wire_7179),
        .dout(new_Jinkela_wire_7180)
    );

    bfr new_Jinkela_buffer_76 (
        .din(N174),
        .dout(new_Jinkela_wire_84)
    );

    bfr new_Jinkela_buffer_5988 (
        .din(new_Jinkela_wire_7255),
        .dout(new_Jinkela_wire_7256)
    );

    bfr new_Jinkela_buffer_0 (
        .din(new_Jinkela_wire_1),
        .dout(new_Jinkela_wire_2)
    );

    bfr new_Jinkela_buffer_3411 (
        .din(new_Jinkela_wire_3972),
        .dout(new_Jinkela_wire_3973)
    );

    bfr new_Jinkela_buffer_4256 (
        .din(new_Jinkela_wire_5024),
        .dout(new_Jinkela_wire_5025)
    );

    bfr new_Jinkela_buffer_7896 (
        .din(new_Jinkela_wire_9963),
        .dout(new_Jinkela_wire_9964)
    );

    bfr new_Jinkela_buffer_4291 (
        .din(new_Jinkela_wire_5073),
        .dout(new_Jinkela_wire_5074)
    );

    bfr new_Jinkela_buffer_7877 (
        .din(new_Jinkela_wire_9938),
        .dout(new_Jinkela_wire_9939)
    );

    bfr new_Jinkela_buffer_3412 (
        .din(new_Jinkela_wire_3973),
        .dout(new_Jinkela_wire_3974)
    );

    bfr new_Jinkela_buffer_4257 (
        .din(new_Jinkela_wire_5025),
        .dout(new_Jinkela_wire_5026)
    );

    bfr new_Jinkela_buffer_7916 (
        .din(new_Jinkela_wire_9985),
        .dout(new_Jinkela_wire_9986)
    );

    bfr new_Jinkela_buffer_3452 (
        .din(new_Jinkela_wire_4024),
        .dout(new_Jinkela_wire_4025)
    );

    bfr new_Jinkela_buffer_4290 (
        .din(new_net_2527),
        .dout(new_Jinkela_wire_5073)
    );

    bfr new_Jinkela_buffer_7878 (
        .din(new_Jinkela_wire_9939),
        .dout(new_Jinkela_wire_9940)
    );

    bfr new_Jinkela_buffer_3413 (
        .din(new_Jinkela_wire_3974),
        .dout(new_Jinkela_wire_3975)
    );

    spl2 new_Jinkela_splitter_295 (
        .a(n_0462_),
        .b(new_Jinkela_wire_5092),
        .c(new_Jinkela_wire_5093)
    );

    bfr new_Jinkela_buffer_4258 (
        .din(new_Jinkela_wire_5026),
        .dout(new_Jinkela_wire_5027)
    );

    bfr new_Jinkela_buffer_7897 (
        .din(new_Jinkela_wire_9964),
        .dout(new_Jinkela_wire_9965)
    );

    bfr new_Jinkela_buffer_3492 (
        .din(new_Jinkela_wire_4070),
        .dout(new_Jinkela_wire_4071)
    );

    bfr new_Jinkela_buffer_7879 (
        .din(new_Jinkela_wire_9940),
        .dout(new_Jinkela_wire_9941)
    );

    bfr new_Jinkela_buffer_3414 (
        .din(new_Jinkela_wire_3975),
        .dout(new_Jinkela_wire_3976)
    );

    spl2 new_Jinkela_splitter_293 (
        .a(n_1348_),
        .b(new_Jinkela_wire_5087),
        .c(new_Jinkela_wire_5088)
    );

    bfr new_Jinkela_buffer_4259 (
        .din(new_Jinkela_wire_5027),
        .dout(new_Jinkela_wire_5028)
    );

    bfr new_Jinkela_buffer_3453 (
        .din(new_Jinkela_wire_4025),
        .dout(new_Jinkela_wire_4026)
    );

    bfr new_Jinkela_buffer_7880 (
        .din(new_Jinkela_wire_9941),
        .dout(new_Jinkela_wire_9942)
    );

    bfr new_Jinkela_buffer_3415 (
        .din(new_Jinkela_wire_3976),
        .dout(new_Jinkela_wire_3977)
    );

    bfr new_Jinkela_buffer_4305 (
        .din(n_1261_),
        .dout(new_Jinkela_wire_5094)
    );

    bfr new_Jinkela_buffer_4260 (
        .din(new_Jinkela_wire_5028),
        .dout(new_Jinkela_wire_5029)
    );

    bfr new_Jinkela_buffer_7960 (
        .din(new_net_2499),
        .dout(new_Jinkela_wire_10033)
    );

    bfr new_Jinkela_buffer_7898 (
        .din(new_Jinkela_wire_9965),
        .dout(new_Jinkela_wire_9966)
    );

    spl3L new_Jinkela_splitter_212 (
        .a(n_0382_),
        .d(new_Jinkela_wire_4088),
        .b(new_Jinkela_wire_4089),
        .c(new_Jinkela_wire_4090)
    );

    spl2 new_Jinkela_splitter_294 (
        .a(new_Jinkela_wire_5088),
        .b(new_Jinkela_wire_5089),
        .c(new_Jinkela_wire_5090)
    );

    bfr new_Jinkela_buffer_7881 (
        .din(new_Jinkela_wire_9942),
        .dout(new_Jinkela_wire_9943)
    );

    bfr new_Jinkela_buffer_3416 (
        .din(new_Jinkela_wire_3977),
        .dout(new_Jinkela_wire_3978)
    );

    bfr new_Jinkela_buffer_4292 (
        .din(new_Jinkela_wire_5074),
        .dout(new_Jinkela_wire_5075)
    );

    bfr new_Jinkela_buffer_4261 (
        .din(new_Jinkela_wire_5029),
        .dout(new_Jinkela_wire_5030)
    );

    bfr new_Jinkela_buffer_3476 (
        .din(new_Jinkela_wire_4052),
        .dout(new_Jinkela_wire_4053)
    );

    spl4L new_Jinkela_splitter_832 (
        .a(n_1280_),
        .d(new_Jinkela_wire_10097),
        .b(new_Jinkela_wire_10098),
        .e(new_Jinkela_wire_10099),
        .c(new_Jinkela_wire_10100)
    );

    bfr new_Jinkela_buffer_3454 (
        .din(new_Jinkela_wire_4026),
        .dout(new_Jinkela_wire_4027)
    );

    bfr new_Jinkela_buffer_7882 (
        .din(new_Jinkela_wire_9943),
        .dout(new_Jinkela_wire_9944)
    );

    bfr new_Jinkela_buffer_3417 (
        .din(new_Jinkela_wire_3978),
        .dout(new_Jinkela_wire_3979)
    );

    bfr new_Jinkela_buffer_4262 (
        .din(new_Jinkela_wire_5030),
        .dout(new_Jinkela_wire_5031)
    );

    bfr new_Jinkela_buffer_8024 (
        .din(n_0802_),
        .dout(new_Jinkela_wire_10101)
    );

    bfr new_Jinkela_buffer_7899 (
        .din(new_Jinkela_wire_9966),
        .dout(new_Jinkela_wire_9967)
    );

    spl3L new_Jinkela_splitter_297 (
        .a(n_0752_),
        .d(new_Jinkela_wire_5097),
        .b(new_Jinkela_wire_5098),
        .c(new_Jinkela_wire_5099)
    );

    bfr new_Jinkela_buffer_7883 (
        .din(new_Jinkela_wire_9944),
        .dout(new_Jinkela_wire_9945)
    );

    bfr new_Jinkela_buffer_3418 (
        .din(new_Jinkela_wire_3979),
        .dout(new_Jinkela_wire_3980)
    );

    bfr new_Jinkela_buffer_4293 (
        .din(new_Jinkela_wire_5075),
        .dout(new_Jinkela_wire_5076)
    );

    bfr new_Jinkela_buffer_4263 (
        .din(new_Jinkela_wire_5031),
        .dout(new_Jinkela_wire_5032)
    );

    bfr new_Jinkela_buffer_7917 (
        .din(new_Jinkela_wire_9986),
        .dout(new_Jinkela_wire_9987)
    );

    bfr new_Jinkela_buffer_3455 (
        .din(new_Jinkela_wire_4027),
        .dout(new_Jinkela_wire_4028)
    );

    bfr new_Jinkela_buffer_7884 (
        .din(new_Jinkela_wire_9945),
        .dout(new_Jinkela_wire_9946)
    );

    bfr new_Jinkela_buffer_3419 (
        .din(new_Jinkela_wire_3980),
        .dout(new_Jinkela_wire_3981)
    );

    spl2 new_Jinkela_splitter_298 (
        .a(new_Jinkela_wire_5099),
        .b(new_Jinkela_wire_5100),
        .c(new_Jinkela_wire_5101)
    );

    bfr new_Jinkela_buffer_4264 (
        .din(new_Jinkela_wire_5032),
        .dout(new_Jinkela_wire_5033)
    );

    bfr new_Jinkela_buffer_7900 (
        .din(new_Jinkela_wire_9967),
        .dout(new_Jinkela_wire_9968)
    );

    bfr new_Jinkela_buffer_3493 (
        .din(new_Jinkela_wire_4071),
        .dout(new_Jinkela_wire_4072)
    );

    bfr new_Jinkela_buffer_7885 (
        .din(new_Jinkela_wire_9946),
        .dout(new_Jinkela_wire_9947)
    );

    bfr new_Jinkela_buffer_3420 (
        .din(new_Jinkela_wire_3981),
        .dout(new_Jinkela_wire_3982)
    );

    bfr new_Jinkela_buffer_4294 (
        .din(new_Jinkela_wire_5076),
        .dout(new_Jinkela_wire_5077)
    );

    bfr new_Jinkela_buffer_4265 (
        .din(new_Jinkela_wire_5033),
        .dout(new_Jinkela_wire_5034)
    );

    bfr new_Jinkela_buffer_3477 (
        .din(new_Jinkela_wire_4053),
        .dout(new_Jinkela_wire_4054)
    );

    bfr new_Jinkela_buffer_7961 (
        .din(new_Jinkela_wire_10033),
        .dout(new_Jinkela_wire_10034)
    );

    bfr new_Jinkela_buffer_3456 (
        .din(new_Jinkela_wire_4028),
        .dout(new_Jinkela_wire_4029)
    );

    bfr new_Jinkela_buffer_7886 (
        .din(new_Jinkela_wire_9947),
        .dout(new_Jinkela_wire_9948)
    );

    bfr new_Jinkela_buffer_3421 (
        .din(new_Jinkela_wire_3982),
        .dout(new_Jinkela_wire_3983)
    );

    bfr new_Jinkela_buffer_4304 (
        .din(new_Jinkela_wire_5090),
        .dout(new_Jinkela_wire_5091)
    );

    bfr new_Jinkela_buffer_4266 (
        .din(new_Jinkela_wire_5034),
        .dout(new_Jinkela_wire_5035)
    );

    bfr new_Jinkela_buffer_7901 (
        .din(new_Jinkela_wire_9968),
        .dout(new_Jinkela_wire_9969)
    );

    bfr new_Jinkela_buffer_7887 (
        .din(new_Jinkela_wire_9948),
        .dout(new_Jinkela_wire_9949)
    );

    bfr new_Jinkela_buffer_3422 (
        .din(new_Jinkela_wire_3983),
        .dout(new_Jinkela_wire_3984)
    );

    bfr new_Jinkela_buffer_4295 (
        .din(new_Jinkela_wire_5077),
        .dout(new_Jinkela_wire_5078)
    );

    bfr new_Jinkela_buffer_4267 (
        .din(new_Jinkela_wire_5035),
        .dout(new_Jinkela_wire_5036)
    );

    bfr new_Jinkela_buffer_7918 (
        .din(new_Jinkela_wire_9987),
        .dout(new_Jinkela_wire_9988)
    );

    bfr new_Jinkela_buffer_3457 (
        .din(new_Jinkela_wire_4029),
        .dout(new_Jinkela_wire_4030)
    );

    bfr new_Jinkela_buffer_7888 (
        .din(new_Jinkela_wire_9949),
        .dout(new_Jinkela_wire_9950)
    );

    bfr new_Jinkela_buffer_3423 (
        .din(new_Jinkela_wire_3984),
        .dout(new_Jinkela_wire_3985)
    );

    bfr new_Jinkela_buffer_4268 (
        .din(new_Jinkela_wire_5036),
        .dout(new_Jinkela_wire_5037)
    );

    bfr new_Jinkela_buffer_7902 (
        .din(new_Jinkela_wire_9969),
        .dout(new_Jinkela_wire_9970)
    );

    bfr new_Jinkela_buffer_7889 (
        .din(new_Jinkela_wire_9950),
        .dout(new_Jinkela_wire_9951)
    );

    bfr new_Jinkela_buffer_3424 (
        .din(new_Jinkela_wire_3985),
        .dout(new_Jinkela_wire_3986)
    );

    bfr new_Jinkela_buffer_4296 (
        .din(new_Jinkela_wire_5078),
        .dout(new_Jinkela_wire_5079)
    );

    bfr new_Jinkela_buffer_4269 (
        .din(new_Jinkela_wire_5037),
        .dout(new_Jinkela_wire_5038)
    );

    bfr new_Jinkela_buffer_3478 (
        .din(new_Jinkela_wire_4054),
        .dout(new_Jinkela_wire_4055)
    );

    bfr new_Jinkela_buffer_3458 (
        .din(new_Jinkela_wire_4030),
        .dout(new_Jinkela_wire_4031)
    );

    bfr new_Jinkela_buffer_7890 (
        .din(new_Jinkela_wire_9951),
        .dout(new_Jinkela_wire_9952)
    );

    bfr new_Jinkela_buffer_3425 (
        .din(new_Jinkela_wire_3986),
        .dout(new_Jinkela_wire_3987)
    );

    spl2 new_Jinkela_splitter_296 (
        .a(n_1132_),
        .b(new_Jinkela_wire_5095),
        .c(new_Jinkela_wire_5096)
    );

    bfr new_Jinkela_buffer_4270 (
        .din(new_Jinkela_wire_5038),
        .dout(new_Jinkela_wire_5039)
    );

    bfr new_Jinkela_buffer_7903 (
        .din(new_Jinkela_wire_9970),
        .dout(new_Jinkela_wire_9971)
    );

    bfr new_Jinkela_buffer_7891 (
        .din(new_Jinkela_wire_9952),
        .dout(new_Jinkela_wire_9953)
    );

    bfr new_Jinkela_buffer_3426 (
        .din(new_Jinkela_wire_3987),
        .dout(new_Jinkela_wire_3988)
    );

    bfr new_Jinkela_buffer_4297 (
        .din(new_Jinkela_wire_5079),
        .dout(new_Jinkela_wire_5080)
    );

    bfr new_Jinkela_buffer_4271 (
        .din(new_Jinkela_wire_5039),
        .dout(new_Jinkela_wire_5040)
    );

    spl3L new_Jinkela_splitter_211 (
        .a(n_1216_),
        .d(new_Jinkela_wire_4085),
        .b(new_Jinkela_wire_4086),
        .c(new_Jinkela_wire_4087)
    );

    bfr new_Jinkela_buffer_7919 (
        .din(new_Jinkela_wire_9988),
        .dout(new_Jinkela_wire_9989)
    );

    bfr new_Jinkela_buffer_3459 (
        .din(new_Jinkela_wire_4031),
        .dout(new_Jinkela_wire_4032)
    );

    bfr new_Jinkela_buffer_7892 (
        .din(new_Jinkela_wire_9953),
        .dout(new_Jinkela_wire_9954)
    );

    bfr new_Jinkela_buffer_3427 (
        .din(new_Jinkela_wire_3988),
        .dout(new_Jinkela_wire_3989)
    );

    bfr new_Jinkela_buffer_4272 (
        .din(new_Jinkela_wire_5040),
        .dout(new_Jinkela_wire_5041)
    );

    bfr new_Jinkela_buffer_7904 (
        .din(new_Jinkela_wire_9971),
        .dout(new_Jinkela_wire_9972)
    );

    bfr new_Jinkela_buffer_3494 (
        .din(new_Jinkela_wire_4072),
        .dout(new_Jinkela_wire_4073)
    );

    bfr new_Jinkela_buffer_3428 (
        .din(new_Jinkela_wire_3989),
        .dout(new_Jinkela_wire_3990)
    );

    bfr new_Jinkela_buffer_4298 (
        .din(new_Jinkela_wire_5080),
        .dout(new_Jinkela_wire_5081)
    );

    spl2 new_Jinkela_splitter_833 (
        .a(n_0629_),
        .b(new_Jinkela_wire_10102),
        .c(new_Jinkela_wire_10103)
    );

    bfr new_Jinkela_buffer_4273 (
        .din(new_Jinkela_wire_5041),
        .dout(new_Jinkela_wire_5042)
    );

    bfr new_Jinkela_buffer_7962 (
        .din(new_Jinkela_wire_10034),
        .dout(new_Jinkela_wire_10035)
    );

    bfr new_Jinkela_buffer_3479 (
        .din(new_Jinkela_wire_4055),
        .dout(new_Jinkela_wire_4056)
    );

    bfr new_Jinkela_buffer_7905 (
        .din(new_Jinkela_wire_9972),
        .dout(new_Jinkela_wire_9973)
    );

    bfr new_Jinkela_buffer_3460 (
        .din(new_Jinkela_wire_4032),
        .dout(new_Jinkela_wire_4033)
    );

    bfr new_Jinkela_buffer_3429 (
        .din(new_Jinkela_wire_3990),
        .dout(new_Jinkela_wire_3991)
    );

    spl2 new_Jinkela_splitter_299 (
        .a(n_1214_),
        .b(new_Jinkela_wire_5102),
        .c(new_Jinkela_wire_5103)
    );

    bfr new_Jinkela_buffer_7920 (
        .din(new_Jinkela_wire_9989),
        .dout(new_Jinkela_wire_9990)
    );

    bfr new_Jinkela_buffer_4274 (
        .din(new_Jinkela_wire_5042),
        .dout(new_Jinkela_wire_5043)
    );

    bfr new_Jinkela_buffer_7906 (
        .din(new_Jinkela_wire_9973),
        .dout(new_Jinkela_wire_9974)
    );

    spl3L new_Jinkela_splitter_300 (
        .a(n_0034_),
        .d(new_Jinkela_wire_5106),
        .b(new_Jinkela_wire_5107),
        .c(new_Jinkela_wire_5108)
    );

    bfr new_Jinkela_buffer_3430 (
        .din(new_Jinkela_wire_3991),
        .dout(new_Jinkela_wire_3992)
    );

    bfr new_Jinkela_buffer_4299 (
        .din(new_Jinkela_wire_5081),
        .dout(new_Jinkela_wire_5082)
    );

    bfr new_Jinkela_buffer_4275 (
        .din(new_Jinkela_wire_5043),
        .dout(new_Jinkela_wire_5044)
    );

    bfr new_Jinkela_buffer_7907 (
        .din(new_Jinkela_wire_9974),
        .dout(new_Jinkela_wire_9975)
    );

    bfr new_Jinkela_buffer_3461 (
        .din(new_Jinkela_wire_4033),
        .dout(new_Jinkela_wire_4034)
    );

    bfr new_Jinkela_buffer_3431 (
        .din(new_Jinkela_wire_3992),
        .dout(new_Jinkela_wire_3993)
    );

    bfr new_Jinkela_buffer_7921 (
        .din(new_Jinkela_wire_9990),
        .dout(new_Jinkela_wire_9991)
    );

    bfr new_Jinkela_buffer_4276 (
        .din(new_Jinkela_wire_5044),
        .dout(new_Jinkela_wire_5045)
    );

    bfr new_Jinkela_buffer_7908 (
        .din(new_Jinkela_wire_9975),
        .dout(new_Jinkela_wire_9976)
    );

    spl2 new_Jinkela_splitter_210 (
        .a(new_Jinkela_wire_4081),
        .b(new_Jinkela_wire_4082),
        .c(new_Jinkela_wire_4083)
    );

    bfr new_Jinkela_buffer_4306 (
        .din(new_Jinkela_wire_5103),
        .dout(new_Jinkela_wire_5104)
    );

    bfr new_Jinkela_buffer_2535 (
        .din(new_Jinkela_wire_2936),
        .dout(new_Jinkela_wire_2937)
    );

    bfr new_Jinkela_buffer_6741 (
        .din(new_Jinkela_wire_8262),
        .dout(new_Jinkela_wire_8263)
    );

    bfr new_Jinkela_buffer_6792 (
        .din(n_0241_),
        .dout(new_Jinkela_wire_8389)
    );

    spl3L new_Jinkela_splitter_633 (
        .a(new_Jinkela_wire_8374),
        .d(new_Jinkela_wire_8375),
        .b(new_Jinkela_wire_8376),
        .c(new_Jinkela_wire_8377)
    );

    bfr new_Jinkela_buffer_2536 (
        .din(new_Jinkela_wire_2937),
        .dout(new_Jinkela_wire_2938)
    );

    bfr new_Jinkela_buffer_6769 (
        .din(new_Jinkela_wire_8344),
        .dout(new_Jinkela_wire_8345)
    );

    bfr new_Jinkela_buffer_2779 (
        .din(N171),
        .dout(new_Jinkela_wire_3194)
    );

    bfr new_Jinkela_buffer_2587 (
        .din(new_Jinkela_wire_2992),
        .dout(new_Jinkela_wire_2993)
    );

    bfr new_Jinkela_buffer_6790 (
        .din(new_Jinkela_wire_8384),
        .dout(new_Jinkela_wire_8385)
    );

    bfr new_Jinkela_buffer_2537 (
        .din(new_Jinkela_wire_2938),
        .dout(new_Jinkela_wire_2939)
    );

    bfr new_Jinkela_buffer_6770 (
        .din(new_Jinkela_wire_8345),
        .dout(new_Jinkela_wire_8346)
    );

    bfr new_Jinkela_buffer_2538 (
        .din(new_Jinkela_wire_2939),
        .dout(new_Jinkela_wire_2940)
    );

    bfr new_Jinkela_buffer_6771 (
        .din(new_Jinkela_wire_8346),
        .dout(new_Jinkela_wire_8347)
    );

    bfr new_Jinkela_buffer_2646 (
        .din(new_Jinkela_wire_3055),
        .dout(new_Jinkela_wire_3056)
    );

    bfr new_Jinkela_buffer_2588 (
        .din(new_Jinkela_wire_2993),
        .dout(new_Jinkela_wire_2994)
    );

    spl4L new_Jinkela_splitter_634 (
        .a(new_Jinkela_wire_8378),
        .d(new_Jinkela_wire_8379),
        .b(new_Jinkela_wire_8380),
        .e(new_Jinkela_wire_8381),
        .c(new_Jinkela_wire_8382)
    );

    bfr new_Jinkela_buffer_2539 (
        .din(new_Jinkela_wire_2940),
        .dout(new_Jinkela_wire_2941)
    );

    bfr new_Jinkela_buffer_6772 (
        .din(new_Jinkela_wire_8347),
        .dout(new_Jinkela_wire_8348)
    );

    bfr new_Jinkela_buffer_6795 (
        .din(n_0870_),
        .dout(new_Jinkela_wire_8392)
    );

    bfr new_Jinkela_buffer_2540 (
        .din(new_Jinkela_wire_2941),
        .dout(new_Jinkela_wire_2942)
    );

    bfr new_Jinkela_buffer_6773 (
        .din(new_Jinkela_wire_8348),
        .dout(new_Jinkela_wire_8349)
    );

    bfr new_Jinkela_buffer_2710 (
        .din(new_Jinkela_wire_3119),
        .dout(new_Jinkela_wire_3120)
    );

    bfr new_Jinkela_buffer_2589 (
        .din(new_Jinkela_wire_2994),
        .dout(new_Jinkela_wire_2995)
    );

    bfr new_Jinkela_buffer_6793 (
        .din(new_Jinkela_wire_8389),
        .dout(new_Jinkela_wire_8390)
    );

    bfr new_Jinkela_buffer_2541 (
        .din(new_Jinkela_wire_2942),
        .dout(new_Jinkela_wire_2943)
    );

    bfr new_Jinkela_buffer_6774 (
        .din(new_Jinkela_wire_8349),
        .dout(new_Jinkela_wire_8350)
    );

    bfr new_Jinkela_buffer_6791 (
        .din(new_Jinkela_wire_8385),
        .dout(new_Jinkela_wire_8386)
    );

    bfr new_Jinkela_buffer_2542 (
        .din(new_Jinkela_wire_2943),
        .dout(new_Jinkela_wire_2944)
    );

    bfr new_Jinkela_buffer_6775 (
        .din(new_Jinkela_wire_8350),
        .dout(new_Jinkela_wire_8351)
    );

    bfr new_Jinkela_buffer_2647 (
        .din(new_Jinkela_wire_3056),
        .dout(new_Jinkela_wire_3057)
    );

    bfr new_Jinkela_buffer_2590 (
        .din(new_Jinkela_wire_2995),
        .dout(new_Jinkela_wire_2996)
    );

    bfr new_Jinkela_buffer_6796 (
        .din(n_0313_),
        .dout(new_Jinkela_wire_8393)
    );

    bfr new_Jinkela_buffer_2543 (
        .din(new_Jinkela_wire_2944),
        .dout(new_Jinkela_wire_2945)
    );

    bfr new_Jinkela_buffer_6776 (
        .din(new_Jinkela_wire_8351),
        .dout(new_Jinkela_wire_8352)
    );

    spl2 new_Jinkela_splitter_635 (
        .a(new_Jinkela_wire_8386),
        .b(new_Jinkela_wire_8387),
        .c(new_Jinkela_wire_8388)
    );

    bfr new_Jinkela_buffer_2544 (
        .din(new_Jinkela_wire_2945),
        .dout(new_Jinkela_wire_2946)
    );

    bfr new_Jinkela_buffer_6777 (
        .din(new_Jinkela_wire_8352),
        .dout(new_Jinkela_wire_8353)
    );

    bfr new_Jinkela_buffer_2591 (
        .din(new_Jinkela_wire_2996),
        .dout(new_Jinkela_wire_2997)
    );

    spl3L new_Jinkela_splitter_636 (
        .a(n_1105_),
        .d(new_Jinkela_wire_8396),
        .b(new_Jinkela_wire_8397),
        .c(new_Jinkela_wire_8398)
    );

    bfr new_Jinkela_buffer_2545 (
        .din(new_Jinkela_wire_2946),
        .dout(new_Jinkela_wire_2947)
    );

    bfr new_Jinkela_buffer_6778 (
        .din(new_Jinkela_wire_8353),
        .dout(new_Jinkela_wire_8354)
    );

    bfr new_Jinkela_buffer_6794 (
        .din(new_Jinkela_wire_8390),
        .dout(new_Jinkela_wire_8391)
    );

    bfr new_Jinkela_buffer_2546 (
        .din(new_Jinkela_wire_2947),
        .dout(new_Jinkela_wire_2948)
    );

    bfr new_Jinkela_buffer_6779 (
        .din(new_Jinkela_wire_8354),
        .dout(new_Jinkela_wire_8355)
    );

    bfr new_Jinkela_buffer_2648 (
        .din(new_Jinkela_wire_3057),
        .dout(new_Jinkela_wire_3058)
    );

    bfr new_Jinkela_buffer_2592 (
        .din(new_Jinkela_wire_2997),
        .dout(new_Jinkela_wire_2998)
    );

    spl2 new_Jinkela_splitter_638 (
        .a(n_0605_),
        .b(new_Jinkela_wire_8401),
        .c(new_Jinkela_wire_8402)
    );

    bfr new_Jinkela_buffer_6797 (
        .din(new_Jinkela_wire_8393),
        .dout(new_Jinkela_wire_8394)
    );

    bfr new_Jinkela_buffer_2547 (
        .din(new_Jinkela_wire_2948),
        .dout(new_Jinkela_wire_2949)
    );

    bfr new_Jinkela_buffer_6780 (
        .din(new_Jinkela_wire_8355),
        .dout(new_Jinkela_wire_8356)
    );

    bfr new_Jinkela_buffer_6799 (
        .din(n_0398_),
        .dout(new_Jinkela_wire_8403)
    );

    bfr new_Jinkela_buffer_2548 (
        .din(new_Jinkela_wire_2949),
        .dout(new_Jinkela_wire_2950)
    );

    bfr new_Jinkela_buffer_6798 (
        .din(new_Jinkela_wire_8394),
        .dout(new_Jinkela_wire_8395)
    );

    bfr new_Jinkela_buffer_2713 (
        .din(new_Jinkela_wire_3122),
        .dout(new_Jinkela_wire_3123)
    );

    bfr new_Jinkela_buffer_2593 (
        .din(new_Jinkela_wire_2998),
        .dout(new_Jinkela_wire_2999)
    );

    bfr new_Jinkela_buffer_2549 (
        .din(new_Jinkela_wire_2950),
        .dout(new_Jinkela_wire_2951)
    );

    spl2 new_Jinkela_splitter_637 (
        .a(new_Jinkela_wire_8398),
        .b(new_Jinkela_wire_8399),
        .c(new_Jinkela_wire_8400)
    );

    bfr new_Jinkela_buffer_2776 (
        .din(new_Jinkela_wire_3190),
        .dout(new_Jinkela_wire_3191)
    );

    bfr new_Jinkela_buffer_6801 (
        .din(new_Jinkela_wire_8404),
        .dout(new_Jinkela_wire_8405)
    );

    bfr new_Jinkela_buffer_2550 (
        .din(new_Jinkela_wire_2951),
        .dout(new_Jinkela_wire_2952)
    );

    bfr new_Jinkela_buffer_6800 (
        .din(new_Jinkela_wire_8403),
        .dout(new_Jinkela_wire_8404)
    );

    bfr new_Jinkela_buffer_2649 (
        .din(new_Jinkela_wire_3058),
        .dout(new_Jinkela_wire_3059)
    );

    bfr new_Jinkela_buffer_2594 (
        .din(new_Jinkela_wire_2999),
        .dout(new_Jinkela_wire_3000)
    );

    bfr new_Jinkela_buffer_6804 (
        .din(n_0180_),
        .dout(new_Jinkela_wire_8410)
    );

    bfr new_Jinkela_buffer_2551 (
        .din(new_Jinkela_wire_2952),
        .dout(new_Jinkela_wire_2953)
    );

    spl2 new_Jinkela_splitter_642 (
        .a(n_0229_),
        .b(new_Jinkela_wire_8439),
        .c(new_Jinkela_wire_8440)
    );

    spl2 new_Jinkela_splitter_641 (
        .a(n_1221_),
        .b(new_Jinkela_wire_8437),
        .c(new_Jinkela_wire_8438)
    );

    bfr new_Jinkela_buffer_2552 (
        .din(new_Jinkela_wire_2953),
        .dout(new_Jinkela_wire_2954)
    );

    bfr new_Jinkela_buffer_6805 (
        .din(new_Jinkela_wire_8410),
        .dout(new_Jinkela_wire_8411)
    );

    bfr new_Jinkela_buffer_2712 (
        .din(new_Jinkela_wire_3121),
        .dout(new_Jinkela_wire_3122)
    );

    bfr new_Jinkela_buffer_2595 (
        .din(new_Jinkela_wire_3000),
        .dout(new_Jinkela_wire_3001)
    );

    bfr new_Jinkela_buffer_6802 (
        .din(new_Jinkela_wire_8405),
        .dout(new_Jinkela_wire_8406)
    );

    bfr new_Jinkela_buffer_2553 (
        .din(new_Jinkela_wire_2954),
        .dout(new_Jinkela_wire_2955)
    );

    bfr new_Jinkela_buffer_6829 (
        .din(n_1159_),
        .dout(new_Jinkela_wire_8443)
    );

    bfr new_Jinkela_buffer_6803 (
        .din(new_Jinkela_wire_8406),
        .dout(new_Jinkela_wire_8407)
    );

    bfr new_Jinkela_buffer_2554 (
        .din(new_Jinkela_wire_2955),
        .dout(new_Jinkela_wire_2956)
    );

    bfr new_Jinkela_buffer_6806 (
        .din(new_Jinkela_wire_8411),
        .dout(new_Jinkela_wire_8412)
    );

    bfr new_Jinkela_buffer_2650 (
        .din(new_Jinkela_wire_3059),
        .dout(new_Jinkela_wire_3060)
    );

    bfr new_Jinkela_buffer_2596 (
        .din(new_Jinkela_wire_3001),
        .dout(new_Jinkela_wire_3002)
    );

    spl2 new_Jinkela_splitter_639 (
        .a(new_Jinkela_wire_8407),
        .b(new_Jinkela_wire_8408),
        .c(new_Jinkela_wire_8409)
    );

    bfr new_Jinkela_buffer_2555 (
        .din(new_Jinkela_wire_2956),
        .dout(new_Jinkela_wire_2957)
    );

    spl2 new_Jinkela_splitter_643 (
        .a(n_0346_),
        .b(new_Jinkela_wire_8441),
        .c(new_Jinkela_wire_8442)
    );

    bfr new_Jinkela_buffer_6807 (
        .din(new_Jinkela_wire_8412),
        .dout(new_Jinkela_wire_8413)
    );

    bfr new_Jinkela_buffer_1830 (
        .din(new_Jinkela_wire_2184),
        .dout(new_Jinkela_wire_2185)
    );

    bfr new_Jinkela_buffer_398 (
        .din(new_Jinkela_wire_429),
        .dout(new_Jinkela_wire_430)
    );

    bfr new_Jinkela_buffer_7756 (
        .din(new_Jinkela_wire_9788),
        .dout(new_Jinkela_wire_9789)
    );

    bfr new_Jinkela_buffer_335 (
        .din(new_Jinkela_wire_366),
        .dout(new_Jinkela_wire_367)
    );

    bfr new_Jinkela_buffer_5128 (
        .din(new_Jinkela_wire_6119),
        .dout(new_Jinkela_wire_6120)
    );

    bfr new_Jinkela_buffer_1785 (
        .din(new_Jinkela_wire_2135),
        .dout(new_Jinkela_wire_2136)
    );

    bfr new_Jinkela_buffer_242 (
        .din(new_Jinkela_wire_261),
        .dout(new_Jinkela_wire_262)
    );

    bfr new_Jinkela_buffer_1947 (
        .din(new_Jinkela_wire_2311),
        .dout(new_Jinkela_wire_2312)
    );

    bfr new_Jinkela_buffer_278 (
        .din(new_Jinkela_wire_302),
        .dout(new_Jinkela_wire_303)
    );

    bfr new_Jinkela_buffer_5175 (
        .din(n_0325_),
        .dout(new_Jinkela_wire_6185)
    );

    bfr new_Jinkela_buffer_1886 (
        .din(new_Jinkela_wire_2246),
        .dout(new_Jinkela_wire_2247)
    );

    bfr new_Jinkela_buffer_5129 (
        .din(new_Jinkela_wire_6120),
        .dout(new_Jinkela_wire_6121)
    );

    bfr new_Jinkela_buffer_7757 (
        .din(new_Jinkela_wire_9789),
        .dout(new_Jinkela_wire_9790)
    );

    bfr new_Jinkela_buffer_1786 (
        .din(new_Jinkela_wire_2136),
        .dout(new_Jinkela_wire_2137)
    );

    bfr new_Jinkela_buffer_243 (
        .din(new_Jinkela_wire_262),
        .dout(new_Jinkela_wire_263)
    );

    bfr new_Jinkela_buffer_7803 (
        .din(new_Jinkela_wire_9837),
        .dout(new_Jinkela_wire_9838)
    );

    bfr new_Jinkela_buffer_7779 (
        .din(new_Jinkela_wire_9811),
        .dout(new_Jinkela_wire_9812)
    );

    bfr new_Jinkela_buffer_5158 (
        .din(new_Jinkela_wire_6167),
        .dout(new_Jinkela_wire_6168)
    );

    bfr new_Jinkela_buffer_1831 (
        .din(new_Jinkela_wire_2185),
        .dout(new_Jinkela_wire_2186)
    );

    bfr new_Jinkela_buffer_7758 (
        .din(new_Jinkela_wire_9790),
        .dout(new_Jinkela_wire_9791)
    );

    bfr new_Jinkela_buffer_5130 (
        .din(new_Jinkela_wire_6121),
        .dout(new_Jinkela_wire_6122)
    );

    bfr new_Jinkela_buffer_1787 (
        .din(new_Jinkela_wire_2137),
        .dout(new_Jinkela_wire_2138)
    );

    bfr new_Jinkela_buffer_244 (
        .din(new_Jinkela_wire_263),
        .dout(new_Jinkela_wire_264)
    );

    bfr new_Jinkela_buffer_5138 (
        .din(new_Jinkela_wire_6143),
        .dout(new_Jinkela_wire_6144)
    );

    bfr new_Jinkela_buffer_7759 (
        .din(new_Jinkela_wire_9791),
        .dout(new_Jinkela_wire_9792)
    );

    bfr new_Jinkela_buffer_279 (
        .din(new_Jinkela_wire_303),
        .dout(new_Jinkela_wire_304)
    );

    bfr new_Jinkela_buffer_5131 (
        .din(new_Jinkela_wire_6122),
        .dout(new_Jinkela_wire_6123)
    );

    bfr new_Jinkela_buffer_1788 (
        .din(new_Jinkela_wire_2138),
        .dout(new_Jinkela_wire_2139)
    );

    bfr new_Jinkela_buffer_245 (
        .din(new_Jinkela_wire_264),
        .dout(new_Jinkela_wire_265)
    );

    bfr new_Jinkela_buffer_5147 (
        .din(new_Jinkela_wire_6156),
        .dout(new_Jinkela_wire_6157)
    );

    bfr new_Jinkela_buffer_7780 (
        .din(new_Jinkela_wire_9812),
        .dout(new_Jinkela_wire_9813)
    );

    bfr new_Jinkela_buffer_1832 (
        .din(new_Jinkela_wire_2186),
        .dout(new_Jinkela_wire_2187)
    );

    bfr new_Jinkela_buffer_407 (
        .din(N289),
        .dout(new_Jinkela_wire_439)
    );

    bfr new_Jinkela_buffer_7760 (
        .din(new_Jinkela_wire_9792),
        .dout(new_Jinkela_wire_9793)
    );

    bfr new_Jinkela_buffer_336 (
        .din(new_Jinkela_wire_367),
        .dout(new_Jinkela_wire_368)
    );

    bfr new_Jinkela_buffer_5132 (
        .din(new_Jinkela_wire_6123),
        .dout(new_Jinkela_wire_6124)
    );

    bfr new_Jinkela_buffer_1789 (
        .din(new_Jinkela_wire_2139),
        .dout(new_Jinkela_wire_2140)
    );

    bfr new_Jinkela_buffer_246 (
        .din(new_Jinkela_wire_265),
        .dout(new_Jinkela_wire_266)
    );

    bfr new_Jinkela_buffer_5139 (
        .din(new_Jinkela_wire_6144),
        .dout(new_Jinkela_wire_6145)
    );

    bfr new_Jinkela_buffer_2011 (
        .din(new_Jinkela_wire_2375),
        .dout(new_Jinkela_wire_2376)
    );

    bfr new_Jinkela_buffer_280 (
        .din(new_Jinkela_wire_304),
        .dout(new_Jinkela_wire_305)
    );

    bfr new_Jinkela_buffer_7761 (
        .din(new_Jinkela_wire_9793),
        .dout(new_Jinkela_wire_9794)
    );

    bfr new_Jinkela_buffer_1887 (
        .din(new_Jinkela_wire_2247),
        .dout(new_Jinkela_wire_2248)
    );

    bfr new_Jinkela_buffer_5133 (
        .din(new_Jinkela_wire_6124),
        .dout(new_Jinkela_wire_6125)
    );

    bfr new_Jinkela_buffer_1790 (
        .din(new_Jinkela_wire_2140),
        .dout(new_Jinkela_wire_2141)
    );

    bfr new_Jinkela_buffer_247 (
        .din(new_Jinkela_wire_266),
        .dout(new_Jinkela_wire_267)
    );

    bfr new_Jinkela_buffer_7804 (
        .din(new_Jinkela_wire_9838),
        .dout(new_Jinkela_wire_9839)
    );

    bfr new_Jinkela_buffer_7781 (
        .din(new_Jinkela_wire_9813),
        .dout(new_Jinkela_wire_9814)
    );

    spl2 new_Jinkela_splitter_389 (
        .a(n_0924_),
        .b(new_Jinkela_wire_6188),
        .c(new_Jinkela_wire_6189)
    );

    bfr new_Jinkela_buffer_1833 (
        .din(new_Jinkela_wire_2187),
        .dout(new_Jinkela_wire_2188)
    );

    bfr new_Jinkela_buffer_7762 (
        .din(new_Jinkela_wire_9794),
        .dout(new_Jinkela_wire_9795)
    );

    bfr new_Jinkela_buffer_5134 (
        .din(new_Jinkela_wire_6125),
        .dout(new_Jinkela_wire_6126)
    );

    bfr new_Jinkela_buffer_1791 (
        .din(new_Jinkela_wire_2141),
        .dout(new_Jinkela_wire_2142)
    );

    bfr new_Jinkela_buffer_281 (
        .din(new_Jinkela_wire_305),
        .dout(new_Jinkela_wire_306)
    );

    bfr new_Jinkela_buffer_5140 (
        .din(new_Jinkela_wire_6145),
        .dout(new_Jinkela_wire_6146)
    );

    bfr new_Jinkela_buffer_7763 (
        .din(new_Jinkela_wire_9795),
        .dout(new_Jinkela_wire_9796)
    );

    bfr new_Jinkela_buffer_401 (
        .din(new_Jinkela_wire_432),
        .dout(new_Jinkela_wire_433)
    );

    bfr new_Jinkela_buffer_337 (
        .din(new_Jinkela_wire_368),
        .dout(new_Jinkela_wire_369)
    );

    bfr new_Jinkela_buffer_5135 (
        .din(new_Jinkela_wire_6126),
        .dout(new_Jinkela_wire_6127)
    );

    bfr new_Jinkela_buffer_1792 (
        .din(new_Jinkela_wire_2142),
        .dout(new_Jinkela_wire_2143)
    );

    bfr new_Jinkela_buffer_282 (
        .din(new_Jinkela_wire_306),
        .dout(new_Jinkela_wire_307)
    );

    bfr new_Jinkela_buffer_7841 (
        .din(n_0949_),
        .dout(new_Jinkela_wire_9886)
    );

    bfr new_Jinkela_buffer_5148 (
        .din(new_Jinkela_wire_6157),
        .dout(new_Jinkela_wire_6158)
    );

    bfr new_Jinkela_buffer_7782 (
        .din(new_Jinkela_wire_9814),
        .dout(new_Jinkela_wire_9815)
    );

    bfr new_Jinkela_buffer_7764 (
        .din(new_Jinkela_wire_9796),
        .dout(new_Jinkela_wire_9797)
    );

    bfr new_Jinkela_buffer_1834 (
        .din(new_Jinkela_wire_2188),
        .dout(new_Jinkela_wire_2189)
    );

    spl2 new_Jinkela_splitter_381 (
        .a(new_Jinkela_wire_6127),
        .b(new_Jinkela_wire_6128),
        .c(new_Jinkela_wire_6129)
    );

    bfr new_Jinkela_buffer_1793 (
        .din(new_Jinkela_wire_2143),
        .dout(new_Jinkela_wire_2144)
    );

    bfr new_Jinkela_buffer_283 (
        .din(new_Jinkela_wire_307),
        .dout(new_Jinkela_wire_308)
    );

    spl2 new_Jinkela_splitter_390 (
        .a(n_0815_),
        .b(new_Jinkela_wire_6190),
        .c(new_Jinkela_wire_6191)
    );

    bfr new_Jinkela_buffer_2013 (
        .din(N349),
        .dout(new_Jinkela_wire_2378)
    );

    bfr new_Jinkela_buffer_404 (
        .din(new_Jinkela_wire_435),
        .dout(new_Jinkela_wire_436)
    );

    bfr new_Jinkela_buffer_5159 (
        .din(new_Jinkela_wire_6168),
        .dout(new_Jinkela_wire_6169)
    );

    bfr new_Jinkela_buffer_338 (
        .din(new_Jinkela_wire_369),
        .dout(new_Jinkela_wire_370)
    );

    bfr new_Jinkela_buffer_1888 (
        .din(new_Jinkela_wire_2248),
        .dout(new_Jinkela_wire_2249)
    );

    bfr new_Jinkela_buffer_5141 (
        .din(new_Jinkela_wire_6146),
        .dout(new_Jinkela_wire_6147)
    );

    bfr new_Jinkela_buffer_1794 (
        .din(new_Jinkela_wire_2144),
        .dout(new_Jinkela_wire_2145)
    );

    bfr new_Jinkela_buffer_284 (
        .din(new_Jinkela_wire_308),
        .dout(new_Jinkela_wire_309)
    );

    bfr new_Jinkela_buffer_7765 (
        .din(new_Jinkela_wire_9797),
        .dout(new_Jinkela_wire_9798)
    );

    bfr new_Jinkela_buffer_5142 (
        .din(new_Jinkela_wire_6147),
        .dout(new_Jinkela_wire_6148)
    );

    bfr new_Jinkela_buffer_7783 (
        .din(new_Jinkela_wire_9815),
        .dout(new_Jinkela_wire_9816)
    );

    bfr new_Jinkela_buffer_7805 (
        .din(new_Jinkela_wire_9839),
        .dout(new_Jinkela_wire_9840)
    );

    bfr new_Jinkela_buffer_7766 (
        .din(new_Jinkela_wire_9798),
        .dout(new_Jinkela_wire_9799)
    );

    bfr new_Jinkela_buffer_1835 (
        .din(new_Jinkela_wire_2189),
        .dout(new_Jinkela_wire_2190)
    );

    bfr new_Jinkela_buffer_5149 (
        .din(new_Jinkela_wire_6158),
        .dout(new_Jinkela_wire_6159)
    );

    bfr new_Jinkela_buffer_1795 (
        .din(new_Jinkela_wire_2145),
        .dout(new_Jinkela_wire_2146)
    );

    bfr new_Jinkela_buffer_285 (
        .din(new_Jinkela_wire_309),
        .dout(new_Jinkela_wire_310)
    );

    bfr new_Jinkela_buffer_5143 (
        .din(new_Jinkela_wire_6148),
        .dout(new_Jinkela_wire_6149)
    );

    bfr new_Jinkela_buffer_7767 (
        .din(new_Jinkela_wire_9799),
        .dout(new_Jinkela_wire_9800)
    );

    bfr new_Jinkela_buffer_402 (
        .din(new_Jinkela_wire_433),
        .dout(new_Jinkela_wire_434)
    );

    bfr new_Jinkela_buffer_339 (
        .din(new_Jinkela_wire_370),
        .dout(new_Jinkela_wire_371)
    );

    bfr new_Jinkela_buffer_2077 (
        .din(N190),
        .dout(new_Jinkela_wire_2447)
    );

    bfr new_Jinkela_buffer_1796 (
        .din(new_Jinkela_wire_2146),
        .dout(new_Jinkela_wire_2147)
    );

    bfr new_Jinkela_buffer_286 (
        .din(new_Jinkela_wire_310),
        .dout(new_Jinkela_wire_311)
    );

    bfr new_Jinkela_buffer_5176 (
        .din(new_Jinkela_wire_6185),
        .dout(new_Jinkela_wire_6186)
    );

    bfr new_Jinkela_buffer_5144 (
        .din(new_Jinkela_wire_6149),
        .dout(new_Jinkela_wire_6150)
    );

    bfr new_Jinkela_buffer_7784 (
        .din(new_Jinkela_wire_9816),
        .dout(new_Jinkela_wire_9817)
    );

    bfr new_Jinkela_buffer_7842 (
        .din(n_0491_),
        .dout(new_Jinkela_wire_9887)
    );

    bfr new_Jinkela_buffer_7768 (
        .din(new_Jinkela_wire_9800),
        .dout(new_Jinkela_wire_9801)
    );

    bfr new_Jinkela_buffer_1836 (
        .din(new_Jinkela_wire_2190),
        .dout(new_Jinkela_wire_2191)
    );

    bfr new_Jinkela_buffer_5150 (
        .din(new_Jinkela_wire_6159),
        .dout(new_Jinkela_wire_6160)
    );

    bfr new_Jinkela_buffer_1797 (
        .din(new_Jinkela_wire_2147),
        .dout(new_Jinkela_wire_2148)
    );

    bfr new_Jinkela_buffer_287 (
        .din(new_Jinkela_wire_311),
        .dout(new_Jinkela_wire_312)
    );

    bfr new_Jinkela_buffer_5145 (
        .din(new_Jinkela_wire_6150),
        .dout(new_Jinkela_wire_6151)
    );

    bfr new_Jinkela_buffer_7806 (
        .din(new_Jinkela_wire_9848),
        .dout(new_Jinkela_wire_9849)
    );

    bfr new_Jinkela_buffer_7769 (
        .din(new_Jinkela_wire_9801),
        .dout(new_Jinkela_wire_9802)
    );

    bfr new_Jinkela_buffer_1948 (
        .din(new_Jinkela_wire_2312),
        .dout(new_Jinkela_wire_2313)
    );

    bfr new_Jinkela_buffer_340 (
        .din(new_Jinkela_wire_371),
        .dout(new_Jinkela_wire_372)
    );

    bfr new_Jinkela_buffer_1889 (
        .din(new_Jinkela_wire_2249),
        .dout(new_Jinkela_wire_2250)
    );

    bfr new_Jinkela_buffer_1798 (
        .din(new_Jinkela_wire_2148),
        .dout(new_Jinkela_wire_2149)
    );

    bfr new_Jinkela_buffer_288 (
        .din(new_Jinkela_wire_312),
        .dout(new_Jinkela_wire_313)
    );

    bfr new_Jinkela_buffer_5160 (
        .din(new_Jinkela_wire_6169),
        .dout(new_Jinkela_wire_6170)
    );

    bfr new_Jinkela_buffer_5151 (
        .din(new_Jinkela_wire_6160),
        .dout(new_Jinkela_wire_6161)
    );

    bfr new_Jinkela_buffer_7785 (
        .din(new_Jinkela_wire_9817),
        .dout(new_Jinkela_wire_9818)
    );

    spl2 new_Jinkela_splitter_816 (
        .a(new_Jinkela_wire_9840),
        .b(new_Jinkela_wire_9841),
        .c(new_Jinkela_wire_9842)
    );

    bfr new_Jinkela_buffer_7770 (
        .din(new_Jinkela_wire_9802),
        .dout(new_Jinkela_wire_9803)
    );

    bfr new_Jinkela_buffer_1837 (
        .din(new_Jinkela_wire_2191),
        .dout(new_Jinkela_wire_2192)
    );

    bfr new_Jinkela_buffer_543 (
        .din(N133),
        .dout(new_Jinkela_wire_585)
    );

    spl2 new_Jinkela_splitter_394 (
        .a(n_1048_),
        .b(new_Jinkela_wire_6245),
        .c(new_Jinkela_wire_6246)
    );

    bfr new_Jinkela_buffer_289 (
        .din(new_Jinkela_wire_313),
        .dout(new_Jinkela_wire_314)
    );

    bfr new_Jinkela_buffer_5152 (
        .din(new_Jinkela_wire_6161),
        .dout(new_Jinkela_wire_6162)
    );

    bfr new_Jinkela_buffer_1838 (
        .din(new_Jinkela_wire_2192),
        .dout(new_Jinkela_wire_2193)
    );

    bfr new_Jinkela_buffer_405 (
        .din(new_Jinkela_wire_436),
        .dout(new_Jinkela_wire_437)
    );

    bfr new_Jinkela_buffer_7864 (
        .din(n_0048_),
        .dout(new_Jinkela_wire_9914)
    );

    bfr new_Jinkela_buffer_341 (
        .din(new_Jinkela_wire_372),
        .dout(new_Jinkela_wire_373)
    );

    bfr new_Jinkela_buffer_7786 (
        .din(new_Jinkela_wire_9818),
        .dout(new_Jinkela_wire_9819)
    );

    bfr new_Jinkela_buffer_2012 (
        .din(new_Jinkela_wire_2376),
        .dout(new_Jinkela_wire_2377)
    );

    bfr new_Jinkela_buffer_290 (
        .din(new_Jinkela_wire_314),
        .dout(new_Jinkela_wire_315)
    );

    bfr new_Jinkela_buffer_5161 (
        .din(new_Jinkela_wire_6170),
        .dout(new_Jinkela_wire_6171)
    );

    bfr new_Jinkela_buffer_1890 (
        .din(new_Jinkela_wire_2250),
        .dout(new_Jinkela_wire_2251)
    );

    bfr new_Jinkela_buffer_5153 (
        .din(new_Jinkela_wire_6162),
        .dout(new_Jinkela_wire_6163)
    );

    bfr new_Jinkela_buffer_7807 (
        .din(new_Jinkela_wire_9849),
        .dout(new_Jinkela_wire_9850)
    );

    spl3L new_Jinkela_splitter_822 (
        .a(n_1319_),
        .d(new_Jinkela_wire_9893),
        .b(new_Jinkela_wire_9894),
        .c(new_Jinkela_wire_9895)
    );

    bfr new_Jinkela_buffer_1839 (
        .din(new_Jinkela_wire_2193),
        .dout(new_Jinkela_wire_2194)
    );

    bfr new_Jinkela_buffer_7787 (
        .din(new_Jinkela_wire_9819),
        .dout(new_Jinkela_wire_9820)
    );

    bfr new_Jinkela_buffer_5177 (
        .din(new_Jinkela_wire_6186),
        .dout(new_Jinkela_wire_6187)
    );

    bfr new_Jinkela_buffer_291 (
        .din(new_Jinkela_wire_315),
        .dout(new_Jinkela_wire_316)
    );

    bfr new_Jinkela_buffer_5154 (
        .din(new_Jinkela_wire_6163),
        .dout(new_Jinkela_wire_6164)
    );

    spl4L new_Jinkela_splitter_824 (
        .a(n_0860_),
        .d(new_Jinkela_wire_9921),
        .b(new_Jinkela_wire_9922),
        .e(new_Jinkela_wire_9923),
        .c(new_Jinkela_wire_9924)
    );

    bfr new_Jinkela_buffer_1840 (
        .din(new_Jinkela_wire_2194),
        .dout(new_Jinkela_wire_2195)
    );

    bfr new_Jinkela_buffer_471 (
        .din(N69),
        .dout(new_Jinkela_wire_508)
    );

    bfr new_Jinkela_buffer_342 (
        .din(new_Jinkela_wire_373),
        .dout(new_Jinkela_wire_374)
    );

    bfr new_Jinkela_buffer_7788 (
        .din(new_Jinkela_wire_9820),
        .dout(new_Jinkela_wire_9821)
    );

    bfr new_Jinkela_buffer_1949 (
        .din(new_Jinkela_wire_2313),
        .dout(new_Jinkela_wire_2314)
    );

    bfr new_Jinkela_buffer_292 (
        .din(new_Jinkela_wire_316),
        .dout(new_Jinkela_wire_317)
    );

    bfr new_Jinkela_buffer_5162 (
        .din(new_Jinkela_wire_6171),
        .dout(new_Jinkela_wire_6172)
    );

    bfr new_Jinkela_buffer_1891 (
        .din(new_Jinkela_wire_2251),
        .dout(new_Jinkela_wire_2252)
    );

    bfr new_Jinkela_buffer_5155 (
        .din(new_Jinkela_wire_6164),
        .dout(new_Jinkela_wire_6165)
    );

    bfr new_Jinkela_buffer_7843 (
        .din(new_Jinkela_wire_9887),
        .dout(new_Jinkela_wire_9888)
    );

    bfr new_Jinkela_buffer_1841 (
        .din(new_Jinkela_wire_2195),
        .dout(new_Jinkela_wire_2196)
    );

    bfr new_Jinkela_buffer_7789 (
        .din(new_Jinkela_wire_9821),
        .dout(new_Jinkela_wire_9822)
    );

    bfr new_Jinkela_buffer_293 (
        .din(new_Jinkela_wire_317),
        .dout(new_Jinkela_wire_318)
    );

    bfr new_Jinkela_buffer_5156 (
        .din(new_Jinkela_wire_6165),
        .dout(new_Jinkela_wire_6166)
    );

    bfr new_Jinkela_buffer_7808 (
        .din(new_Jinkela_wire_9850),
        .dout(new_Jinkela_wire_9851)
    );

    bfr new_Jinkela_buffer_1842 (
        .din(new_Jinkela_wire_2196),
        .dout(new_Jinkela_wire_2197)
    );

    bfr new_Jinkela_buffer_406 (
        .din(new_Jinkela_wire_437),
        .dout(new_Jinkela_wire_438)
    );

    bfr new_Jinkela_buffer_343 (
        .din(new_Jinkela_wire_374),
        .dout(new_Jinkela_wire_375)
    );

    bfr new_Jinkela_buffer_7790 (
        .din(new_Jinkela_wire_9822),
        .dout(new_Jinkela_wire_9823)
    );

    bfr new_Jinkela_buffer_5163 (
        .din(new_Jinkela_wire_6172),
        .dout(new_Jinkela_wire_6173)
    );

    bfr new_Jinkela_buffer_294 (
        .din(new_Jinkela_wire_318),
        .dout(new_Jinkela_wire_319)
    );

    bfr new_Jinkela_buffer_1892 (
        .din(new_Jinkela_wire_2252),
        .dout(new_Jinkela_wire_2253)
    );

    spl2 new_Jinkela_splitter_391 (
        .a(n_0108_),
        .b(new_Jinkela_wire_6192),
        .c(new_Jinkela_wire_6195)
    );

    bfr new_Jinkela_buffer_1843 (
        .din(new_Jinkela_wire_2197),
        .dout(new_Jinkela_wire_2198)
    );

    bfr new_Jinkela_buffer_5216 (
        .din(new_net_2537),
        .dout(new_Jinkela_wire_6238)
    );

    bfr new_Jinkela_buffer_7791 (
        .din(new_Jinkela_wire_9823),
        .dout(new_Jinkela_wire_9824)
    );

    bfr new_Jinkela_buffer_5164 (
        .din(new_Jinkela_wire_6173),
        .dout(new_Jinkela_wire_6174)
    );

    bfr new_Jinkela_buffer_295 (
        .din(new_Jinkela_wire_319),
        .dout(new_Jinkela_wire_320)
    );

    bfr new_Jinkela_buffer_7809 (
        .din(new_Jinkela_wire_9851),
        .dout(new_Jinkela_wire_9852)
    );

    and_bi n_2706_ (
        .a(new_Jinkela_wire_10146),
        .b(new_Jinkela_wire_7225),
        .c(n_0563_)
    );

    or_bb n_2707_ (
        .a(n_0563_),
        .b(new_Jinkela_wire_8757),
        .c(n_0564_)
    );

    and_ii n_2708_ (
        .a(new_Jinkela_wire_8880),
        .b(new_Jinkela_wire_3699),
        .c(n_0565_)
    );

    and_bb n_2709_ (
        .a(new_Jinkela_wire_8879),
        .b(new_Jinkela_wire_3698),
        .c(n_0566_)
    );

    and_ii n_2710_ (
        .a(n_0566_),
        .b(n_0565_),
        .c(n_0567_)
    );

    or_bb n_2711_ (
        .a(new_Jinkela_wire_8314),
        .b(new_Jinkela_wire_6133),
        .c(n_0568_)
    );

    and_bb n_2712_ (
        .a(new_Jinkela_wire_8313),
        .b(new_Jinkela_wire_6132),
        .c(n_0569_)
    );

    or_bi n_2713_ (
        .a(n_0569_),
        .b(n_0568_),
        .c(n_0570_)
    );

    and_bi n_2714_ (
        .a(new_Jinkela_wire_9015),
        .b(new_Jinkela_wire_9429),
        .c(n_0571_)
    );

    and_ii n_2715_ (
        .a(n_0571_),
        .b(n_0558_),
        .c(n_0572_)
    );

    and_ii n_2716_ (
        .a(new_Jinkela_wire_5980),
        .b(new_Jinkela_wire_8624),
        .c(n_0573_)
    );

    or_bi n_2717_ (
        .a(new_Jinkela_wire_3718),
        .b(new_Jinkela_wire_4435),
        .c(n_0574_)
    );

    and_bb n_2718_ (
        .a(new_Jinkela_wire_7405),
        .b(new_Jinkela_wire_8926),
        .c(n_0575_)
    );

    and_ii n_2719_ (
        .a(new_Jinkela_wire_7404),
        .b(new_Jinkela_wire_8925),
        .c(n_0576_)
    );

    and_ii n_2720_ (
        .a(n_0576_),
        .b(n_0575_),
        .c(n_0577_)
    );

    and_ii n_2721_ (
        .a(new_Jinkela_wire_7188),
        .b(new_Jinkela_wire_7252),
        .c(n_0578_)
    );

    and_bb n_2722_ (
        .a(new_Jinkela_wire_7187),
        .b(new_Jinkela_wire_7251),
        .c(n_0579_)
    );

    or_bb n_2723_ (
        .a(n_0579_),
        .b(n_0578_),
        .c(new_net_2539)
    );

    and_ii n_2724_ (
        .a(new_Jinkela_wire_9351),
        .b(new_Jinkela_wire_8514),
        .c(n_0580_)
    );

    and_bi n_2725_ (
        .a(new_Jinkela_wire_9345),
        .b(new_Jinkela_wire_8844),
        .c(n_0581_)
    );

    and_ii n_2726_ (
        .a(new_Jinkela_wire_9609),
        .b(n_0580_),
        .c(n_0582_)
    );

    and_ii n_2727_ (
        .a(new_Jinkela_wire_9484),
        .b(new_Jinkela_wire_6137),
        .c(n_0583_)
    );

    and_bb n_2728_ (
        .a(new_Jinkela_wire_9483),
        .b(new_Jinkela_wire_6138),
        .c(n_0584_)
    );

    or_bb n_2729_ (
        .a(n_0584_),
        .b(n_0583_),
        .c(n_0585_)
    );

    and_ii n_2730_ (
        .a(new_Jinkela_wire_6745),
        .b(new_Jinkela_wire_5879),
        .c(n_0586_)
    );

    and_bi n_2731_ (
        .a(new_Jinkela_wire_4523),
        .b(new_Jinkela_wire_10341),
        .c(n_0587_)
    );

    or_bb n_2732_ (
        .a(new_Jinkela_wire_3912),
        .b(new_Jinkela_wire_10508),
        .c(n_0588_)
    );

    and_bi n_2733_ (
        .a(new_Jinkela_wire_3911),
        .b(new_Jinkela_wire_9623),
        .c(n_0589_)
    );

    and_bi n_2734_ (
        .a(n_0588_),
        .b(n_0589_),
        .c(n_0590_)
    );

    and_ii n_2735_ (
        .a(new_Jinkela_wire_6946),
        .b(new_Jinkela_wire_8884),
        .c(n_0591_)
    );

    and_bb n_2736_ (
        .a(new_Jinkela_wire_6945),
        .b(new_Jinkela_wire_8883),
        .c(n_0592_)
    );

    and_ii n_2737_ (
        .a(n_0592_),
        .b(n_0591_),
        .c(n_0593_)
    );

    or_bb n_2738_ (
        .a(new_Jinkela_wire_9769),
        .b(new_Jinkela_wire_4917),
        .c(n_0594_)
    );

    and_bi n_2739_ (
        .a(new_Jinkela_wire_5089),
        .b(new_Jinkela_wire_6407),
        .c(n_0595_)
    );

    and_bi n_2740_ (
        .a(new_Jinkela_wire_6406),
        .b(new_Jinkela_wire_8847),
        .c(n_0596_)
    );

    or_bb n_2741_ (
        .a(n_0596_),
        .b(n_0595_),
        .c(n_0597_)
    );

    or_bi n_2742_ (
        .a(new_Jinkela_wire_8849),
        .b(new_Jinkela_wire_3729),
        .c(n_0598_)
    );

    and_bi n_2743_ (
        .a(new_Jinkela_wire_6135),
        .b(new_Jinkela_wire_8511),
        .c(n_0599_)
    );

    and_bb n_2744_ (
        .a(new_Jinkela_wire_8509),
        .b(new_Jinkela_wire_7205),
        .c(n_0600_)
    );

    and_bi n_2745_ (
        .a(new_Jinkela_wire_3822),
        .b(new_Jinkela_wire_6141),
        .c(n_0601_)
    );

    and_ii n_2746_ (
        .a(n_0601_),
        .b(new_Jinkela_wire_4970),
        .c(n_0602_)
    );

    and_ii n_2747_ (
        .a(new_Jinkela_wire_8176),
        .b(new_Jinkela_wire_3920),
        .c(n_0603_)
    );

    bfr new_Jinkela_buffer_5941 (
        .din(new_Jinkela_wire_7180),
        .dout(new_Jinkela_wire_7181)
    );

    bfr new_Jinkela_buffer_4300 (
        .din(new_Jinkela_wire_5082),
        .dout(new_Jinkela_wire_5083)
    );

    and_ii n_1989_ (
        .a(new_Jinkela_wire_9641),
        .b(new_Jinkela_wire_7370),
        .c(n_1255_)
    );

    bfr new_Jinkela_buffer_4277 (
        .din(new_Jinkela_wire_5045),
        .dout(new_Jinkela_wire_5046)
    );

    bfr new_Jinkela_buffer_7792 (
        .din(new_Jinkela_wire_9824),
        .dout(new_Jinkela_wire_9825)
    );

    spl4L new_Jinkela_splitter_502 (
        .a(n_1178_),
        .d(new_Jinkela_wire_7276),
        .b(new_Jinkela_wire_7277),
        .e(new_Jinkela_wire_7278),
        .c(new_Jinkela_wire_7279)
    );

    and_ii n_1990_ (
        .a(new_Jinkela_wire_7272),
        .b(new_Jinkela_wire_5641),
        .c(n_1256_)
    );

    spl2 new_Jinkela_splitter_501 (
        .a(n_0803_),
        .b(new_Jinkela_wire_7274),
        .c(new_Jinkela_wire_7275)
    );

    bfr new_Jinkela_buffer_7844 (
        .din(new_Jinkela_wire_9888),
        .dout(new_Jinkela_wire_9889)
    );

    bfr new_Jinkela_buffer_5942 (
        .din(new_Jinkela_wire_7181),
        .dout(new_Jinkela_wire_7182)
    );

    and_bb n_1991_ (
        .a(new_Jinkela_wire_7270),
        .b(new_Jinkela_wire_5642),
        .c(n_1257_)
    );

    bfr new_Jinkela_buffer_4278 (
        .din(new_Jinkela_wire_5046),
        .dout(new_Jinkela_wire_5047)
    );

    bfr new_Jinkela_buffer_7793 (
        .din(new_Jinkela_wire_9825),
        .dout(new_Jinkela_wire_9826)
    );

    bfr new_Jinkela_buffer_5989 (
        .din(new_Jinkela_wire_7256),
        .dout(new_Jinkela_wire_7257)
    );

    and_ii n_1992_ (
        .a(n_1257_),
        .b(n_1256_),
        .c(n_1258_)
    );

    spl2 new_Jinkela_splitter_302 (
        .a(n_0726_),
        .b(new_Jinkela_wire_5146),
        .c(new_Jinkela_wire_5147)
    );

    bfr new_Jinkela_buffer_7810 (
        .din(new_Jinkela_wire_9852),
        .dout(new_Jinkela_wire_9853)
    );

    bfr new_Jinkela_buffer_5943 (
        .din(new_Jinkela_wire_7182),
        .dout(new_Jinkela_wire_7183)
    );

    bfr new_Jinkela_buffer_4301 (
        .din(new_Jinkela_wire_5083),
        .dout(new_Jinkela_wire_5084)
    );

    and_bb n_1993_ (
        .a(new_Jinkela_wire_779),
        .b(new_Jinkela_wire_1186),
        .c(n_1259_)
    );

    bfr new_Jinkela_buffer_4279 (
        .din(new_Jinkela_wire_5047),
        .dout(new_Jinkela_wire_5048)
    );

    bfr new_Jinkela_buffer_7794 (
        .din(new_Jinkela_wire_9826),
        .dout(new_Jinkela_wire_9827)
    );

    and_ii n_1994_ (
        .a(new_Jinkela_wire_9983),
        .b(new_Jinkela_wire_6152),
        .c(n_1260_)
    );

    bfr new_Jinkela_buffer_5994 (
        .din(n_0415_),
        .dout(new_Jinkela_wire_7280)
    );

    bfr new_Jinkela_buffer_5944 (
        .din(new_Jinkela_wire_7183),
        .dout(new_Jinkela_wire_7184)
    );

    and_bb n_1995_ (
        .a(new_Jinkela_wire_3048),
        .b(new_Jinkela_wire_1215),
        .c(n_1261_)
    );

    bfr new_Jinkela_buffer_4280 (
        .din(new_Jinkela_wire_5048),
        .dout(new_Jinkela_wire_5049)
    );

    bfr new_Jinkela_buffer_7795 (
        .din(new_Jinkela_wire_9827),
        .dout(new_Jinkela_wire_9828)
    );

    bfr new_Jinkela_buffer_5990 (
        .din(new_Jinkela_wire_7257),
        .dout(new_Jinkela_wire_7258)
    );

    and_ii n_1996_ (
        .a(new_Jinkela_wire_5094),
        .b(new_Jinkela_wire_4187),
        .c(n_1262_)
    );

    spl3L new_Jinkela_splitter_301 (
        .a(n_0076_),
        .d(new_Jinkela_wire_5143),
        .b(new_Jinkela_wire_5144),
        .c(new_Jinkela_wire_5145)
    );

    bfr new_Jinkela_buffer_7811 (
        .din(new_Jinkela_wire_9853),
        .dout(new_Jinkela_wire_9854)
    );

    bfr new_Jinkela_buffer_4302 (
        .din(new_Jinkela_wire_5084),
        .dout(new_Jinkela_wire_5085)
    );

    and_bi n_1997_ (
        .a(new_Jinkela_wire_10421),
        .b(new_Jinkela_wire_3868),
        .c(n_1263_)
    );

    bfr new_Jinkela_buffer_4281 (
        .din(new_Jinkela_wire_5049),
        .dout(new_Jinkela_wire_5050)
    );

    bfr new_Jinkela_buffer_5995 (
        .din(new_Jinkela_wire_7280),
        .dout(new_Jinkela_wire_7281)
    );

    bfr new_Jinkela_buffer_7796 (
        .din(new_Jinkela_wire_9828),
        .dout(new_Jinkela_wire_9829)
    );

    bfr new_Jinkela_buffer_5991 (
        .din(new_Jinkela_wire_7258),
        .dout(new_Jinkela_wire_7259)
    );

    and_bi n_1998_ (
        .a(new_Jinkela_wire_3869),
        .b(new_Jinkela_wire_10420),
        .c(n_1264_)
    );

    bfr new_Jinkela_buffer_7845 (
        .din(new_Jinkela_wire_9889),
        .dout(new_Jinkela_wire_9890)
    );

    bfr new_Jinkela_buffer_4308 (
        .din(new_Jinkela_wire_5108),
        .dout(new_Jinkela_wire_5109)
    );

    and_ii n_1999_ (
        .a(n_1264_),
        .b(n_1263_),
        .c(n_1265_)
    );

    bfr new_Jinkela_buffer_4282 (
        .din(new_Jinkela_wire_5050),
        .dout(new_Jinkela_wire_5051)
    );

    bfr new_Jinkela_buffer_7797 (
        .din(new_Jinkela_wire_9829),
        .dout(new_Jinkela_wire_9830)
    );

    bfr new_Jinkela_buffer_5992 (
        .din(new_Jinkela_wire_7259),
        .dout(new_Jinkela_wire_7260)
    );

    and_bi n_2000_ (
        .a(new_Jinkela_wire_8477),
        .b(new_Jinkela_wire_9643),
        .c(n_1266_)
    );

    bfr new_Jinkela_buffer_4307 (
        .din(new_Jinkela_wire_5104),
        .dout(new_Jinkela_wire_5105)
    );

    bfr new_Jinkela_buffer_7812 (
        .din(new_Jinkela_wire_9854),
        .dout(new_Jinkela_wire_9855)
    );

    bfr new_Jinkela_buffer_4303 (
        .din(new_Jinkela_wire_5085),
        .dout(new_Jinkela_wire_5086)
    );

    and_bi n_2001_ (
        .a(new_Jinkela_wire_9642),
        .b(new_Jinkela_wire_8476),
        .c(n_1267_)
    );

    bfr new_Jinkela_buffer_4283 (
        .din(new_Jinkela_wire_5051),
        .dout(new_Jinkela_wire_5052)
    );

    spl2 new_Jinkela_splitter_504 (
        .a(n_1173_),
        .b(new_Jinkela_wire_7297),
        .c(new_Jinkela_wire_7298)
    );

    bfr new_Jinkela_buffer_7798 (
        .din(new_Jinkela_wire_9830),
        .dout(new_Jinkela_wire_9831)
    );

    bfr new_Jinkela_buffer_5993 (
        .din(new_Jinkela_wire_7260),
        .dout(new_Jinkela_wire_7261)
    );

    and_ii n_2002_ (
        .a(n_1267_),
        .b(n_1266_),
        .c(n_1268_)
    );

    bfr new_Jinkela_buffer_7846 (
        .din(new_Jinkela_wire_9895),
        .dout(new_Jinkela_wire_9896)
    );

    and_ii n_2003_ (
        .a(new_Jinkela_wire_8886),
        .b(new_Jinkela_wire_7351),
        .c(n_1269_)
    );

    bfr new_Jinkela_buffer_4284 (
        .din(new_Jinkela_wire_5052),
        .dout(new_Jinkela_wire_5053)
    );

    spl2 new_Jinkela_splitter_503 (
        .a(n_1081_),
        .b(new_Jinkela_wire_7295),
        .c(new_Jinkela_wire_7296)
    );

    bfr new_Jinkela_buffer_7813 (
        .din(new_Jinkela_wire_9855),
        .dout(new_Jinkela_wire_9856)
    );

    and_bb n_2004_ (
        .a(new_Jinkela_wire_8885),
        .b(new_Jinkela_wire_7350),
        .c(n_1270_)
    );

    spl2 new_Jinkela_splitter_303 (
        .a(n_0938_),
        .b(new_Jinkela_wire_5150),
        .c(new_Jinkela_wire_5151)
    );

    spl2 new_Jinkela_splitter_506 (
        .a(n_0403_),
        .b(new_Jinkela_wire_7301),
        .c(new_Jinkela_wire_7302)
    );

    spl2 new_Jinkela_splitter_821 (
        .a(new_Jinkela_wire_9890),
        .b(new_Jinkela_wire_9891),
        .c(new_Jinkela_wire_9892)
    );

    bfr new_Jinkela_buffer_5996 (
        .din(new_Jinkela_wire_7281),
        .dout(new_Jinkela_wire_7282)
    );

    bfr new_Jinkela_buffer_7869 (
        .din(n_0212_),
        .dout(new_Jinkela_wire_9925)
    );

    and_ii n_2005_ (
        .a(n_1270_),
        .b(n_1269_),
        .c(n_1271_)
    );

    bfr new_Jinkela_buffer_7814 (
        .din(new_Jinkela_wire_9856),
        .dout(new_Jinkela_wire_9857)
    );

    and_bb n_2006_ (
        .a(new_Jinkela_wire_2080),
        .b(new_Jinkela_wire_1199),
        .c(n_1272_)
    );

    bfr new_Jinkela_buffer_4309 (
        .din(new_Jinkela_wire_5109),
        .dout(new_Jinkela_wire_5110)
    );

    bfr new_Jinkela_buffer_7865 (
        .din(new_Jinkela_wire_9914),
        .dout(new_Jinkela_wire_9915)
    );

    bfr new_Jinkela_buffer_5997 (
        .din(new_Jinkela_wire_7282),
        .dout(new_Jinkela_wire_7283)
    );

    and_ii n_2007_ (
        .a(new_Jinkela_wire_8180),
        .b(new_Jinkela_wire_7274),
        .c(n_1273_)
    );

    bfr new_Jinkela_buffer_7815 (
        .din(new_Jinkela_wire_9857),
        .dout(new_Jinkela_wire_9858)
    );

    spl2 new_Jinkela_splitter_505 (
        .a(n_0033_),
        .b(new_Jinkela_wire_7299),
        .c(new_Jinkela_wire_7300)
    );

    bfr new_Jinkela_buffer_4348 (
        .din(n_1157_),
        .dout(new_Jinkela_wire_5156)
    );

    and_bb n_2008_ (
        .a(new_Jinkela_wire_2555),
        .b(new_Jinkela_wire_1341),
        .c(n_1274_)
    );

    bfr new_Jinkela_buffer_4310 (
        .din(new_Jinkela_wire_5110),
        .dout(new_Jinkela_wire_5111)
    );

    spl2 new_Jinkela_splitter_508 (
        .a(n_0806_),
        .b(new_Jinkela_wire_7305),
        .c(new_Jinkela_wire_7306)
    );

    bfr new_Jinkela_buffer_7847 (
        .din(new_Jinkela_wire_9896),
        .dout(new_Jinkela_wire_9897)
    );

    bfr new_Jinkela_buffer_5998 (
        .din(new_Jinkela_wire_7283),
        .dout(new_Jinkela_wire_7284)
    );

    and_ii n_2009_ (
        .a(new_Jinkela_wire_5054),
        .b(new_Jinkela_wire_7081),
        .c(n_1275_)
    );

    bfr new_Jinkela_buffer_4342 (
        .din(new_Jinkela_wire_5147),
        .dout(new_Jinkela_wire_5148)
    );

    bfr new_Jinkela_buffer_7816 (
        .din(new_Jinkela_wire_9858),
        .dout(new_Jinkela_wire_9859)
    );

    and_bi n_2010_ (
        .a(new_Jinkela_wire_8292),
        .b(new_Jinkela_wire_3696),
        .c(n_1276_)
    );

    bfr new_Jinkela_buffer_4311 (
        .din(new_Jinkela_wire_5111),
        .dout(new_Jinkela_wire_5112)
    );

    bfr new_Jinkela_buffer_7848 (
        .din(new_Jinkela_wire_9897),
        .dout(new_Jinkela_wire_9898)
    );

    bfr new_Jinkela_buffer_5999 (
        .din(new_Jinkela_wire_7284),
        .dout(new_Jinkela_wire_7285)
    );

    and_bi n_2011_ (
        .a(new_Jinkela_wire_3697),
        .b(new_Jinkela_wire_8290),
        .c(n_1277_)
    );

    bfr new_Jinkela_buffer_7817 (
        .din(new_Jinkela_wire_9859),
        .dout(new_Jinkela_wire_9860)
    );

    spl2 new_Jinkela_splitter_507 (
        .a(n_0088_),
        .b(new_Jinkela_wire_7303),
        .c(new_Jinkela_wire_7304)
    );

    and_ii n_2012_ (
        .a(n_1277_),
        .b(n_1276_),
        .c(n_1278_)
    );

    bfr new_Jinkela_buffer_4312 (
        .din(new_Jinkela_wire_5112),
        .dout(new_Jinkela_wire_5113)
    );

    bfr new_Jinkela_buffer_6000 (
        .din(new_Jinkela_wire_7285),
        .dout(new_Jinkela_wire_7286)
    );

    and_bb n_2013_ (
        .a(new_Jinkela_wire_1981),
        .b(new_Jinkela_wire_1297),
        .c(n_1279_)
    );

    bfr new_Jinkela_buffer_4343 (
        .din(new_Jinkela_wire_5148),
        .dout(new_Jinkela_wire_5149)
    );

    bfr new_Jinkela_buffer_7818 (
        .din(new_Jinkela_wire_9860),
        .dout(new_Jinkela_wire_9861)
    );

    and_ii n_2014_ (
        .a(new_Jinkela_wire_9956),
        .b(new_Jinkela_wire_10360),
        .c(n_1280_)
    );

    bfr new_Jinkela_buffer_4313 (
        .din(new_Jinkela_wire_5113),
        .dout(new_Jinkela_wire_5114)
    );

    spl2 new_Jinkela_splitter_825 (
        .a(n_1320_),
        .b(new_Jinkela_wire_9926),
        .c(new_Jinkela_wire_9928)
    );

    bfr new_Jinkela_buffer_7849 (
        .din(new_Jinkela_wire_9898),
        .dout(new_Jinkela_wire_9899)
    );

    bfr new_Jinkela_buffer_6001 (
        .din(new_Jinkela_wire_7286),
        .dout(new_Jinkela_wire_7287)
    );

    and_bb n_2015_ (
        .a(new_Jinkela_wire_1690),
        .b(new_Jinkela_wire_1278),
        .c(n_1281_)
    );

    bfr new_Jinkela_buffer_4344 (
        .din(new_Jinkela_wire_5151),
        .dout(new_Jinkela_wire_5152)
    );

    bfr new_Jinkela_buffer_7819 (
        .din(new_Jinkela_wire_9861),
        .dout(new_Jinkela_wire_9862)
    );

    spl3L new_Jinkela_splitter_509 (
        .a(n_1124_),
        .d(new_Jinkela_wire_7307),
        .b(new_Jinkela_wire_7308),
        .c(new_Jinkela_wire_7309)
    );

    spl4L new_Jinkela_splitter_304 (
        .a(n_0758_),
        .d(new_Jinkela_wire_5157),
        .b(new_Jinkela_wire_5158),
        .e(new_Jinkela_wire_5159),
        .c(new_Jinkela_wire_5160)
    );

    and_ii n_2016_ (
        .a(new_Jinkela_wire_5298),
        .b(new_Jinkela_wire_9392),
        .c(n_1282_)
    );

    bfr new_Jinkela_buffer_4314 (
        .din(new_Jinkela_wire_5114),
        .dout(new_Jinkela_wire_5115)
    );

    spl3L new_Jinkela_splitter_512 (
        .a(n_0701_),
        .d(new_Jinkela_wire_7322),
        .b(new_Jinkela_wire_7323),
        .c(new_Jinkela_wire_7324)
    );

    bfr new_Jinkela_buffer_7866 (
        .din(new_Jinkela_wire_9915),
        .dout(new_Jinkela_wire_9916)
    );

    bfr new_Jinkela_buffer_6002 (
        .din(new_Jinkela_wire_7287),
        .dout(new_Jinkela_wire_7288)
    );

    and_ii n_2017_ (
        .a(new_Jinkela_wire_8576),
        .b(new_Jinkela_wire_10099),
        .c(n_1283_)
    );

    spl3L new_Jinkela_splitter_305 (
        .a(n_0012_),
        .d(new_Jinkela_wire_5161),
        .b(new_Jinkela_wire_5162),
        .c(new_Jinkela_wire_5163)
    );

    bfr new_Jinkela_buffer_7820 (
        .din(new_Jinkela_wire_9862),
        .dout(new_Jinkela_wire_9863)
    );

    bfr new_Jinkela_buffer_6009 (
        .din(n_1339_),
        .dout(new_Jinkela_wire_7310)
    );

    and_bb n_2018_ (
        .a(new_Jinkela_wire_8575),
        .b(new_Jinkela_wire_10097),
        .c(n_1284_)
    );

    bfr new_Jinkela_buffer_4315 (
        .din(new_Jinkela_wire_5115),
        .dout(new_Jinkela_wire_5116)
    );

    bfr new_Jinkela_buffer_7850 (
        .din(new_Jinkela_wire_9899),
        .dout(new_Jinkela_wire_9900)
    );

    bfr new_Jinkela_buffer_6003 (
        .din(new_Jinkela_wire_7288),
        .dout(new_Jinkela_wire_7289)
    );

    and_ii n_2019_ (
        .a(n_1284_),
        .b(n_1283_),
        .c(n_1285_)
    );

    bfr new_Jinkela_buffer_4345 (
        .din(new_Jinkela_wire_5152),
        .dout(new_Jinkela_wire_5153)
    );

    bfr new_Jinkela_buffer_7821 (
        .din(new_Jinkela_wire_9863),
        .dout(new_Jinkela_wire_9864)
    );

    bfr new_Jinkela_buffer_6010 (
        .din(new_Jinkela_wire_7310),
        .dout(new_Jinkela_wire_7311)
    );

    and_bi n_2020_ (
        .a(new_Jinkela_wire_8092),
        .b(new_Jinkela_wire_3732),
        .c(n_1286_)
    );

    bfr new_Jinkela_buffer_4316 (
        .din(new_Jinkela_wire_5116),
        .dout(new_Jinkela_wire_5117)
    );

    spl2 new_Jinkela_splitter_514 (
        .a(n_1212_),
        .b(new_Jinkela_wire_7330),
        .c(new_Jinkela_wire_7331)
    );

    bfr new_Jinkela_buffer_7893 (
        .din(n_1225_),
        .dout(new_Jinkela_wire_9955)
    );

    bfr new_Jinkela_buffer_6004 (
        .din(new_Jinkela_wire_7289),
        .dout(new_Jinkela_wire_7290)
    );

    and_bi n_2021_ (
        .a(new_Jinkela_wire_3731),
        .b(new_Jinkela_wire_8091),
        .c(n_1287_)
    );

    bfr new_Jinkela_buffer_4349 (
        .din(n_0262_),
        .dout(new_Jinkela_wire_5164)
    );

    bfr new_Jinkela_buffer_7822 (
        .din(new_Jinkela_wire_9864),
        .dout(new_Jinkela_wire_9865)
    );

    bfr new_Jinkela_buffer_4350 (
        .din(new_Jinkela_wire_5164),
        .dout(new_Jinkela_wire_5165)
    );

    and_ii n_2022_ (
        .a(n_1287_),
        .b(n_1286_),
        .c(n_1288_)
    );

    bfr new_Jinkela_buffer_4317 (
        .din(new_Jinkela_wire_5117),
        .dout(new_Jinkela_wire_5118)
    );

    bfr new_Jinkela_buffer_7851 (
        .din(new_Jinkela_wire_9900),
        .dout(new_Jinkela_wire_9901)
    );

    bfr new_Jinkela_buffer_6005 (
        .din(new_Jinkela_wire_7290),
        .dout(new_Jinkela_wire_7291)
    );

    and_bb n_2023_ (
        .a(new_Jinkela_wire_9117),
        .b(new_Jinkela_wire_8324),
        .c(n_1289_)
    );

    bfr new_Jinkela_buffer_4346 (
        .din(new_Jinkela_wire_5153),
        .dout(new_Jinkela_wire_5154)
    );

    bfr new_Jinkela_buffer_7823 (
        .din(new_Jinkela_wire_9865),
        .dout(new_Jinkela_wire_9866)
    );

    bfr new_Jinkela_buffer_6017 (
        .din(new_Jinkela_wire_7324),
        .dout(new_Jinkela_wire_7325)
    );

    and_ii n_2024_ (
        .a(new_Jinkela_wire_9116),
        .b(new_Jinkela_wire_8323),
        .c(n_1290_)
    );

    bfr new_Jinkela_buffer_4318 (
        .din(new_Jinkela_wire_5118),
        .dout(new_Jinkela_wire_5119)
    );

    bfr new_Jinkela_buffer_7867 (
        .din(new_Jinkela_wire_9916),
        .dout(new_Jinkela_wire_9917)
    );

    bfr new_Jinkela_buffer_6006 (
        .din(new_Jinkela_wire_7291),
        .dout(new_Jinkela_wire_7292)
    );

    or_bb n_2025_ (
        .a(n_1290_),
        .b(n_1289_),
        .c(n_1291_)
    );

    bfr new_Jinkela_buffer_4377 (
        .din(n_0668_),
        .dout(new_Jinkela_wire_5197)
    );

    bfr new_Jinkela_buffer_7824 (
        .din(new_Jinkela_wire_9866),
        .dout(new_Jinkela_wire_9867)
    );

    bfr new_Jinkela_buffer_6011 (
        .din(new_Jinkela_wire_7311),
        .dout(new_Jinkela_wire_7312)
    );

    or_bb n_2026_ (
        .a(n_1291_),
        .b(n_1244_),
        .c(n_1292_)
    );

    bfr new_Jinkela_buffer_4319 (
        .din(new_Jinkela_wire_5119),
        .dout(new_Jinkela_wire_5120)
    );

    bfr new_Jinkela_buffer_7852 (
        .din(new_Jinkela_wire_9901),
        .dout(new_Jinkela_wire_9902)
    );

    bfr new_Jinkela_buffer_6007 (
        .din(new_Jinkela_wire_7292),
        .dout(new_Jinkela_wire_7293)
    );

    or_bb n_2027_ (
        .a(n_1292_),
        .b(n_1197_),
        .c(new_net_5)
    );

    bfr new_Jinkela_buffer_4347 (
        .din(new_Jinkela_wire_5154),
        .dout(new_Jinkela_wire_5155)
    );

    bfr new_Jinkela_buffer_7825 (
        .din(new_Jinkela_wire_9867),
        .dout(new_Jinkela_wire_9868)
    );

    spl4L new_Jinkela_splitter_513 (
        .a(n_1226_),
        .d(new_Jinkela_wire_7326),
        .b(new_Jinkela_wire_7327),
        .e(new_Jinkela_wire_7328),
        .c(new_Jinkela_wire_7329)
    );

    inv n_2028_ (
        .din(new_Jinkela_wire_2591),
        .dout(n_1293_)
    );

    bfr new_Jinkela_buffer_4320 (
        .din(new_Jinkela_wire_5120),
        .dout(new_Jinkela_wire_5121)
    );

    spl4L new_Jinkela_splitter_826 (
        .a(new_Jinkela_wire_9928),
        .d(new_Jinkela_wire_9929),
        .b(new_Jinkela_wire_9930),
        .e(new_Jinkela_wire_9931),
        .c(new_Jinkela_wire_9932)
    );

    bfr new_Jinkela_buffer_6008 (
        .din(new_Jinkela_wire_7293),
        .dout(new_Jinkela_wire_7294)
    );

    and_bi n_2029_ (
        .a(new_Jinkela_wire_8704),
        .b(new_Jinkela_wire_5058),
        .c(n_1294_)
    );

    bfr new_Jinkela_buffer_7826 (
        .din(new_Jinkela_wire_9868),
        .dout(new_Jinkela_wire_9869)
    );

    bfr new_Jinkela_buffer_6012 (
        .din(new_Jinkela_wire_7312),
        .dout(new_Jinkela_wire_7313)
    );

    spl3L new_Jinkela_splitter_306 (
        .a(n_0385_),
        .d(new_Jinkela_wire_5166),
        .b(new_Jinkela_wire_5167),
        .c(new_Jinkela_wire_5168)
    );

    and_bi n_2030_ (
        .a(new_Jinkela_wire_5056),
        .b(new_Jinkela_wire_8703),
        .c(n_1295_)
    );

    bfr new_Jinkela_buffer_4321 (
        .din(new_Jinkela_wire_5121),
        .dout(new_Jinkela_wire_5122)
    );

    bfr new_Jinkela_buffer_3432 (
        .din(new_Jinkela_wire_3993),
        .dout(new_Jinkela_wire_3994)
    );

    bfr new_Jinkela_buffer_2556 (
        .din(new_Jinkela_wire_2957),
        .dout(new_Jinkela_wire_2958)
    );

    bfr new_Jinkela_buffer_3480 (
        .din(new_Jinkela_wire_4056),
        .dout(new_Jinkela_wire_4057)
    );

    bfr new_Jinkela_buffer_2597 (
        .din(new_Jinkela_wire_3002),
        .dout(new_Jinkela_wire_3003)
    );

    bfr new_Jinkela_buffer_3462 (
        .din(new_Jinkela_wire_4034),
        .dout(new_Jinkela_wire_4035)
    );

    bfr new_Jinkela_buffer_3433 (
        .din(new_Jinkela_wire_3994),
        .dout(new_Jinkela_wire_3995)
    );

    bfr new_Jinkela_buffer_2557 (
        .din(new_Jinkela_wire_2958),
        .dout(new_Jinkela_wire_2959)
    );

    spl2 new_Jinkela_splitter_138 (
        .a(new_Jinkela_wire_3123),
        .b(new_Jinkela_wire_3124),
        .c(new_Jinkela_wire_3125)
    );

    bfr new_Jinkela_buffer_3434 (
        .din(new_Jinkela_wire_3995),
        .dout(new_Jinkela_wire_3996)
    );

    bfr new_Jinkela_buffer_2558 (
        .din(new_Jinkela_wire_2959),
        .dout(new_Jinkela_wire_2960)
    );

    bfr new_Jinkela_buffer_3573 (
        .din(n_0625_),
        .dout(new_Jinkela_wire_4171)
    );

    bfr new_Jinkela_buffer_2651 (
        .din(new_Jinkela_wire_3060),
        .dout(new_Jinkela_wire_3061)
    );

    bfr new_Jinkela_buffer_2598 (
        .din(new_Jinkela_wire_3003),
        .dout(new_Jinkela_wire_3004)
    );

    bfr new_Jinkela_buffer_3463 (
        .din(new_Jinkela_wire_4035),
        .dout(new_Jinkela_wire_4036)
    );

    bfr new_Jinkela_buffer_3435 (
        .din(new_Jinkela_wire_3996),
        .dout(new_Jinkela_wire_3997)
    );

    bfr new_Jinkela_buffer_2559 (
        .din(new_Jinkela_wire_2960),
        .dout(new_Jinkela_wire_2961)
    );

    bfr new_Jinkela_buffer_3495 (
        .din(new_Jinkela_wire_4073),
        .dout(new_Jinkela_wire_4074)
    );

    bfr new_Jinkela_buffer_3436 (
        .din(new_Jinkela_wire_3997),
        .dout(new_Jinkela_wire_3998)
    );

    bfr new_Jinkela_buffer_2560 (
        .din(new_Jinkela_wire_2961),
        .dout(new_Jinkela_wire_2962)
    );

    bfr new_Jinkela_buffer_3481 (
        .din(new_Jinkela_wire_4057),
        .dout(new_Jinkela_wire_4058)
    );

    bfr new_Jinkela_buffer_2714 (
        .din(new_Jinkela_wire_3125),
        .dout(new_Jinkela_wire_3126)
    );

    bfr new_Jinkela_buffer_2599 (
        .din(new_Jinkela_wire_3004),
        .dout(new_Jinkela_wire_3005)
    );

    bfr new_Jinkela_buffer_3464 (
        .din(new_Jinkela_wire_4036),
        .dout(new_Jinkela_wire_4037)
    );

    bfr new_Jinkela_buffer_3437 (
        .din(new_Jinkela_wire_3998),
        .dout(new_Jinkela_wire_3999)
    );

    bfr new_Jinkela_buffer_2561 (
        .din(new_Jinkela_wire_2962),
        .dout(new_Jinkela_wire_2963)
    );

    bfr new_Jinkela_buffer_3438 (
        .din(new_Jinkela_wire_3999),
        .dout(new_Jinkela_wire_4000)
    );

    bfr new_Jinkela_buffer_2562 (
        .din(new_Jinkela_wire_2963),
        .dout(new_Jinkela_wire_2964)
    );

    bfr new_Jinkela_buffer_2652 (
        .din(new_Jinkela_wire_3061),
        .dout(new_Jinkela_wire_3062)
    );

    bfr new_Jinkela_buffer_2600 (
        .din(new_Jinkela_wire_3005),
        .dout(new_Jinkela_wire_3006)
    );

    bfr new_Jinkela_buffer_3465 (
        .din(new_Jinkela_wire_4037),
        .dout(new_Jinkela_wire_4038)
    );

    bfr new_Jinkela_buffer_7014 (
        .din(new_Jinkela_wire_8666),
        .dout(new_Jinkela_wire_8667)
    );

    bfr new_Jinkela_buffer_3439 (
        .din(new_Jinkela_wire_4000),
        .dout(new_Jinkela_wire_4001)
    );

    bfr new_Jinkela_buffer_2563 (
        .din(new_Jinkela_wire_2964),
        .dout(new_Jinkela_wire_2965)
    );

    bfr new_Jinkela_buffer_3440 (
        .din(new_Jinkela_wire_4001),
        .dout(new_Jinkela_wire_4002)
    );

    bfr new_Jinkela_buffer_2564 (
        .din(new_Jinkela_wire_2965),
        .dout(new_Jinkela_wire_2966)
    );

    bfr new_Jinkela_buffer_3482 (
        .din(new_Jinkela_wire_4058),
        .dout(new_Jinkela_wire_4059)
    );

    bfr new_Jinkela_buffer_2783 (
        .din(N56),
        .dout(new_Jinkela_wire_3198)
    );

    bfr new_Jinkela_buffer_2601 (
        .din(new_Jinkela_wire_3006),
        .dout(new_Jinkela_wire_3007)
    );

    bfr new_Jinkela_buffer_3466 (
        .din(new_Jinkela_wire_4038),
        .dout(new_Jinkela_wire_4039)
    );

    bfr new_Jinkela_buffer_3441 (
        .din(new_Jinkela_wire_4002),
        .dout(new_Jinkela_wire_4003)
    );

    bfr new_Jinkela_buffer_2565 (
        .din(new_Jinkela_wire_2966),
        .dout(new_Jinkela_wire_2967)
    );

    bfr new_Jinkela_buffer_3442 (
        .din(new_Jinkela_wire_4003),
        .dout(new_Jinkela_wire_4004)
    );

    bfr new_Jinkela_buffer_2653 (
        .din(new_Jinkela_wire_3062),
        .dout(new_Jinkela_wire_3063)
    );

    bfr new_Jinkela_buffer_2602 (
        .din(new_Jinkela_wire_3007),
        .dout(new_Jinkela_wire_3008)
    );

    bfr new_Jinkela_buffer_3497 (
        .din(new_Jinkela_wire_4083),
        .dout(new_Jinkela_wire_4084)
    );

    bfr new_Jinkela_buffer_3467 (
        .din(new_Jinkela_wire_4039),
        .dout(new_Jinkela_wire_4040)
    );

    bfr new_Jinkela_buffer_3443 (
        .din(new_Jinkela_wire_4004),
        .dout(new_Jinkela_wire_4005)
    );

    bfr new_Jinkela_buffer_2777 (
        .din(new_Jinkela_wire_3191),
        .dout(new_Jinkela_wire_3192)
    );

    bfr new_Jinkela_buffer_2603 (
        .din(new_Jinkela_wire_3008),
        .dout(new_Jinkela_wire_3009)
    );

    bfr new_Jinkela_buffer_3496 (
        .din(new_Jinkela_wire_4074),
        .dout(new_Jinkela_wire_4075)
    );

    bfr new_Jinkela_buffer_3444 (
        .din(new_Jinkela_wire_4005),
        .dout(new_Jinkela_wire_4006)
    );

    bfr new_Jinkela_buffer_2654 (
        .din(new_Jinkela_wire_3063),
        .dout(new_Jinkela_wire_3064)
    );

    bfr new_Jinkela_buffer_2604 (
        .din(new_Jinkela_wire_3009),
        .dout(new_Jinkela_wire_3010)
    );

    bfr new_Jinkela_buffer_3483 (
        .din(new_Jinkela_wire_4059),
        .dout(new_Jinkela_wire_4060)
    );

    bfr new_Jinkela_buffer_3468 (
        .din(new_Jinkela_wire_4040),
        .dout(new_Jinkela_wire_4041)
    );

    bfr new_Jinkela_buffer_2780 (
        .din(new_Jinkela_wire_3194),
        .dout(new_Jinkela_wire_3195)
    );

    bfr new_Jinkela_buffer_2605 (
        .din(new_Jinkela_wire_3010),
        .dout(new_Jinkela_wire_3011)
    );

    bfr new_Jinkela_buffer_3469 (
        .din(new_Jinkela_wire_4041),
        .dout(new_Jinkela_wire_4042)
    );

    bfr new_Jinkela_buffer_2655 (
        .din(new_Jinkela_wire_3064),
        .dout(new_Jinkela_wire_3065)
    );

    bfr new_Jinkela_buffer_2606 (
        .din(new_Jinkela_wire_3011),
        .dout(new_Jinkela_wire_3012)
    );

    bfr new_Jinkela_buffer_3484 (
        .din(new_Jinkela_wire_4060),
        .dout(new_Jinkela_wire_4061)
    );

    bfr new_Jinkela_buffer_3470 (
        .din(new_Jinkela_wire_4042),
        .dout(new_Jinkela_wire_4043)
    );

    bfr new_Jinkela_buffer_2715 (
        .din(new_Jinkela_wire_3126),
        .dout(new_Jinkela_wire_3127)
    );

    bfr new_Jinkela_buffer_2607 (
        .din(new_Jinkela_wire_3012),
        .dout(new_Jinkela_wire_3013)
    );

    bfr new_Jinkela_buffer_3523 (
        .din(new_net_2507),
        .dout(new_Jinkela_wire_4121)
    );

    bfr new_Jinkela_buffer_3471 (
        .din(new_Jinkela_wire_4043),
        .dout(new_Jinkela_wire_4044)
    );

    bfr new_Jinkela_buffer_2656 (
        .din(new_Jinkela_wire_3065),
        .dout(new_Jinkela_wire_3066)
    );

    bfr new_Jinkela_buffer_2608 (
        .din(new_Jinkela_wire_3013),
        .dout(new_Jinkela_wire_3014)
    );

    spl2 new_Jinkela_splitter_207 (
        .a(new_Jinkela_wire_4075),
        .b(new_Jinkela_wire_4076),
        .c(new_Jinkela_wire_4077)
    );

    bfr new_Jinkela_buffer_3485 (
        .din(new_Jinkela_wire_4061),
        .dout(new_Jinkela_wire_4062)
    );

    bfr new_Jinkela_buffer_2778 (
        .din(new_Jinkela_wire_3192),
        .dout(new_Jinkela_wire_3193)
    );

    bfr new_Jinkela_buffer_2609 (
        .din(new_Jinkela_wire_3014),
        .dout(new_Jinkela_wire_3015)
    );

    bfr new_Jinkela_buffer_3486 (
        .din(new_Jinkela_wire_4062),
        .dout(new_Jinkela_wire_4063)
    );

    bfr new_Jinkela_buffer_3524 (
        .din(new_Jinkela_wire_4121),
        .dout(new_Jinkela_wire_4122)
    );

    bfr new_Jinkela_buffer_2657 (
        .din(new_Jinkela_wire_3066),
        .dout(new_Jinkela_wire_3067)
    );

    bfr new_Jinkela_buffer_2610 (
        .din(new_Jinkela_wire_3015),
        .dout(new_Jinkela_wire_3016)
    );

    bfr new_Jinkela_buffer_3487 (
        .din(new_Jinkela_wire_4063),
        .dout(new_Jinkela_wire_4064)
    );

    bfr new_Jinkela_buffer_2716 (
        .din(new_Jinkela_wire_3127),
        .dout(new_Jinkela_wire_3128)
    );

    bfr new_Jinkela_buffer_2611 (
        .din(new_Jinkela_wire_3016),
        .dout(new_Jinkela_wire_3017)
    );

    bfr new_Jinkela_buffer_3488 (
        .din(new_Jinkela_wire_4064),
        .dout(new_Jinkela_wire_4065)
    );

    bfr new_Jinkela_buffer_3498 (
        .din(new_Jinkela_wire_4090),
        .dout(new_Jinkela_wire_4091)
    );

    bfr new_Jinkela_buffer_2658 (
        .din(new_Jinkela_wire_3067),
        .dout(new_Jinkela_wire_3068)
    );

    bfr new_Jinkela_buffer_2612 (
        .din(new_Jinkela_wire_3017),
        .dout(new_Jinkela_wire_3018)
    );

    bfr new_Jinkela_buffer_3489 (
        .din(new_Jinkela_wire_4065),
        .dout(new_Jinkela_wire_4066)
    );

    bfr new_Jinkela_buffer_344 (
        .din(new_Jinkela_wire_375),
        .dout(new_Jinkela_wire_376)
    );

    bfr new_Jinkela_buffer_296 (
        .din(new_Jinkela_wire_320),
        .dout(new_Jinkela_wire_321)
    );

    bfr new_Jinkela_buffer_297 (
        .din(new_Jinkela_wire_321),
        .dout(new_Jinkela_wire_322)
    );

    bfr new_Jinkela_buffer_409 (
        .din(new_Jinkela_wire_440),
        .dout(new_Jinkela_wire_441)
    );

    bfr new_Jinkela_buffer_345 (
        .din(new_Jinkela_wire_376),
        .dout(new_Jinkela_wire_377)
    );

    bfr new_Jinkela_buffer_298 (
        .din(new_Jinkela_wire_322),
        .dout(new_Jinkela_wire_323)
    );

    bfr new_Jinkela_buffer_472 (
        .din(new_Jinkela_wire_508),
        .dout(new_Jinkela_wire_509)
    );

    bfr new_Jinkela_buffer_299 (
        .din(new_Jinkela_wire_323),
        .dout(new_Jinkela_wire_324)
    );

    bfr new_Jinkela_buffer_408 (
        .din(new_Jinkela_wire_439),
        .dout(new_Jinkela_wire_440)
    );

    bfr new_Jinkela_buffer_346 (
        .din(new_Jinkela_wire_377),
        .dout(new_Jinkela_wire_378)
    );

    bfr new_Jinkela_buffer_300 (
        .din(new_Jinkela_wire_324),
        .dout(new_Jinkela_wire_325)
    );

    bfr new_Jinkela_buffer_539 (
        .din(N44),
        .dout(new_Jinkela_wire_581)
    );

    bfr new_Jinkela_buffer_301 (
        .din(new_Jinkela_wire_325),
        .dout(new_Jinkela_wire_326)
    );

    bfr new_Jinkela_buffer_347 (
        .din(new_Jinkela_wire_378),
        .dout(new_Jinkela_wire_379)
    );

    bfr new_Jinkela_buffer_302 (
        .din(new_Jinkela_wire_326),
        .dout(new_Jinkela_wire_327)
    );

    bfr new_Jinkela_buffer_303 (
        .din(new_Jinkela_wire_327),
        .dout(new_Jinkela_wire_328)
    );

    spl2 new_Jinkela_splitter_14 (
        .a(new_Jinkela_wire_441),
        .b(new_Jinkela_wire_442),
        .c(new_Jinkela_wire_443)
    );

    bfr new_Jinkela_buffer_348 (
        .din(new_Jinkela_wire_379),
        .dout(new_Jinkela_wire_380)
    );

    bfr new_Jinkela_buffer_304 (
        .din(new_Jinkela_wire_328),
        .dout(new_Jinkela_wire_329)
    );

    bfr new_Jinkela_buffer_475 (
        .din(N352),
        .dout(new_Jinkela_wire_512)
    );

    bfr new_Jinkela_buffer_305 (
        .din(new_Jinkela_wire_329),
        .dout(new_Jinkela_wire_330)
    );

    bfr new_Jinkela_buffer_410 (
        .din(new_Jinkela_wire_443),
        .dout(new_Jinkela_wire_444)
    );

    bfr new_Jinkela_buffer_349 (
        .din(new_Jinkela_wire_380),
        .dout(new_Jinkela_wire_381)
    );

    bfr new_Jinkela_buffer_306 (
        .din(new_Jinkela_wire_330),
        .dout(new_Jinkela_wire_331)
    );

    bfr new_Jinkela_buffer_307 (
        .din(new_Jinkela_wire_331),
        .dout(new_Jinkela_wire_332)
    );

    bfr new_Jinkela_buffer_473 (
        .din(new_Jinkela_wire_509),
        .dout(new_Jinkela_wire_510)
    );

    bfr new_Jinkela_buffer_350 (
        .din(new_Jinkela_wire_381),
        .dout(new_Jinkela_wire_382)
    );

    bfr new_Jinkela_buffer_308 (
        .din(new_Jinkela_wire_332),
        .dout(new_Jinkela_wire_333)
    );

    bfr new_Jinkela_buffer_309 (
        .din(new_Jinkela_wire_333),
        .dout(new_Jinkela_wire_334)
    );

    bfr new_Jinkela_buffer_351 (
        .din(new_Jinkela_wire_382),
        .dout(new_Jinkela_wire_383)
    );

    bfr new_Jinkela_buffer_310 (
        .din(new_Jinkela_wire_334),
        .dout(new_Jinkela_wire_335)
    );

    bfr new_Jinkela_buffer_311 (
        .din(new_Jinkela_wire_335),
        .dout(new_Jinkela_wire_336)
    );

    bfr new_Jinkela_buffer_411 (
        .din(new_Jinkela_wire_444),
        .dout(new_Jinkela_wire_445)
    );

    bfr new_Jinkela_buffer_352 (
        .din(new_Jinkela_wire_383),
        .dout(new_Jinkela_wire_384)
    );

    bfr new_Jinkela_buffer_312 (
        .din(new_Jinkela_wire_336),
        .dout(new_Jinkela_wire_337)
    );

    bfr new_Jinkela_buffer_313 (
        .din(new_Jinkela_wire_337),
        .dout(new_Jinkela_wire_338)
    );

    bfr new_Jinkela_buffer_474 (
        .din(new_Jinkela_wire_510),
        .dout(new_Jinkela_wire_511)
    );

    bfr new_Jinkela_buffer_353 (
        .din(new_Jinkela_wire_384),
        .dout(new_Jinkela_wire_385)
    );

    bfr new_Jinkela_buffer_314 (
        .din(new_Jinkela_wire_338),
        .dout(new_Jinkela_wire_339)
    );

    bfr new_Jinkela_buffer_315 (
        .din(new_Jinkela_wire_339),
        .dout(new_Jinkela_wire_340)
    );

    or_bb n_2589_ (
        .a(n_0447_),
        .b(n_0446_),
        .c(n_0448_)
    );

    and_bi n_1418_ (
        .a(new_Jinkela_wire_2745),
        .b(new_Jinkela_wire_7266),
        .c(n_0690_)
    );

    spl3L new_Jinkela_splitter_15 (
        .a(new_Jinkela_wire_445),
        .d(new_Jinkela_wire_446),
        .b(new_Jinkela_wire_447),
        .c(new_Jinkela_wire_448)
    );

    bfr new_Jinkela_buffer_354 (
        .din(new_Jinkela_wire_385),
        .dout(new_Jinkela_wire_386)
    );

    bfr new_Jinkela_buffer_1844 (
        .din(new_Jinkela_wire_2198),
        .dout(new_Jinkela_wire_2199)
    );

    bfr new_Jinkela_buffer_1950 (
        .din(new_Jinkela_wire_2314),
        .dout(new_Jinkela_wire_2315)
    );

    bfr new_Jinkela_buffer_1893 (
        .din(new_Jinkela_wire_2253),
        .dout(new_Jinkela_wire_2254)
    );

    bfr new_Jinkela_buffer_1845 (
        .din(new_Jinkela_wire_2199),
        .dout(new_Jinkela_wire_2200)
    );

    bfr new_Jinkela_buffer_1846 (
        .din(new_Jinkela_wire_2200),
        .dout(new_Jinkela_wire_2201)
    );

    bfr new_Jinkela_buffer_1894 (
        .din(new_Jinkela_wire_2254),
        .dout(new_Jinkela_wire_2255)
    );

    bfr new_Jinkela_buffer_1847 (
        .din(new_Jinkela_wire_2201),
        .dout(new_Jinkela_wire_2202)
    );

    bfr new_Jinkela_buffer_2015 (
        .din(new_Jinkela_wire_2379),
        .dout(new_Jinkela_wire_2380)
    );

    bfr new_Jinkela_buffer_1848 (
        .din(new_Jinkela_wire_2202),
        .dout(new_Jinkela_wire_2203)
    );

    bfr new_Jinkela_buffer_1951 (
        .din(new_Jinkela_wire_2315),
        .dout(new_Jinkela_wire_2316)
    );

    bfr new_Jinkela_buffer_1895 (
        .din(new_Jinkela_wire_2255),
        .dout(new_Jinkela_wire_2256)
    );

    bfr new_Jinkela_buffer_1849 (
        .din(new_Jinkela_wire_2203),
        .dout(new_Jinkela_wire_2204)
    );

    bfr new_Jinkela_buffer_1850 (
        .din(new_Jinkela_wire_2204),
        .dout(new_Jinkela_wire_2205)
    );

    bfr new_Jinkela_buffer_2078 (
        .din(new_Jinkela_wire_2447),
        .dout(new_Jinkela_wire_2448)
    );

    bfr new_Jinkela_buffer_1896 (
        .din(new_Jinkela_wire_2256),
        .dout(new_Jinkela_wire_2257)
    );

    bfr new_Jinkela_buffer_1851 (
        .din(new_Jinkela_wire_2205),
        .dout(new_Jinkela_wire_2206)
    );

    bfr new_Jinkela_buffer_1852 (
        .din(new_Jinkela_wire_2206),
        .dout(new_Jinkela_wire_2207)
    );

    and_bi n_1397_ (
        .a(new_Jinkela_wire_8934),
        .b(new_Jinkela_wire_7931),
        .c(new_net_2531)
    );

    bfr new_Jinkela_buffer_1952 (
        .din(new_Jinkela_wire_2316),
        .dout(new_Jinkela_wire_2317)
    );

    bfr new_Jinkela_buffer_1897 (
        .din(new_Jinkela_wire_2257),
        .dout(new_Jinkela_wire_2258)
    );

    or_bb n_1375_ (
        .a(n_0654_),
        .b(n_0653_),
        .c(new_net_1)
    );

    bfr new_Jinkela_buffer_1853 (
        .din(new_Jinkela_wire_2207),
        .dout(new_Jinkela_wire_2208)
    );

    or_ii n_1373_ (
        .a(N184),
        .b(N150),
        .c(n_0653_)
    );

    or_ii n_1374_ (
        .a(N240),
        .b(N228),
        .c(n_0654_)
    );

    bfr new_Jinkela_buffer_1854 (
        .din(new_Jinkela_wire_2208),
        .dout(new_Jinkela_wire_2209)
    );

    or_bb n_1372_ (
        .a(new_Jinkela_wire_3538),
        .b(new_Jinkela_wire_96),
        .c(new_net_2562)
    );

    or_ii n_1376_ (
        .a(N152),
        .b(N210),
        .c(n_0655_)
    );

    bfr new_Jinkela_buffer_1898 (
        .din(new_Jinkela_wire_2258),
        .dout(new_Jinkela_wire_2259)
    );

    or_ii n_1380_ (
        .a(N186),
        .b(N185),
        .c(n_0658_)
    );

    bfr new_Jinkela_buffer_1855 (
        .din(new_Jinkela_wire_2209),
        .dout(new_Jinkela_wire_2210)
    );

    or_ii n_1379_ (
        .a(N182),
        .b(N183),
        .c(n_0657_)
    );

    spl2 new_Jinkela_splitter_119 (
        .a(new_Jinkela_wire_2380),
        .b(new_Jinkela_wire_2381),
        .c(new_Jinkela_wire_2382)
    );

    or_ii n_1377_ (
        .a(N230),
        .b(N218),
        .c(n_0656_)
    );

    bfr new_Jinkela_buffer_1856 (
        .din(new_Jinkela_wire_2210),
        .dout(new_Jinkela_wire_2211)
    );

    bfr new_Jinkela_buffer_1953 (
        .din(new_Jinkela_wire_2317),
        .dout(new_Jinkela_wire_2318)
    );

    or_bi n_1389_ (
        .a(new_Jinkela_wire_1312),
        .b(new_Jinkela_wire_181),
        .c(n_0662_)
    );

    bfr new_Jinkela_buffer_1899 (
        .din(new_Jinkela_wire_2259),
        .dout(new_Jinkela_wire_2260)
    );

    or_bb n_1378_ (
        .a(n_0656_),
        .b(n_0655_),
        .c(new_net_0)
    );

    bfr new_Jinkela_buffer_1857 (
        .din(new_Jinkela_wire_2211),
        .dout(new_Jinkela_wire_2212)
    );

    or_bb n_1381_ (
        .a(n_0658_),
        .b(n_0657_),
        .c(new_net_3)
    );

    or_ii n_1382_ (
        .a(N172),
        .b(N162),
        .c(n_0659_)
    );

    bfr new_Jinkela_buffer_1858 (
        .din(new_Jinkela_wire_2212),
        .dout(new_Jinkela_wire_2213)
    );

    or_ii n_1383_ (
        .a(N199),
        .b(N188),
        .c(n_0660_)
    );

    bfr new_Jinkela_buffer_2016 (
        .din(new_Jinkela_wire_2382),
        .dout(new_Jinkela_wire_2383)
    );

    or_bb n_1384_ (
        .a(n_0660_),
        .b(n_0659_),
        .c(new_net_2)
    );

    bfr new_Jinkela_buffer_1900 (
        .din(new_Jinkela_wire_2260),
        .dout(new_Jinkela_wire_2261)
    );

    bfr new_Jinkela_buffer_1859 (
        .din(new_Jinkela_wire_2213),
        .dout(new_Jinkela_wire_2214)
    );

    or_bi n_1385_ (
        .a(new_Jinkela_wire_3536),
        .b(new_Jinkela_wire_609),
        .c(new_net_10)
    );

    inv n_1386_ (
        .din(N15),
        .dout(new_net_11)
    );

    bfr new_Jinkela_buffer_1860 (
        .din(new_Jinkela_wire_2214),
        .dout(new_Jinkela_wire_2215)
    );

    and_bi n_1387_ (
        .a(new_Jinkela_wire_1609),
        .b(new_Jinkela_wire_3537),
        .c(n_0661_)
    );

    bfr new_Jinkela_buffer_1954 (
        .din(new_Jinkela_wire_2318),
        .dout(new_Jinkela_wire_2319)
    );

    or_ii n_1388_ (
        .a(n_0661_),
        .b(new_Jinkela_wire_586),
        .c(new_net_12)
    );

    bfr new_Jinkela_buffer_1901 (
        .din(new_Jinkela_wire_2261),
        .dout(new_Jinkela_wire_2262)
    );

    bfr new_Jinkela_buffer_1861 (
        .din(new_Jinkela_wire_2215),
        .dout(new_Jinkela_wire_2216)
    );

    or_bb n_1390_ (
        .a(new_Jinkela_wire_8364),
        .b(new_Jinkela_wire_2244),
        .c(n_0663_)
    );

    or_bb n_1391_ (
        .a(new_Jinkela_wire_180),
        .b(new_Jinkela_wire_1187),
        .c(n_0664_)
    );

    bfr new_Jinkela_buffer_1862 (
        .din(new_Jinkela_wire_2216),
        .dout(new_Jinkela_wire_2217)
    );

    and_bi n_1392_ (
        .a(new_Jinkela_wire_2242),
        .b(n_0664_),
        .c(n_0665_)
    );

    bfr new_Jinkela_buffer_2085 (
        .din(N47),
        .dout(new_Jinkela_wire_2455)
    );

    bfr new_Jinkela_buffer_1902 (
        .din(new_Jinkela_wire_2262),
        .dout(new_Jinkela_wire_2263)
    );

    or_bi n_1393_ (
        .a(new_Jinkela_wire_5450),
        .b(new_Jinkela_wire_3921),
        .c(n_0666_)
    );

    bfr new_Jinkela_buffer_1863 (
        .din(new_Jinkela_wire_2217),
        .dout(new_Jinkela_wire_2218)
    );

    and_bi n_1394_ (
        .a(new_Jinkela_wire_2566),
        .b(new_Jinkela_wire_6100),
        .c(n_0667_)
    );

    inv n_1395_ (
        .din(new_Jinkela_wire_2556),
        .dout(n_0668_)
    );

    bfr new_Jinkela_buffer_1864 (
        .din(new_Jinkela_wire_2218),
        .dout(new_Jinkela_wire_2219)
    );

    or_ii n_1396_ (
        .a(new_Jinkela_wire_6099),
        .b(new_Jinkela_wire_5204),
        .c(n_0669_)
    );

    bfr new_Jinkela_buffer_1955 (
        .din(new_Jinkela_wire_2319),
        .dout(new_Jinkela_wire_2320)
    );

    bfr new_Jinkela_buffer_1903 (
        .din(new_Jinkela_wire_2263),
        .dout(new_Jinkela_wire_2264)
    );

    bfr new_Jinkela_buffer_5223 (
        .din(n_0303_),
        .dout(new_Jinkela_wire_6247)
    );

    bfr new_Jinkela_buffer_7853 (
        .din(new_Jinkela_wire_9902),
        .dout(new_Jinkela_wire_9903)
    );

    bfr new_Jinkela_buffer_7827 (
        .din(new_Jinkela_wire_9869),
        .dout(new_Jinkela_wire_9870)
    );

    bfr new_Jinkela_buffer_5165 (
        .din(new_Jinkela_wire_6174),
        .dout(new_Jinkela_wire_6175)
    );

    bfr new_Jinkela_buffer_7868 (
        .din(new_Jinkela_wire_9917),
        .dout(new_Jinkela_wire_9918)
    );

    spl4L new_Jinkela_splitter_393 (
        .a(new_Jinkela_wire_6195),
        .d(new_Jinkela_wire_6196),
        .b(new_Jinkela_wire_6197),
        .e(new_Jinkela_wire_6198),
        .c(new_Jinkela_wire_6199)
    );

    bfr new_Jinkela_buffer_7828 (
        .din(new_Jinkela_wire_9870),
        .dout(new_Jinkela_wire_9871)
    );

    bfr new_Jinkela_buffer_5166 (
        .din(new_Jinkela_wire_6175),
        .dout(new_Jinkela_wire_6176)
    );

    spl2 new_Jinkela_splitter_392 (
        .a(new_Jinkela_wire_6192),
        .b(new_Jinkela_wire_6193),
        .c(new_Jinkela_wire_6194)
    );

    bfr new_Jinkela_buffer_7854 (
        .din(new_Jinkela_wire_9903),
        .dout(new_Jinkela_wire_9904)
    );

    bfr new_Jinkela_buffer_7829 (
        .din(new_Jinkela_wire_9871),
        .dout(new_Jinkela_wire_9872)
    );

    bfr new_Jinkela_buffer_5167 (
        .din(new_Jinkela_wire_6176),
        .dout(new_Jinkela_wire_6177)
    );

    bfr new_Jinkela_buffer_5178 (
        .din(new_Jinkela_wire_6199),
        .dout(new_Jinkela_wire_6200)
    );

    bfr new_Jinkela_buffer_7830 (
        .din(new_Jinkela_wire_9872),
        .dout(new_Jinkela_wire_9873)
    );

    bfr new_Jinkela_buffer_5168 (
        .din(new_Jinkela_wire_6177),
        .dout(new_Jinkela_wire_6178)
    );

    bfr new_Jinkela_buffer_7870 (
        .din(new_Jinkela_wire_9926),
        .dout(new_Jinkela_wire_9927)
    );

    bfr new_Jinkela_buffer_5217 (
        .din(new_Jinkela_wire_6238),
        .dout(new_Jinkela_wire_6239)
    );

    bfr new_Jinkela_buffer_7855 (
        .din(new_Jinkela_wire_9904),
        .dout(new_Jinkela_wire_9905)
    );

    bfr new_Jinkela_buffer_7831 (
        .din(new_Jinkela_wire_9873),
        .dout(new_Jinkela_wire_9874)
    );

    bfr new_Jinkela_buffer_5169 (
        .din(new_Jinkela_wire_6178),
        .dout(new_Jinkela_wire_6179)
    );

    spl2 new_Jinkela_splitter_823 (
        .a(new_Jinkela_wire_9918),
        .b(new_Jinkela_wire_9919),
        .c(new_Jinkela_wire_9920)
    );

    spl4L new_Jinkela_splitter_395 (
        .a(n_0750_),
        .d(new_Jinkela_wire_6250),
        .b(new_Jinkela_wire_6251),
        .e(new_Jinkela_wire_6252),
        .c(new_Jinkela_wire_6253)
    );

    bfr new_Jinkela_buffer_7832 (
        .din(new_Jinkela_wire_9874),
        .dout(new_Jinkela_wire_9875)
    );

    bfr new_Jinkela_buffer_5170 (
        .din(new_Jinkela_wire_6179),
        .dout(new_Jinkela_wire_6180)
    );

    bfr new_Jinkela_buffer_5218 (
        .din(new_Jinkela_wire_6239),
        .dout(new_Jinkela_wire_6240)
    );

    bfr new_Jinkela_buffer_7856 (
        .din(new_Jinkela_wire_9905),
        .dout(new_Jinkela_wire_9906)
    );

    bfr new_Jinkela_buffer_5179 (
        .din(new_Jinkela_wire_6200),
        .dout(new_Jinkela_wire_6201)
    );

    bfr new_Jinkela_buffer_7833 (
        .din(new_Jinkela_wire_9875),
        .dout(new_Jinkela_wire_9876)
    );

    bfr new_Jinkela_buffer_5171 (
        .din(new_Jinkela_wire_6180),
        .dout(new_Jinkela_wire_6181)
    );

    bfr new_Jinkela_buffer_7834 (
        .din(new_Jinkela_wire_9876),
        .dout(new_Jinkela_wire_9877)
    );

    bfr new_Jinkela_buffer_5172 (
        .din(new_Jinkela_wire_6181),
        .dout(new_Jinkela_wire_6182)
    );

    bfr new_Jinkela_buffer_7871 (
        .din(new_Jinkela_wire_9932),
        .dout(new_Jinkela_wire_9933)
    );

    bfr new_Jinkela_buffer_7857 (
        .din(new_Jinkela_wire_9906),
        .dout(new_Jinkela_wire_9907)
    );

    bfr new_Jinkela_buffer_5180 (
        .din(new_Jinkela_wire_6201),
        .dout(new_Jinkela_wire_6202)
    );

    bfr new_Jinkela_buffer_7835 (
        .din(new_Jinkela_wire_9877),
        .dout(new_Jinkela_wire_9878)
    );

    bfr new_Jinkela_buffer_5173 (
        .din(new_Jinkela_wire_6182),
        .dout(new_Jinkela_wire_6183)
    );

    bfr new_Jinkela_buffer_7894 (
        .din(n_1279_),
        .dout(new_Jinkela_wire_9956)
    );

    bfr new_Jinkela_buffer_7836 (
        .din(new_Jinkela_wire_9878),
        .dout(new_Jinkela_wire_9879)
    );

    bfr new_Jinkela_buffer_5174 (
        .din(new_Jinkela_wire_6183),
        .dout(new_Jinkela_wire_6184)
    );

    bfr new_Jinkela_buffer_5219 (
        .din(new_Jinkela_wire_6240),
        .dout(new_Jinkela_wire_6241)
    );

    bfr new_Jinkela_buffer_7858 (
        .din(new_Jinkela_wire_9907),
        .dout(new_Jinkela_wire_9908)
    );

    bfr new_Jinkela_buffer_5181 (
        .din(new_Jinkela_wire_6202),
        .dout(new_Jinkela_wire_6203)
    );

    bfr new_Jinkela_buffer_7837 (
        .din(new_Jinkela_wire_9879),
        .dout(new_Jinkela_wire_9880)
    );

    bfr new_Jinkela_buffer_5224 (
        .din(n_0340_),
        .dout(new_Jinkela_wire_6248)
    );

    bfr new_Jinkela_buffer_5182 (
        .din(new_Jinkela_wire_6203),
        .dout(new_Jinkela_wire_6204)
    );

    bfr new_Jinkela_buffer_7838 (
        .din(new_Jinkela_wire_9880),
        .dout(new_Jinkela_wire_9881)
    );

    bfr new_Jinkela_buffer_5226 (
        .din(n_1331_),
        .dout(new_Jinkela_wire_6254)
    );

    spl2 new_Jinkela_splitter_827 (
        .a(n_0741_),
        .b(new_Jinkela_wire_9957),
        .c(new_Jinkela_wire_9958)
    );

    bfr new_Jinkela_buffer_5220 (
        .din(new_Jinkela_wire_6241),
        .dout(new_Jinkela_wire_6242)
    );

    bfr new_Jinkela_buffer_7859 (
        .din(new_Jinkela_wire_9908),
        .dout(new_Jinkela_wire_9909)
    );

    bfr new_Jinkela_buffer_5183 (
        .din(new_Jinkela_wire_6204),
        .dout(new_Jinkela_wire_6205)
    );

    bfr new_Jinkela_buffer_7839 (
        .din(new_Jinkela_wire_9881),
        .dout(new_Jinkela_wire_9882)
    );

    bfr new_Jinkela_buffer_5225 (
        .din(new_Jinkela_wire_6248),
        .dout(new_Jinkela_wire_6249)
    );

    spl2 new_Jinkela_splitter_828 (
        .a(n_0467_),
        .b(new_Jinkela_wire_9959),
        .c(new_Jinkela_wire_9960)
    );

    bfr new_Jinkela_buffer_5184 (
        .din(new_Jinkela_wire_6205),
        .dout(new_Jinkela_wire_6206)
    );

    bfr new_Jinkela_buffer_7840 (
        .din(new_Jinkela_wire_9882),
        .dout(new_Jinkela_wire_9883)
    );

    bfr new_Jinkela_buffer_5221 (
        .din(new_Jinkela_wire_6242),
        .dout(new_Jinkela_wire_6243)
    );

    bfr new_Jinkela_buffer_7860 (
        .din(new_Jinkela_wire_9909),
        .dout(new_Jinkela_wire_9910)
    );

    bfr new_Jinkela_buffer_5185 (
        .din(new_Jinkela_wire_6206),
        .dout(new_Jinkela_wire_6207)
    );

    spl2 new_Jinkela_splitter_820 (
        .a(new_Jinkela_wire_9883),
        .b(new_Jinkela_wire_9884),
        .c(new_Jinkela_wire_9885)
    );

    bfr new_Jinkela_buffer_7872 (
        .din(new_Jinkela_wire_9933),
        .dout(new_Jinkela_wire_9934)
    );

    bfr new_Jinkela_buffer_7861 (
        .din(new_Jinkela_wire_9910),
        .dout(new_Jinkela_wire_9911)
    );

    bfr new_Jinkela_buffer_5186 (
        .din(new_Jinkela_wire_6207),
        .dout(new_Jinkela_wire_6208)
    );

    spl3L new_Jinkela_splitter_397 (
        .a(n_0788_),
        .d(new_Jinkela_wire_6261),
        .b(new_Jinkela_wire_6262),
        .c(new_Jinkela_wire_6263)
    );

    bfr new_Jinkela_buffer_5222 (
        .din(new_Jinkela_wire_6243),
        .dout(new_Jinkela_wire_6244)
    );

    bfr new_Jinkela_buffer_5187 (
        .din(new_Jinkela_wire_6208),
        .dout(new_Jinkela_wire_6209)
    );

    bfr new_Jinkela_buffer_7862 (
        .din(new_Jinkela_wire_9911),
        .dout(new_Jinkela_wire_9912)
    );

    bfr new_Jinkela_buffer_5188 (
        .din(new_Jinkela_wire_6209),
        .dout(new_Jinkela_wire_6210)
    );

    bfr new_Jinkela_buffer_7873 (
        .din(new_Jinkela_wire_9934),
        .dout(new_Jinkela_wire_9935)
    );

    bfr new_Jinkela_buffer_7863 (
        .din(new_Jinkela_wire_9912),
        .dout(new_Jinkela_wire_9913)
    );

    spl2 new_Jinkela_splitter_398 (
        .a(n_1238_),
        .b(new_Jinkela_wire_6264),
        .c(new_Jinkela_wire_6265)
    );

    bfr new_Jinkela_buffer_5189 (
        .din(new_Jinkela_wire_6210),
        .dout(new_Jinkela_wire_6211)
    );

    spl2 new_Jinkela_splitter_829 (
        .a(n_0060_),
        .b(new_Jinkela_wire_9961),
        .c(new_Jinkela_wire_9962)
    );

    bfr new_Jinkela_buffer_5231 (
        .din(new_net_2560),
        .dout(new_Jinkela_wire_6266)
    );

    bfr new_Jinkela_buffer_7874 (
        .din(new_Jinkela_wire_9935),
        .dout(new_Jinkela_wire_9936)
    );

    bfr new_Jinkela_buffer_5227 (
        .din(new_Jinkela_wire_6254),
        .dout(new_Jinkela_wire_6255)
    );

    bfr new_Jinkela_buffer_5190 (
        .din(new_Jinkela_wire_6211),
        .dout(new_Jinkela_wire_6212)
    );

    bfr new_Jinkela_buffer_7915 (
        .din(n_1259_),
        .dout(new_Jinkela_wire_9983)
    );

    bfr new_Jinkela_buffer_7895 (
        .din(new_Jinkela_wire_9962),
        .dout(new_Jinkela_wire_9963)
    );

    bfr new_Jinkela_buffer_7875 (
        .din(new_Jinkela_wire_9936),
        .dout(new_Jinkela_wire_9937)
    );

    bfr new_Jinkela_buffer_5228 (
        .din(new_Jinkela_wire_6255),
        .dout(new_Jinkela_wire_6256)
    );

    bfr new_Jinkela_buffer_5191 (
        .din(new_Jinkela_wire_6212),
        .dout(new_Jinkela_wire_6213)
    );

    spl2 new_Jinkela_splitter_830 (
        .a(new_net_4),
        .b(new_Jinkela_wire_9984),
        .c(new_Jinkela_wire_9985)
    );

    spl3L new_Jinkela_splitter_831 (
        .a(n_0140_),
        .d(new_Jinkela_wire_10030),
        .b(new_Jinkela_wire_10031),
        .c(new_Jinkela_wire_10032)
    );

    bfr new_Jinkela_buffer_7876 (
        .din(new_Jinkela_wire_9937),
        .dout(new_Jinkela_wire_9938)
    );

    bfr new_Jinkela_buffer_1865 (
        .din(new_Jinkela_wire_2219),
        .dout(new_Jinkela_wire_2220)
    );

    bfr new_Jinkela_buffer_1866 (
        .din(new_Jinkela_wire_2220),
        .dout(new_Jinkela_wire_2221)
    );

    bfr new_Jinkela_buffer_2079 (
        .din(new_Jinkela_wire_2448),
        .dout(new_Jinkela_wire_2449)
    );

    bfr new_Jinkela_buffer_1904 (
        .din(new_Jinkela_wire_2264),
        .dout(new_Jinkela_wire_2265)
    );

    bfr new_Jinkela_buffer_1867 (
        .din(new_Jinkela_wire_2221),
        .dout(new_Jinkela_wire_2222)
    );

    bfr new_Jinkela_buffer_1868 (
        .din(new_Jinkela_wire_2222),
        .dout(new_Jinkela_wire_2223)
    );

    bfr new_Jinkela_buffer_1956 (
        .din(new_Jinkela_wire_2320),
        .dout(new_Jinkela_wire_2321)
    );

    bfr new_Jinkela_buffer_1905 (
        .din(new_Jinkela_wire_2265),
        .dout(new_Jinkela_wire_2266)
    );

    bfr new_Jinkela_buffer_1869 (
        .din(new_Jinkela_wire_2223),
        .dout(new_Jinkela_wire_2224)
    );

    bfr new_Jinkela_buffer_1870 (
        .din(new_Jinkela_wire_2224),
        .dout(new_Jinkela_wire_2225)
    );

    bfr new_Jinkela_buffer_2082 (
        .din(new_Jinkela_wire_2451),
        .dout(new_Jinkela_wire_2452)
    );

    bfr new_Jinkela_buffer_1906 (
        .din(new_Jinkela_wire_2266),
        .dout(new_Jinkela_wire_2267)
    );

    bfr new_Jinkela_buffer_1871 (
        .din(new_Jinkela_wire_2225),
        .dout(new_Jinkela_wire_2226)
    );

    bfr new_Jinkela_buffer_1872 (
        .din(new_Jinkela_wire_2226),
        .dout(new_Jinkela_wire_2227)
    );

    bfr new_Jinkela_buffer_1957 (
        .din(new_Jinkela_wire_2321),
        .dout(new_Jinkela_wire_2322)
    );

    bfr new_Jinkela_buffer_1907 (
        .din(new_Jinkela_wire_2267),
        .dout(new_Jinkela_wire_2268)
    );

    bfr new_Jinkela_buffer_1873 (
        .din(new_Jinkela_wire_2227),
        .dout(new_Jinkela_wire_2228)
    );

    bfr new_Jinkela_buffer_1874 (
        .din(new_Jinkela_wire_2228),
        .dout(new_Jinkela_wire_2229)
    );

    bfr new_Jinkela_buffer_2017 (
        .din(new_Jinkela_wire_2383),
        .dout(new_Jinkela_wire_2384)
    );

    bfr new_Jinkela_buffer_1908 (
        .din(new_Jinkela_wire_2268),
        .dout(new_Jinkela_wire_2269)
    );

    bfr new_Jinkela_buffer_1875 (
        .din(new_Jinkela_wire_2229),
        .dout(new_Jinkela_wire_2230)
    );

    bfr new_Jinkela_buffer_1876 (
        .din(new_Jinkela_wire_2230),
        .dout(new_Jinkela_wire_2231)
    );

    bfr new_Jinkela_buffer_1958 (
        .din(new_Jinkela_wire_2322),
        .dout(new_Jinkela_wire_2323)
    );

    bfr new_Jinkela_buffer_1909 (
        .din(new_Jinkela_wire_2269),
        .dout(new_Jinkela_wire_2270)
    );

    bfr new_Jinkela_buffer_1877 (
        .din(new_Jinkela_wire_2231),
        .dout(new_Jinkela_wire_2232)
    );

    bfr new_Jinkela_buffer_2080 (
        .din(new_Jinkela_wire_2449),
        .dout(new_Jinkela_wire_2450)
    );

    bfr new_Jinkela_buffer_1910 (
        .din(new_Jinkela_wire_2270),
        .dout(new_Jinkela_wire_2271)
    );

    bfr new_Jinkela_buffer_1959 (
        .din(new_Jinkela_wire_2323),
        .dout(new_Jinkela_wire_2324)
    );

    bfr new_Jinkela_buffer_1911 (
        .din(new_Jinkela_wire_2271),
        .dout(new_Jinkela_wire_2272)
    );

    bfr new_Jinkela_buffer_2018 (
        .din(new_Jinkela_wire_2384),
        .dout(new_Jinkela_wire_2385)
    );

    bfr new_Jinkela_buffer_1912 (
        .din(new_Jinkela_wire_2272),
        .dout(new_Jinkela_wire_2273)
    );

    bfr new_Jinkela_buffer_1960 (
        .din(new_Jinkela_wire_2324),
        .dout(new_Jinkela_wire_2325)
    );

    bfr new_Jinkela_buffer_1913 (
        .din(new_Jinkela_wire_2273),
        .dout(new_Jinkela_wire_2274)
    );

    bfr new_Jinkela_buffer_2089 (
        .din(N221),
        .dout(new_Jinkela_wire_2459)
    );

    bfr new_Jinkela_buffer_1914 (
        .din(new_Jinkela_wire_2274),
        .dout(new_Jinkela_wire_2275)
    );

    bfr new_Jinkela_buffer_1961 (
        .din(new_Jinkela_wire_2325),
        .dout(new_Jinkela_wire_2326)
    );

    bfr new_Jinkela_buffer_1915 (
        .din(new_Jinkela_wire_2275),
        .dout(new_Jinkela_wire_2276)
    );

    spl3L new_Jinkela_splitter_120 (
        .a(new_Jinkela_wire_2385),
        .d(new_Jinkela_wire_2386),
        .b(new_Jinkela_wire_2387),
        .c(new_Jinkela_wire_2388)
    );

    bfr new_Jinkela_buffer_1916 (
        .din(new_Jinkela_wire_2276),
        .dout(new_Jinkela_wire_2277)
    );

    bfr new_Jinkela_buffer_1962 (
        .din(new_Jinkela_wire_2326),
        .dout(new_Jinkela_wire_2327)
    );

    bfr new_Jinkela_buffer_1917 (
        .din(new_Jinkela_wire_2277),
        .dout(new_Jinkela_wire_2278)
    );

    and_bb n_2748_ (
        .a(new_Jinkela_wire_8175),
        .b(new_Jinkela_wire_3919),
        .c(n_0604_)
    );

    and_ii n_2031_ (
        .a(new_Jinkela_wire_9343),
        .b(new_Jinkela_wire_7463),
        .c(n_1296_)
    );

    or_bb n_2749_ (
        .a(n_0604_),
        .b(n_0603_),
        .c(n_0605_)
    );

    bfr new_Jinkela_buffer_2787 (
        .din(N340),
        .dout(new_Jinkela_wire_3202)
    );

    inv n_2032_ (
        .din(new_Jinkela_wire_1018),
        .dout(n_1297_)
    );

    bfr new_Jinkela_buffer_355 (
        .din(new_Jinkela_wire_386),
        .dout(new_Jinkela_wire_387)
    );

    and_bi n_2750_ (
        .a(new_Jinkela_wire_4920),
        .b(new_Jinkela_wire_8402),
        .c(n_0606_)
    );

    and_bi n_2033_ (
        .a(new_Jinkela_wire_8009),
        .b(new_Jinkela_wire_5295),
        .c(n_1298_)
    );

    bfr new_Jinkela_buffer_545 (
        .din(N214),
        .dout(new_Jinkela_wire_587)
    );

    or_bb n_2751_ (
        .a(n_0606_),
        .b(new_Jinkela_wire_5224),
        .c(n_0607_)
    );

    bfr new_Jinkela_buffer_2659 (
        .din(new_Jinkela_wire_3068),
        .dout(new_Jinkela_wire_3069)
    );

    bfr new_Jinkela_buffer_412 (
        .din(new_Jinkela_wire_448),
        .dout(new_Jinkela_wire_449)
    );

    and_bi n_2034_ (
        .a(new_Jinkela_wire_5293),
        .b(new_Jinkela_wire_8008),
        .c(n_1299_)
    );

    bfr new_Jinkela_buffer_356 (
        .din(new_Jinkela_wire_387),
        .dout(new_Jinkela_wire_388)
    );

    and_bi n_2752_ (
        .a(new_Jinkela_wire_6311),
        .b(n_0607_),
        .c(n_0608_)
    );

    inv n_2035_ (
        .din(new_Jinkela_wire_800),
        .dout(n_1300_)
    );

    and_bb n_2753_ (
        .a(new_Jinkela_wire_9768),
        .b(new_Jinkela_wire_4781),
        .c(n_0609_)
    );

    spl3L new_Jinkela_splitter_139 (
        .a(new_Jinkela_wire_3128),
        .d(new_Jinkela_wire_3129),
        .b(new_Jinkela_wire_3130),
        .c(new_Jinkela_wire_3131)
    );

    bfr new_Jinkela_buffer_477 (
        .din(new_Jinkela_wire_513),
        .dout(new_Jinkela_wire_514)
    );

    and_bi n_2036_ (
        .a(new_Jinkela_wire_5229),
        .b(new_Jinkela_wire_7233),
        .c(n_1301_)
    );

    bfr new_Jinkela_buffer_357 (
        .din(new_Jinkela_wire_388),
        .dout(new_Jinkela_wire_389)
    );

    or_ii n_2754_ (
        .a(new_Jinkela_wire_5069),
        .b(new_Jinkela_wire_5217),
        .c(n_0610_)
    );

    and_bi n_2037_ (
        .a(new_Jinkela_wire_7232),
        .b(new_Jinkela_wire_5228),
        .c(n_1302_)
    );

    bfr new_Jinkela_buffer_540 (
        .din(new_Jinkela_wire_581),
        .dout(new_Jinkela_wire_582)
    );

    and_bi n_2755_ (
        .a(new_Jinkela_wire_8401),
        .b(new_Jinkela_wire_5873),
        .c(n_0611_)
    );

    inv n_2038_ (
        .din(new_Jinkela_wire_6535),
        .dout(n_1303_)
    );

    bfr new_Jinkela_buffer_2616 (
        .din(new_Jinkela_wire_3021),
        .dout(new_Jinkela_wire_3022)
    );

    bfr new_Jinkela_buffer_358 (
        .din(new_Jinkela_wire_389),
        .dout(new_Jinkela_wire_390)
    );

    or_bb n_2756_ (
        .a(n_0611_),
        .b(new_Jinkela_wire_5572),
        .c(n_0612_)
    );

    inv n_2039_ (
        .din(new_Jinkela_wire_1541),
        .dout(n_1304_)
    );

    or_bb n_2757_ (
        .a(new_Jinkela_wire_6790),
        .b(n_0608_),
        .c(n_0613_)
    );

    bfr new_Jinkela_buffer_2781 (
        .din(new_Jinkela_wire_3195),
        .dout(new_Jinkela_wire_3196)
    );

    and_bi n_2040_ (
        .a(new_Jinkela_wire_7684),
        .b(new_Jinkela_wire_9842),
        .c(n_1305_)
    );

    bfr new_Jinkela_buffer_2617 (
        .din(new_Jinkela_wire_3022),
        .dout(new_Jinkela_wire_3023)
    );

    bfr new_Jinkela_buffer_359 (
        .din(new_Jinkela_wire_390),
        .dout(new_Jinkela_wire_391)
    );

    and_bb n_2758_ (
        .a(new_Jinkela_wire_5560),
        .b(new_Jinkela_wire_9738),
        .c(n_0614_)
    );

    and_bi n_2041_ (
        .a(new_Jinkela_wire_9841),
        .b(new_Jinkela_wire_7683),
        .c(n_1306_)
    );

    bfr new_Jinkela_buffer_476 (
        .din(new_Jinkela_wire_512),
        .dout(new_Jinkela_wire_513)
    );

    or_bb n_2759_ (
        .a(new_Jinkela_wire_9135),
        .b(new_Jinkela_wire_7322),
        .c(n_0615_)
    );

    bfr new_Jinkela_buffer_2661 (
        .din(new_Jinkela_wire_3070),
        .dout(new_Jinkela_wire_3071)
    );

    bfr new_Jinkela_buffer_414 (
        .din(new_Jinkela_wire_450),
        .dout(new_Jinkela_wire_451)
    );

    inv n_2042_ (
        .din(new_Jinkela_wire_2306),
        .dout(n_1307_)
    );

    and_bi n_2760_ (
        .a(new_Jinkela_wire_8170),
        .b(new_Jinkela_wire_4661),
        .c(n_0616_)
    );

    and_bi n_2043_ (
        .a(new_Jinkela_wire_8656),
        .b(new_Jinkela_wire_9469),
        .c(n_1308_)
    );

    and_bb n_2761_ (
        .a(new_Jinkela_wire_8936),
        .b(new_Jinkela_wire_6104),
        .c(n_0617_)
    );

    bfr new_Jinkela_buffer_2717 (
        .din(new_Jinkela_wire_3131),
        .dout(new_Jinkela_wire_3132)
    );

    spl2 new_Jinkela_splitter_16 (
        .a(new_Jinkela_wire_514),
        .b(new_Jinkela_wire_515),
        .c(new_Jinkela_wire_516)
    );

    and_ii n_2044_ (
        .a(new_Jinkela_wire_4309),
        .b(new_Jinkela_wire_3781),
        .c(n_1309_)
    );

    and_bi n_2762_ (
        .a(new_Jinkela_wire_8277),
        .b(new_Jinkela_wire_5280),
        .c(n_0618_)
    );

    and_ii n_2045_ (
        .a(new_Jinkela_wire_8708),
        .b(new_Jinkela_wire_8873),
        .c(n_1310_)
    );

    and_bi n_2763_ (
        .a(new_Jinkela_wire_8748),
        .b(new_Jinkela_wire_7757),
        .c(n_0619_)
    );

    bfr new_Jinkela_buffer_2662 (
        .din(new_Jinkela_wire_3071),
        .dout(new_Jinkela_wire_3072)
    );

    bfr new_Jinkela_buffer_415 (
        .din(new_Jinkela_wire_451),
        .dout(new_Jinkela_wire_452)
    );

    and_bi n_2046_ (
        .a(new_Jinkela_wire_3875),
        .b(new_Jinkela_wire_10528),
        .c(n_1311_)
    );

    and_bi n_2764_ (
        .a(new_Jinkela_wire_7758),
        .b(new_Jinkela_wire_8747),
        .c(n_0620_)
    );

    or_bb n_2047_ (
        .a(n_1311_),
        .b(new_Jinkela_wire_6813),
        .c(n_1312_)
    );

    and_ii n_2765_ (
        .a(n_0620_),
        .b(n_0619_),
        .c(n_0621_)
    );

    inv n_2048_ (
        .din(new_Jinkela_wire_6806),
        .dout(n_1313_)
    );

    bfr new_Jinkela_buffer_2621 (
        .din(new_Jinkela_wire_3026),
        .dout(new_Jinkela_wire_3027)
    );

    bfr new_Jinkela_buffer_363 (
        .din(new_Jinkela_wire_394),
        .dout(new_Jinkela_wire_395)
    );

    and_bi n_2766_ (
        .a(new_Jinkela_wire_4958),
        .b(new_Jinkela_wire_6330),
        .c(n_0622_)
    );

    and_ii n_2049_ (
        .a(new_Jinkela_wire_3782),
        .b(new_Jinkela_wire_8870),
        .c(n_1314_)
    );

    and_bi n_2767_ (
        .a(new_Jinkela_wire_6329),
        .b(new_Jinkela_wire_4957),
        .c(n_0623_)
    );

    and_bi n_2050_ (
        .a(new_Jinkela_wire_9472),
        .b(new_Jinkela_wire_8655),
        .c(n_1315_)
    );

    bfr new_Jinkela_buffer_2622 (
        .din(new_Jinkela_wire_3027),
        .dout(new_Jinkela_wire_3028)
    );

    bfr new_Jinkela_buffer_364 (
        .din(new_Jinkela_wire_395),
        .dout(new_Jinkela_wire_396)
    );

    or_bb n_2768_ (
        .a(n_0623_),
        .b(n_0622_),
        .c(n_0624_)
    );

    or_bb n_2051_ (
        .a(new_Jinkela_wire_9773),
        .b(new_Jinkela_wire_4308),
        .c(n_1316_)
    );

    and_ii n_2769_ (
        .a(new_Jinkela_wire_6131),
        .b(new_Jinkela_wire_7920),
        .c(n_0625_)
    );

    and_bi n_2052_ (
        .a(new_Jinkela_wire_3793),
        .b(new_Jinkela_wire_10390),
        .c(n_1317_)
    );

    bfr new_Jinkela_buffer_2623 (
        .din(new_Jinkela_wire_3028),
        .dout(new_Jinkela_wire_3029)
    );

    bfr new_Jinkela_buffer_365 (
        .din(new_Jinkela_wire_396),
        .dout(new_Jinkela_wire_397)
    );

    and_bb n_2770_ (
        .a(new_Jinkela_wire_6130),
        .b(new_Jinkela_wire_7919),
        .c(n_0626_)
    );

    or_ii n_2053_ (
        .a(new_Jinkela_wire_5731),
        .b(new_Jinkela_wire_6533),
        .c(n_1318_)
    );

    or_bb n_2771_ (
        .a(n_0626_),
        .b(new_Jinkela_wire_2581),
        .c(n_0627_)
    );

    bfr new_Jinkela_buffer_2664 (
        .din(new_Jinkela_wire_3073),
        .dout(new_Jinkela_wire_3074)
    );

    bfr new_Jinkela_buffer_417 (
        .din(new_Jinkela_wire_453),
        .dout(new_Jinkela_wire_454)
    );

    or_ii n_2054_ (
        .a(new_Jinkela_wire_7729),
        .b(new_Jinkela_wire_5343),
        .c(n_1319_)
    );

    bfr new_Jinkela_buffer_2624 (
        .din(new_Jinkela_wire_3029),
        .dout(new_Jinkela_wire_3030)
    );

    bfr new_Jinkela_buffer_366 (
        .din(new_Jinkela_wire_397),
        .dout(new_Jinkela_wire_398)
    );

    or_bb n_2772_ (
        .a(n_0627_),
        .b(new_Jinkela_wire_4171),
        .c(n_0628_)
    );

    or_bb n_2055_ (
        .a(new_Jinkela_wire_9764),
        .b(new_Jinkela_wire_3210),
        .c(n_1320_)
    );

    and_ii n_2773_ (
        .a(new_Jinkela_wire_5563),
        .b(new_Jinkela_wire_7992),
        .c(n_0629_)
    );

    bfr new_Jinkela_buffer_2782 (
        .din(new_Jinkela_wire_3196),
        .dout(new_Jinkela_wire_3197)
    );

    bfr new_Jinkela_buffer_541 (
        .din(new_Jinkela_wire_582),
        .dout(new_Jinkela_wire_583)
    );

    inv n_2056_ (
        .din(new_Jinkela_wire_105),
        .dout(n_1321_)
    );

    bfr new_Jinkela_buffer_2625 (
        .din(new_Jinkela_wire_3030),
        .dout(new_Jinkela_wire_3031)
    );

    and_ii n_2774_ (
        .a(new_Jinkela_wire_4509),
        .b(new_Jinkela_wire_5453),
        .c(n_0630_)
    );

    and_bi n_2057_ (
        .a(new_Jinkela_wire_10365),
        .b(new_Jinkela_wire_7223),
        .c(n_1322_)
    );

    or_bi n_2775_ (
        .a(new_Jinkela_wire_7752),
        .b(new_Jinkela_wire_8171),
        .c(n_0631_)
    );

    bfr new_Jinkela_buffer_2665 (
        .din(new_Jinkela_wire_3074),
        .dout(new_Jinkela_wire_3075)
    );

    bfr new_Jinkela_buffer_418 (
        .din(new_Jinkela_wire_454),
        .dout(new_Jinkela_wire_455)
    );

    and_bi n_2058_ (
        .a(new_Jinkela_wire_9927),
        .b(new_Jinkela_wire_4082),
        .c(n_1323_)
    );

    bfr new_Jinkela_buffer_2626 (
        .din(new_Jinkela_wire_3031),
        .dout(new_Jinkela_wire_3032)
    );

    bfr new_Jinkela_buffer_368 (
        .din(new_Jinkela_wire_399),
        .dout(new_Jinkela_wire_400)
    );

    and_bi n_2776_ (
        .a(new_Jinkela_wire_5457),
        .b(n_0631_),
        .c(n_0632_)
    );

    and_bb n_2059_ (
        .a(new_Jinkela_wire_9763),
        .b(new_Jinkela_wire_3211),
        .c(n_1324_)
    );

    and_ii n_2777_ (
        .a(n_0632_),
        .b(new_Jinkela_wire_7085),
        .c(n_0633_)
    );

    bfr new_Jinkela_buffer_2719 (
        .din(new_Jinkela_wire_3133),
        .dout(new_Jinkela_wire_3134)
    );

    bfr new_Jinkela_buffer_544 (
        .din(new_Jinkela_wire_585),
        .dout(new_Jinkela_wire_586)
    );

    and_bi n_2060_ (
        .a(new_Jinkela_wire_7222),
        .b(new_Jinkela_wire_10363),
        .c(n_1325_)
    );

    bfr new_Jinkela_buffer_2627 (
        .din(new_Jinkela_wire_3032),
        .dout(new_Jinkela_wire_3033)
    );

    bfr new_Jinkela_buffer_369 (
        .din(new_Jinkela_wire_400),
        .dout(new_Jinkela_wire_401)
    );

    or_bi n_2778_ (
        .a(new_Jinkela_wire_10103),
        .b(new_Jinkela_wire_9647),
        .c(n_0634_)
    );

    and_ii n_2061_ (
        .a(new_Jinkela_wire_8759),
        .b(new_Jinkela_wire_9395),
        .c(n_1326_)
    );

    and_bi n_2779_ (
        .a(new_Jinkela_wire_10102),
        .b(new_Jinkela_wire_9646),
        .c(n_0635_)
    );

    bfr new_Jinkela_buffer_2666 (
        .din(new_Jinkela_wire_3075),
        .dout(new_Jinkela_wire_3076)
    );

    bfr new_Jinkela_buffer_419 (
        .din(new_Jinkela_wire_455),
        .dout(new_Jinkela_wire_456)
    );

    and_bb n_2062_ (
        .a(new_Jinkela_wire_7226),
        .b(new_Jinkela_wire_10147),
        .c(n_1327_)
    );

    bfr new_Jinkela_buffer_2628 (
        .din(new_Jinkela_wire_3033),
        .dout(new_Jinkela_wire_3034)
    );

    bfr new_Jinkela_buffer_370 (
        .din(new_Jinkela_wire_401),
        .dout(new_Jinkela_wire_402)
    );

    and_bi n_2780_ (
        .a(n_0634_),
        .b(n_0635_),
        .c(n_0636_)
    );

    and_bi n_2063_ (
        .a(new_Jinkela_wire_2387),
        .b(new_Jinkela_wire_10140),
        .c(n_1328_)
    );

    and_bi n_2781_ (
        .a(new_Jinkela_wire_8182),
        .b(new_Jinkela_wire_4961),
        .c(n_0637_)
    );

    bfr new_Jinkela_buffer_479 (
        .din(new_Jinkela_wire_517),
        .dout(new_Jinkela_wire_518)
    );

    and_bi n_2064_ (
        .a(new_Jinkela_wire_10138),
        .b(new_Jinkela_wire_2386),
        .c(n_1329_)
    );

    bfr new_Jinkela_buffer_2629 (
        .din(new_Jinkela_wire_3034),
        .dout(new_Jinkela_wire_3035)
    );

    bfr new_Jinkela_buffer_371 (
        .din(new_Jinkela_wire_402),
        .dout(new_Jinkela_wire_403)
    );

    and_bi n_2782_ (
        .a(new_Jinkela_wire_4962),
        .b(new_Jinkela_wire_8181),
        .c(n_0638_)
    );

    and_ii n_2065_ (
        .a(new_Jinkela_wire_5577),
        .b(new_Jinkela_wire_6087),
        .c(n_1330_)
    );

    spl2 new_Jinkela_splitter_142 (
        .a(N322),
        .b(new_Jinkela_wire_3271),
        .c(new_Jinkela_wire_3272)
    );

    or_bb n_2783_ (
        .a(n_0638_),
        .b(n_0637_),
        .c(n_0639_)
    );

    bfr new_Jinkela_buffer_420 (
        .din(new_Jinkela_wire_456),
        .dout(new_Jinkela_wire_457)
    );

    inv n_2066_ (
        .din(new_Jinkela_wire_200),
        .dout(n_1331_)
    );

    bfr new_Jinkela_buffer_2630 (
        .din(new_Jinkela_wire_3035),
        .dout(new_Jinkela_wire_3036)
    );

    bfr new_Jinkela_buffer_372 (
        .din(new_Jinkela_wire_403),
        .dout(new_Jinkela_wire_404)
    );

    or_bi n_2784_ (
        .a(new_Jinkela_wire_4660),
        .b(new_Jinkela_wire_6322),
        .c(n_0640_)
    );

    and_bi n_2067_ (
        .a(new_Jinkela_wire_9921),
        .b(new_Jinkela_wire_6260),
        .c(n_1332_)
    );

    and_bi n_2785_ (
        .a(new_Jinkela_wire_4659),
        .b(new_Jinkela_wire_6321),
        .c(n_0641_)
    );

    bfr new_Jinkela_buffer_542 (
        .din(new_Jinkela_wire_583),
        .dout(new_Jinkela_wire_584)
    );

    and_bi n_2068_ (
        .a(new_Jinkela_wire_6259),
        .b(new_Jinkela_wire_9922),
        .c(n_1333_)
    );

    bfr new_Jinkela_buffer_2631 (
        .din(new_Jinkela_wire_3036),
        .dout(new_Jinkela_wire_3037)
    );

    bfr new_Jinkela_buffer_373 (
        .din(new_Jinkela_wire_404),
        .dout(new_Jinkela_wire_405)
    );

    or_bb n_2786_ (
        .a(n_0641_),
        .b(new_Jinkela_wire_5222),
        .c(n_0642_)
    );

    and_ii n_2069_ (
        .a(new_Jinkela_wire_5918),
        .b(new_Jinkela_wire_7730),
        .c(n_1334_)
    );

    and_bi n_2787_ (
        .a(new_Jinkela_wire_8924),
        .b(n_0642_),
        .c(n_0643_)
    );

    bfr new_Jinkela_buffer_2668 (
        .din(new_Jinkela_wire_3077),
        .dout(new_Jinkela_wire_3078)
    );

    bfr new_Jinkela_buffer_421 (
        .din(new_Jinkela_wire_457),
        .dout(new_Jinkela_wire_458)
    );

    or_ii n_2070_ (
        .a(new_Jinkela_wire_5979),
        .b(new_Jinkela_wire_8625),
        .c(n_1335_)
    );

    bfr new_Jinkela_buffer_2632 (
        .din(new_Jinkela_wire_3037),
        .dout(new_Jinkela_wire_3038)
    );

    bfr new_Jinkela_buffer_374 (
        .din(new_Jinkela_wire_405),
        .dout(new_Jinkela_wire_406)
    );

    and_bi n_2788_ (
        .a(new_Jinkela_wire_9391),
        .b(n_0643_),
        .c(n_0644_)
    );

    or_bi n_2071_ (
        .a(new_Jinkela_wire_4437),
        .b(new_Jinkela_wire_7839),
        .c(n_1336_)
    );

    or_bi n_2789_ (
        .a(new_Jinkela_wire_8813),
        .b(new_Jinkela_wire_9585),
        .c(n_0645_)
    );

    bfr new_Jinkela_buffer_2785 (
        .din(new_Jinkela_wire_3199),
        .dout(new_Jinkela_wire_3200)
    );

    bfr new_Jinkela_buffer_480 (
        .din(new_Jinkela_wire_518),
        .dout(new_Jinkela_wire_519)
    );

    and_ii n_2072_ (
        .a(new_Jinkela_wire_4648),
        .b(new_Jinkela_wire_520),
        .c(n_1337_)
    );

    bfr new_Jinkela_buffer_2633 (
        .din(new_Jinkela_wire_3038),
        .dout(new_Jinkela_wire_3039)
    );

    bfr new_Jinkela_buffer_375 (
        .din(new_Jinkela_wire_406),
        .dout(new_Jinkela_wire_407)
    );

    bfr new_Jinkela_buffer_6834 (
        .din(n_1186_),
        .dout(new_Jinkela_wire_8450)
    );

    and_bi n_1419_ (
        .a(new_Jinkela_wire_7265),
        .b(new_Jinkela_wire_2744),
        .c(n_0691_)
    );

    bfr new_Jinkela_buffer_4322 (
        .din(new_Jinkela_wire_5122),
        .dout(new_Jinkela_wire_5123)
    );

    bfr new_Jinkela_buffer_6808 (
        .din(new_Jinkela_wire_8413),
        .dout(new_Jinkela_wire_8414)
    );

    spl2 new_Jinkela_splitter_311 (
        .a(n_0364_),
        .b(new_Jinkela_wire_5226),
        .c(new_Jinkela_wire_5227)
    );

    bfr new_Jinkela_buffer_6830 (
        .din(n_0409_),
        .dout(new_Jinkela_wire_8444)
    );

    bfr new_Jinkela_buffer_4323 (
        .din(new_Jinkela_wire_5123),
        .dout(new_Jinkela_wire_5124)
    );

    bfr new_Jinkela_buffer_6809 (
        .din(new_Jinkela_wire_8414),
        .dout(new_Jinkela_wire_8415)
    );

    spl4L new_Jinkela_splitter_312 (
        .a(n_0878_),
        .d(new_Jinkela_wire_5228),
        .b(new_Jinkela_wire_5229),
        .e(new_Jinkela_wire_5230),
        .c(new_Jinkela_wire_5231)
    );

    bfr new_Jinkela_buffer_6835 (
        .din(new_net_2509),
        .dout(new_Jinkela_wire_8451)
    );

    bfr new_Jinkela_buffer_4324 (
        .din(new_Jinkela_wire_5124),
        .dout(new_Jinkela_wire_5125)
    );

    bfr new_Jinkela_buffer_6810 (
        .din(new_Jinkela_wire_8415),
        .dout(new_Jinkela_wire_8416)
    );

    bfr new_Jinkela_buffer_4381 (
        .din(new_Jinkela_wire_5200),
        .dout(new_Jinkela_wire_5201)
    );

    bfr new_Jinkela_buffer_6831 (
        .din(new_Jinkela_wire_8444),
        .dout(new_Jinkela_wire_8445)
    );

    bfr new_Jinkela_buffer_4398 (
        .din(n_0276_),
        .dout(new_Jinkela_wire_5225)
    );

    bfr new_Jinkela_buffer_4325 (
        .din(new_Jinkela_wire_5125),
        .dout(new_Jinkela_wire_5126)
    );

    bfr new_Jinkela_buffer_6811 (
        .din(new_Jinkela_wire_8416),
        .dout(new_Jinkela_wire_8417)
    );

    spl2 new_Jinkela_splitter_645 (
        .a(n_1265_),
        .b(new_Jinkela_wire_8476),
        .c(new_Jinkela_wire_8477)
    );

    bfr new_Jinkela_buffer_4352 (
        .din(new_Jinkela_wire_5169),
        .dout(new_Jinkela_wire_5170)
    );

    bfr new_Jinkela_buffer_4326 (
        .din(new_Jinkela_wire_5126),
        .dout(new_Jinkela_wire_5127)
    );

    bfr new_Jinkela_buffer_6812 (
        .din(new_Jinkela_wire_8417),
        .dout(new_Jinkela_wire_8418)
    );

    bfr new_Jinkela_buffer_6832 (
        .din(new_Jinkela_wire_8445),
        .dout(new_Jinkela_wire_8446)
    );

    bfr new_Jinkela_buffer_4327 (
        .din(new_Jinkela_wire_5127),
        .dout(new_Jinkela_wire_5128)
    );

    bfr new_Jinkela_buffer_6813 (
        .din(new_Jinkela_wire_8418),
        .dout(new_Jinkela_wire_8419)
    );

    spl2 new_Jinkela_splitter_646 (
        .a(n_0120_),
        .b(new_Jinkela_wire_8478),
        .c(new_Jinkela_wire_8479)
    );

    bfr new_Jinkela_buffer_4353 (
        .din(new_Jinkela_wire_5170),
        .dout(new_Jinkela_wire_5171)
    );

    bfr new_Jinkela_buffer_6836 (
        .din(new_Jinkela_wire_8451),
        .dout(new_Jinkela_wire_8452)
    );

    bfr new_Jinkela_buffer_4328 (
        .din(new_Jinkela_wire_5128),
        .dout(new_Jinkela_wire_5129)
    );

    bfr new_Jinkela_buffer_6814 (
        .din(new_Jinkela_wire_8419),
        .dout(new_Jinkela_wire_8420)
    );

    bfr new_Jinkela_buffer_6833 (
        .din(new_Jinkela_wire_8446),
        .dout(new_Jinkela_wire_8447)
    );

    bfr new_Jinkela_buffer_4329 (
        .din(new_Jinkela_wire_5129),
        .dout(new_Jinkela_wire_5130)
    );

    bfr new_Jinkela_buffer_6815 (
        .din(new_Jinkela_wire_8420),
        .dout(new_Jinkela_wire_8421)
    );

    bfr new_Jinkela_buffer_4379 (
        .din(new_Jinkela_wire_5198),
        .dout(new_Jinkela_wire_5199)
    );

    bfr new_Jinkela_buffer_4354 (
        .din(new_Jinkela_wire_5171),
        .dout(new_Jinkela_wire_5172)
    );

    bfr new_Jinkela_buffer_4330 (
        .din(new_Jinkela_wire_5130),
        .dout(new_Jinkela_wire_5131)
    );

    bfr new_Jinkela_buffer_6816 (
        .din(new_Jinkela_wire_8421),
        .dout(new_Jinkela_wire_8422)
    );

    spl2 new_Jinkela_splitter_644 (
        .a(new_Jinkela_wire_8447),
        .b(new_Jinkela_wire_8448),
        .c(new_Jinkela_wire_8449)
    );

    bfr new_Jinkela_buffer_4331 (
        .din(new_Jinkela_wire_5131),
        .dout(new_Jinkela_wire_5132)
    );

    bfr new_Jinkela_buffer_6817 (
        .din(new_Jinkela_wire_8422),
        .dout(new_Jinkela_wire_8423)
    );

    bfr new_Jinkela_buffer_4355 (
        .din(new_Jinkela_wire_5172),
        .dout(new_Jinkela_wire_5173)
    );

    bfr new_Jinkela_buffer_4332 (
        .din(new_Jinkela_wire_5132),
        .dout(new_Jinkela_wire_5133)
    );

    bfr new_Jinkela_buffer_6818 (
        .din(new_Jinkela_wire_8423),
        .dout(new_Jinkela_wire_8424)
    );

    bfr new_Jinkela_buffer_6837 (
        .din(new_Jinkela_wire_8452),
        .dout(new_Jinkela_wire_8453)
    );

    bfr new_Jinkela_buffer_4333 (
        .din(new_Jinkela_wire_5133),
        .dout(new_Jinkela_wire_5134)
    );

    bfr new_Jinkela_buffer_6819 (
        .din(new_Jinkela_wire_8424),
        .dout(new_Jinkela_wire_8425)
    );

    spl4L new_Jinkela_splitter_647 (
        .a(n_0059_),
        .d(new_Jinkela_wire_8480),
        .b(new_Jinkela_wire_8481),
        .e(new_Jinkela_wire_8482),
        .c(new_Jinkela_wire_8483)
    );

    bfr new_Jinkela_buffer_4356 (
        .din(new_Jinkela_wire_5173),
        .dout(new_Jinkela_wire_5174)
    );

    bfr new_Jinkela_buffer_6838 (
        .din(new_Jinkela_wire_8453),
        .dout(new_Jinkela_wire_8454)
    );

    bfr new_Jinkela_buffer_4334 (
        .din(new_Jinkela_wire_5134),
        .dout(new_Jinkela_wire_5135)
    );

    bfr new_Jinkela_buffer_6820 (
        .din(new_Jinkela_wire_8425),
        .dout(new_Jinkela_wire_8426)
    );

    bfr new_Jinkela_buffer_4378 (
        .din(new_Jinkela_wire_5197),
        .dout(new_Jinkela_wire_5198)
    );

    spl2 new_Jinkela_splitter_649 (
        .a(n_0006_),
        .b(new_Jinkela_wire_8512),
        .c(new_Jinkela_wire_8513)
    );

    bfr new_Jinkela_buffer_4335 (
        .din(new_Jinkela_wire_5135),
        .dout(new_Jinkela_wire_5136)
    );

    bfr new_Jinkela_buffer_6821 (
        .din(new_Jinkela_wire_8426),
        .dout(new_Jinkela_wire_8427)
    );

    spl2 new_Jinkela_splitter_314 (
        .a(n_1093_),
        .b(new_Jinkela_wire_5235),
        .c(new_Jinkela_wire_5236)
    );

    spl2 new_Jinkela_splitter_648 (
        .a(n_0598_),
        .b(new_Jinkela_wire_8509),
        .c(new_Jinkela_wire_8510)
    );

    bfr new_Jinkela_buffer_4357 (
        .din(new_Jinkela_wire_5174),
        .dout(new_Jinkela_wire_5175)
    );

    bfr new_Jinkela_buffer_6839 (
        .din(new_Jinkela_wire_8454),
        .dout(new_Jinkela_wire_8455)
    );

    bfr new_Jinkela_buffer_4336 (
        .din(new_Jinkela_wire_5136),
        .dout(new_Jinkela_wire_5137)
    );

    bfr new_Jinkela_buffer_6822 (
        .din(new_Jinkela_wire_8427),
        .dout(new_Jinkela_wire_8428)
    );

    bfr new_Jinkela_buffer_6860 (
        .din(new_Jinkela_wire_8483),
        .dout(new_Jinkela_wire_8484)
    );

    bfr new_Jinkela_buffer_4337 (
        .din(new_Jinkela_wire_5137),
        .dout(new_Jinkela_wire_5138)
    );

    bfr new_Jinkela_buffer_6823 (
        .din(new_Jinkela_wire_8428),
        .dout(new_Jinkela_wire_8429)
    );

    bfr new_Jinkela_buffer_4358 (
        .din(new_Jinkela_wire_5175),
        .dout(new_Jinkela_wire_5176)
    );

    bfr new_Jinkela_buffer_4351 (
        .din(new_Jinkela_wire_5168),
        .dout(new_Jinkela_wire_5169)
    );

    bfr new_Jinkela_buffer_6840 (
        .din(new_Jinkela_wire_8455),
        .dout(new_Jinkela_wire_8456)
    );

    bfr new_Jinkela_buffer_4338 (
        .din(new_Jinkela_wire_5138),
        .dout(new_Jinkela_wire_5139)
    );

    bfr new_Jinkela_buffer_6824 (
        .din(new_Jinkela_wire_8429),
        .dout(new_Jinkela_wire_8430)
    );

    bfr new_Jinkela_buffer_4339 (
        .din(new_Jinkela_wire_5139),
        .dout(new_Jinkela_wire_5140)
    );

    bfr new_Jinkela_buffer_6825 (
        .din(new_Jinkela_wire_8430),
        .dout(new_Jinkela_wire_8431)
    );

    bfr new_Jinkela_buffer_4380 (
        .din(new_Jinkela_wire_5199),
        .dout(new_Jinkela_wire_5200)
    );

    bfr new_Jinkela_buffer_6885 (
        .din(new_Jinkela_wire_8510),
        .dout(new_Jinkela_wire_8511)
    );

    bfr new_Jinkela_buffer_4359 (
        .din(new_Jinkela_wire_5176),
        .dout(new_Jinkela_wire_5177)
    );

    bfr new_Jinkela_buffer_6841 (
        .din(new_Jinkela_wire_8456),
        .dout(new_Jinkela_wire_8457)
    );

    bfr new_Jinkela_buffer_4340 (
        .din(new_Jinkela_wire_5140),
        .dout(new_Jinkela_wire_5141)
    );

    bfr new_Jinkela_buffer_6826 (
        .din(new_Jinkela_wire_8431),
        .dout(new_Jinkela_wire_8432)
    );

    spl2 new_Jinkela_splitter_313 (
        .a(n_0275_),
        .b(new_Jinkela_wire_5232),
        .c(new_Jinkela_wire_5233)
    );

    bfr new_Jinkela_buffer_4341 (
        .din(new_Jinkela_wire_5141),
        .dout(new_Jinkela_wire_5142)
    );

    bfr new_Jinkela_buffer_6827 (
        .din(new_Jinkela_wire_8432),
        .dout(new_Jinkela_wire_8433)
    );

    bfr new_Jinkela_buffer_4399 (
        .din(new_Jinkela_wire_5233),
        .dout(new_Jinkela_wire_5234)
    );

    bfr new_Jinkela_buffer_6861 (
        .din(new_Jinkela_wire_8484),
        .dout(new_Jinkela_wire_8485)
    );

    bfr new_Jinkela_buffer_4360 (
        .din(new_Jinkela_wire_5177),
        .dout(new_Jinkela_wire_5178)
    );

    bfr new_Jinkela_buffer_6842 (
        .din(new_Jinkela_wire_8457),
        .dout(new_Jinkela_wire_8458)
    );

    bfr new_Jinkela_buffer_6828 (
        .din(new_Jinkela_wire_8433),
        .dout(new_Jinkela_wire_8434)
    );

    bfr new_Jinkela_buffer_6020 (
        .din(new_Jinkela_wire_7337),
        .dout(new_Jinkela_wire_7338)
    );

    bfr new_Jinkela_buffer_3574 (
        .din(n_0849_),
        .dout(new_Jinkela_wire_4172)
    );

    bfr new_Jinkela_buffer_3499 (
        .din(new_Jinkela_wire_4091),
        .dout(new_Jinkela_wire_4092)
    );

    spl2 new_Jinkela_splitter_516 (
        .a(n_0733_),
        .b(new_Jinkela_wire_7340),
        .c(new_Jinkela_wire_7341)
    );

    bfr new_Jinkela_buffer_6013 (
        .din(new_Jinkela_wire_7313),
        .dout(new_Jinkela_wire_7314)
    );

    bfr new_Jinkela_buffer_3490 (
        .din(new_Jinkela_wire_4066),
        .dout(new_Jinkela_wire_4067)
    );

    bfr new_Jinkela_buffer_6018 (
        .din(new_Jinkela_wire_7331),
        .dout(new_Jinkela_wire_7332)
    );

    bfr new_Jinkela_buffer_3525 (
        .din(new_Jinkela_wire_4122),
        .dout(new_Jinkela_wire_4123)
    );

    spl2 new_Jinkela_splitter_510 (
        .a(new_Jinkela_wire_7314),
        .b(new_Jinkela_wire_7315),
        .c(new_Jinkela_wire_7316)
    );

    spl2 new_Jinkela_splitter_206 (
        .a(new_Jinkela_wire_4067),
        .b(new_Jinkela_wire_4068),
        .c(new_Jinkela_wire_4069)
    );

    bfr new_Jinkela_buffer_6014 (
        .din(new_Jinkela_wire_7316),
        .dout(new_Jinkela_wire_7317)
    );

    spl2 new_Jinkela_splitter_217 (
        .a(n_0672_),
        .b(new_Jinkela_wire_4187),
        .c(new_Jinkela_wire_4188)
    );

    spl4L new_Jinkela_splitter_515 (
        .a(n_0052_),
        .d(new_Jinkela_wire_7334),
        .b(new_Jinkela_wire_7335),
        .e(new_Jinkela_wire_7336),
        .c(new_Jinkela_wire_7337)
    );

    spl3L new_Jinkela_splitter_215 (
        .a(n_0772_),
        .d(new_Jinkela_wire_4173),
        .b(new_Jinkela_wire_4174),
        .c(new_Jinkela_wire_4175)
    );

    bfr new_Jinkela_buffer_3501 (
        .din(new_Jinkela_wire_4093),
        .dout(new_Jinkela_wire_4094)
    );

    bfr new_Jinkela_buffer_6019 (
        .din(new_Jinkela_wire_7332),
        .dout(new_Jinkela_wire_7333)
    );

    bfr new_Jinkela_buffer_6015 (
        .din(new_Jinkela_wire_7317),
        .dout(new_Jinkela_wire_7318)
    );

    bfr new_Jinkela_buffer_3575 (
        .din(new_net_2552),
        .dout(new_Jinkela_wire_4176)
    );

    bfr new_Jinkela_buffer_3526 (
        .din(new_Jinkela_wire_4123),
        .dout(new_Jinkela_wire_4124)
    );

    spl3L new_Jinkela_splitter_213 (
        .a(new_Jinkela_wire_4094),
        .d(new_Jinkela_wire_4095),
        .b(new_Jinkela_wire_4096),
        .c(new_Jinkela_wire_4097)
    );

    bfr new_Jinkela_buffer_6016 (
        .din(new_Jinkela_wire_7318),
        .dout(new_Jinkela_wire_7319)
    );

    bfr new_Jinkela_buffer_3502 (
        .din(new_Jinkela_wire_4097),
        .dout(new_Jinkela_wire_4098)
    );

    bfr new_Jinkela_buffer_6022 (
        .din(n_1060_),
        .dout(new_Jinkela_wire_7342)
    );

    spl2 new_Jinkela_splitter_511 (
        .a(new_Jinkela_wire_7319),
        .b(new_Jinkela_wire_7320),
        .c(new_Jinkela_wire_7321)
    );

    bfr new_Jinkela_buffer_3576 (
        .din(n_0101_),
        .dout(new_Jinkela_wire_4177)
    );

    bfr new_Jinkela_buffer_3527 (
        .din(new_Jinkela_wire_4124),
        .dout(new_Jinkela_wire_4125)
    );

    bfr new_Jinkela_buffer_3503 (
        .din(new_Jinkela_wire_4098),
        .dout(new_Jinkela_wire_4099)
    );

    bfr new_Jinkela_buffer_6021 (
        .din(new_Jinkela_wire_7338),
        .dout(new_Jinkela_wire_7339)
    );

    bfr new_Jinkela_buffer_6025 (
        .din(n_1251_),
        .dout(new_Jinkela_wire_7347)
    );

    bfr new_Jinkela_buffer_3504 (
        .din(new_Jinkela_wire_4099),
        .dout(new_Jinkela_wire_4100)
    );

    bfr new_Jinkela_buffer_6023 (
        .din(new_Jinkela_wire_7342),
        .dout(new_Jinkela_wire_7343)
    );

    bfr new_Jinkela_buffer_3528 (
        .din(new_Jinkela_wire_4125),
        .dout(new_Jinkela_wire_4126)
    );

    bfr new_Jinkela_buffer_6033 (
        .din(n_0770_),
        .dout(new_Jinkela_wire_7359)
    );

    spl2 new_Jinkela_splitter_519 (
        .a(n_0696_),
        .b(new_Jinkela_wire_7352),
        .c(new_Jinkela_wire_7353)
    );

    bfr new_Jinkela_buffer_3500 (
        .din(new_Jinkela_wire_4092),
        .dout(new_Jinkela_wire_4093)
    );

    bfr new_Jinkela_buffer_3505 (
        .din(new_Jinkela_wire_4100),
        .dout(new_Jinkela_wire_4101)
    );

    bfr new_Jinkela_buffer_6024 (
        .din(new_Jinkela_wire_7343),
        .dout(new_Jinkela_wire_7344)
    );

    bfr new_Jinkela_buffer_6026 (
        .din(new_Jinkela_wire_7347),
        .dout(new_Jinkela_wire_7348)
    );

    spl2 new_Jinkela_splitter_216 (
        .a(n_0051_),
        .b(new_Jinkela_wire_4181),
        .c(new_Jinkela_wire_4182)
    );

    bfr new_Jinkela_buffer_3506 (
        .din(new_Jinkela_wire_4101),
        .dout(new_Jinkela_wire_4102)
    );

    spl2 new_Jinkela_splitter_517 (
        .a(new_Jinkela_wire_7344),
        .b(new_Jinkela_wire_7345),
        .c(new_Jinkela_wire_7346)
    );

    bfr new_Jinkela_buffer_6027 (
        .din(new_Jinkela_wire_7348),
        .dout(new_Jinkela_wire_7349)
    );

    bfr new_Jinkela_buffer_3529 (
        .din(new_Jinkela_wire_4126),
        .dout(new_Jinkela_wire_4127)
    );

    bfr new_Jinkela_buffer_3507 (
        .din(new_Jinkela_wire_4102),
        .dout(new_Jinkela_wire_4103)
    );

    bfr new_Jinkela_buffer_6036 (
        .din(n_0257_),
        .dout(new_Jinkela_wire_7364)
    );

    bfr new_Jinkela_buffer_6028 (
        .din(new_Jinkela_wire_7353),
        .dout(new_Jinkela_wire_7354)
    );

    bfr new_Jinkela_buffer_3577 (
        .din(new_Jinkela_wire_4177),
        .dout(new_Jinkela_wire_4178)
    );

    bfr new_Jinkela_buffer_3508 (
        .din(new_Jinkela_wire_4103),
        .dout(new_Jinkela_wire_4104)
    );

    spl2 new_Jinkela_splitter_518 (
        .a(new_Jinkela_wire_7349),
        .b(new_Jinkela_wire_7350),
        .c(new_Jinkela_wire_7351)
    );

    bfr new_Jinkela_buffer_6029 (
        .din(new_Jinkela_wire_7354),
        .dout(new_Jinkela_wire_7355)
    );

    bfr new_Jinkela_buffer_3530 (
        .din(new_Jinkela_wire_4127),
        .dout(new_Jinkela_wire_4128)
    );

    bfr new_Jinkela_buffer_3509 (
        .din(new_Jinkela_wire_4104),
        .dout(new_Jinkela_wire_4105)
    );

    spl2 new_Jinkela_splitter_521 (
        .a(n_0682_),
        .b(new_Jinkela_wire_7370),
        .c(new_Jinkela_wire_7371)
    );

    bfr new_Jinkela_buffer_6034 (
        .din(new_Jinkela_wire_7359),
        .dout(new_Jinkela_wire_7360)
    );

    spl2 new_Jinkela_splitter_522 (
        .a(n_1342_),
        .b(new_Jinkela_wire_7372),
        .c(new_Jinkela_wire_7373)
    );

    bfr new_Jinkela_buffer_3580 (
        .din(new_Jinkela_wire_4182),
        .dout(new_Jinkela_wire_4183)
    );

    bfr new_Jinkela_buffer_3510 (
        .din(new_Jinkela_wire_4105),
        .dout(new_Jinkela_wire_4106)
    );

    bfr new_Jinkela_buffer_6030 (
        .din(new_Jinkela_wire_7355),
        .dout(new_Jinkela_wire_7356)
    );

    bfr new_Jinkela_buffer_6037 (
        .din(new_Jinkela_wire_7364),
        .dout(new_Jinkela_wire_7365)
    );

    bfr new_Jinkela_buffer_3531 (
        .din(new_Jinkela_wire_4128),
        .dout(new_Jinkela_wire_4129)
    );

    bfr new_Jinkela_buffer_3511 (
        .din(new_Jinkela_wire_4106),
        .dout(new_Jinkela_wire_4107)
    );

    bfr new_Jinkela_buffer_6031 (
        .din(new_Jinkela_wire_7356),
        .dout(new_Jinkela_wire_7357)
    );

    bfr new_Jinkela_buffer_6035 (
        .din(new_Jinkela_wire_7360),
        .dout(new_Jinkela_wire_7361)
    );

    bfr new_Jinkela_buffer_3578 (
        .din(new_Jinkela_wire_4178),
        .dout(new_Jinkela_wire_4179)
    );

    bfr new_Jinkela_buffer_3512 (
        .din(new_Jinkela_wire_4107),
        .dout(new_Jinkela_wire_4108)
    );

    bfr new_Jinkela_buffer_6032 (
        .din(new_Jinkela_wire_7357),
        .dout(new_Jinkela_wire_7358)
    );

    bfr new_Jinkela_buffer_3532 (
        .din(new_Jinkela_wire_4129),
        .dout(new_Jinkela_wire_4130)
    );

    bfr new_Jinkela_buffer_3513 (
        .din(new_Jinkela_wire_4108),
        .dout(new_Jinkela_wire_4109)
    );

    spl2 new_Jinkela_splitter_520 (
        .a(new_Jinkela_wire_7361),
        .b(new_Jinkela_wire_7362),
        .c(new_Jinkela_wire_7363)
    );

    bfr new_Jinkela_buffer_3514 (
        .din(new_Jinkela_wire_4109),
        .dout(new_Jinkela_wire_4110)
    );

    bfr new_Jinkela_buffer_6051 (
        .din(n_0397_),
        .dout(new_Jinkela_wire_7385)
    );

    bfr new_Jinkela_buffer_6038 (
        .din(new_Jinkela_wire_7365),
        .dout(new_Jinkela_wire_7366)
    );

    bfr new_Jinkela_buffer_6039 (
        .din(new_Jinkela_wire_7366),
        .dout(new_Jinkela_wire_7367)
    );

    bfr new_Jinkela_buffer_3533 (
        .din(new_Jinkela_wire_4130),
        .dout(new_Jinkela_wire_4131)
    );

    bfr new_Jinkela_buffer_3515 (
        .din(new_Jinkela_wire_4110),
        .dout(new_Jinkela_wire_4111)
    );

    spl2 new_Jinkela_splitter_523 (
        .a(n_1183_),
        .b(new_Jinkela_wire_7383),
        .c(new_Jinkela_wire_7384)
    );

    bfr new_Jinkela_buffer_6042 (
        .din(new_Jinkela_wire_7373),
        .dout(new_Jinkela_wire_7374)
    );

    bfr new_Jinkela_buffer_6040 (
        .din(new_Jinkela_wire_7367),
        .dout(new_Jinkela_wire_7368)
    );

    bfr new_Jinkela_buffer_3579 (
        .din(new_Jinkela_wire_4179),
        .dout(new_Jinkela_wire_4180)
    );

    bfr new_Jinkela_buffer_3516 (
        .din(new_Jinkela_wire_4111),
        .dout(new_Jinkela_wire_4112)
    );

    bfr new_Jinkela_buffer_6052 (
        .din(n_0574_),
        .dout(new_Jinkela_wire_7386)
    );

    bfr new_Jinkela_buffer_6041 (
        .din(new_Jinkela_wire_7368),
        .dout(new_Jinkela_wire_7369)
    );

    bfr new_Jinkela_buffer_3534 (
        .din(new_Jinkela_wire_4131),
        .dout(new_Jinkela_wire_4132)
    );

    bfr new_Jinkela_buffer_3517 (
        .din(new_Jinkela_wire_4112),
        .dout(new_Jinkela_wire_4113)
    );

    bfr new_Jinkela_buffer_6043 (
        .din(new_Jinkela_wire_7374),
        .dout(new_Jinkela_wire_7375)
    );

    bfr new_Jinkela_buffer_2083 (
        .din(new_Jinkela_wire_2452),
        .dout(new_Jinkela_wire_2453)
    );

    bfr new_Jinkela_buffer_422 (
        .din(new_Jinkela_wire_458),
        .dout(new_Jinkela_wire_459)
    );

    bfr new_Jinkela_buffer_376 (
        .din(new_Jinkela_wire_407),
        .dout(new_Jinkela_wire_408)
    );

    bfr new_Jinkela_buffer_1918 (
        .din(new_Jinkela_wire_2278),
        .dout(new_Jinkela_wire_2279)
    );

    bfr new_Jinkela_buffer_5192 (
        .din(new_Jinkela_wire_6213),
        .dout(new_Jinkela_wire_6214)
    );

    bfr new_Jinkela_buffer_1963 (
        .din(new_Jinkela_wire_2327),
        .dout(new_Jinkela_wire_2328)
    );

    bfr new_Jinkela_buffer_549 (
        .din(N109),
        .dout(new_Jinkela_wire_591)
    );

    bfr new_Jinkela_buffer_5273 (
        .din(n_0594_),
        .dout(new_Jinkela_wire_6310)
    );

    bfr new_Jinkela_buffer_377 (
        .din(new_Jinkela_wire_408),
        .dout(new_Jinkela_wire_409)
    );

    bfr new_Jinkela_buffer_1919 (
        .din(new_Jinkela_wire_2279),
        .dout(new_Jinkela_wire_2280)
    );

    bfr new_Jinkela_buffer_5193 (
        .din(new_Jinkela_wire_6214),
        .dout(new_Jinkela_wire_6215)
    );

    bfr new_Jinkela_buffer_5229 (
        .din(new_Jinkela_wire_6256),
        .dout(new_Jinkela_wire_6257)
    );

    bfr new_Jinkela_buffer_2019 (
        .din(new_Jinkela_wire_2388),
        .dout(new_Jinkela_wire_2389)
    );

    bfr new_Jinkela_buffer_423 (
        .din(new_Jinkela_wire_459),
        .dout(new_Jinkela_wire_460)
    );

    bfr new_Jinkela_buffer_378 (
        .din(new_Jinkela_wire_409),
        .dout(new_Jinkela_wire_410)
    );

    bfr new_Jinkela_buffer_1920 (
        .din(new_Jinkela_wire_2280),
        .dout(new_Jinkela_wire_2281)
    );

    bfr new_Jinkela_buffer_5194 (
        .din(new_Jinkela_wire_6215),
        .dout(new_Jinkela_wire_6216)
    );

    spl2 new_Jinkela_splitter_399 (
        .a(n_0474_),
        .b(new_Jinkela_wire_6308),
        .c(new_Jinkela_wire_6309)
    );

    bfr new_Jinkela_buffer_1964 (
        .din(new_Jinkela_wire_2328),
        .dout(new_Jinkela_wire_2329)
    );

    spl3L new_Jinkela_splitter_17 (
        .a(new_Jinkela_wire_519),
        .d(new_Jinkela_wire_520),
        .b(new_Jinkela_wire_521),
        .c(new_Jinkela_wire_522)
    );

    bfr new_Jinkela_buffer_5232 (
        .din(new_Jinkela_wire_6266),
        .dout(new_Jinkela_wire_6267)
    );

    bfr new_Jinkela_buffer_379 (
        .din(new_Jinkela_wire_410),
        .dout(new_Jinkela_wire_411)
    );

    bfr new_Jinkela_buffer_1921 (
        .din(new_Jinkela_wire_2281),
        .dout(new_Jinkela_wire_2282)
    );

    bfr new_Jinkela_buffer_5195 (
        .din(new_Jinkela_wire_6216),
        .dout(new_Jinkela_wire_6217)
    );

    bfr new_Jinkela_buffer_5230 (
        .din(new_Jinkela_wire_6257),
        .dout(new_Jinkela_wire_6258)
    );

    bfr new_Jinkela_buffer_2086 (
        .din(new_Jinkela_wire_2455),
        .dout(new_Jinkela_wire_2456)
    );

    bfr new_Jinkela_buffer_424 (
        .din(new_Jinkela_wire_460),
        .dout(new_Jinkela_wire_461)
    );

    bfr new_Jinkela_buffer_380 (
        .din(new_Jinkela_wire_411),
        .dout(new_Jinkela_wire_412)
    );

    bfr new_Jinkela_buffer_1922 (
        .din(new_Jinkela_wire_2282),
        .dout(new_Jinkela_wire_2283)
    );

    bfr new_Jinkela_buffer_5196 (
        .din(new_Jinkela_wire_6217),
        .dout(new_Jinkela_wire_6218)
    );

    bfr new_Jinkela_buffer_1965 (
        .din(new_Jinkela_wire_2329),
        .dout(new_Jinkela_wire_2330)
    );

    bfr new_Jinkela_buffer_546 (
        .din(new_Jinkela_wire_587),
        .dout(new_Jinkela_wire_588)
    );

    spl2 new_Jinkela_splitter_401 (
        .a(n_0695_),
        .b(new_Jinkela_wire_6315),
        .c(new_Jinkela_wire_6316)
    );

    bfr new_Jinkela_buffer_381 (
        .din(new_Jinkela_wire_412),
        .dout(new_Jinkela_wire_413)
    );

    bfr new_Jinkela_buffer_1923 (
        .din(new_Jinkela_wire_2283),
        .dout(new_Jinkela_wire_2284)
    );

    bfr new_Jinkela_buffer_5197 (
        .din(new_Jinkela_wire_6218),
        .dout(new_Jinkela_wire_6219)
    );

    spl2 new_Jinkela_splitter_396 (
        .a(new_Jinkela_wire_6258),
        .b(new_Jinkela_wire_6259),
        .c(new_Jinkela_wire_6260)
    );

    bfr new_Jinkela_buffer_2020 (
        .din(new_Jinkela_wire_2389),
        .dout(new_Jinkela_wire_2390)
    );

    bfr new_Jinkela_buffer_425 (
        .din(new_Jinkela_wire_461),
        .dout(new_Jinkela_wire_462)
    );

    bfr new_Jinkela_buffer_382 (
        .din(new_Jinkela_wire_413),
        .dout(new_Jinkela_wire_414)
    );

    bfr new_Jinkela_buffer_1924 (
        .din(new_Jinkela_wire_2284),
        .dout(new_Jinkela_wire_2285)
    );

    bfr new_Jinkela_buffer_5198 (
        .din(new_Jinkela_wire_6219),
        .dout(new_Jinkela_wire_6220)
    );

    bfr new_Jinkela_buffer_1966 (
        .din(new_Jinkela_wire_2330),
        .dout(new_Jinkela_wire_2331)
    );

    bfr new_Jinkela_buffer_481 (
        .din(new_Jinkela_wire_522),
        .dout(new_Jinkela_wire_523)
    );

    bfr new_Jinkela_buffer_383 (
        .din(new_Jinkela_wire_414),
        .dout(new_Jinkela_wire_415)
    );

    bfr new_Jinkela_buffer_1925 (
        .din(new_Jinkela_wire_2285),
        .dout(new_Jinkela_wire_2286)
    );

    bfr new_Jinkela_buffer_5199 (
        .din(new_Jinkela_wire_6220),
        .dout(new_Jinkela_wire_6221)
    );

    bfr new_Jinkela_buffer_5274 (
        .din(new_Jinkela_wire_6310),
        .dout(new_Jinkela_wire_6311)
    );

    bfr new_Jinkela_buffer_2084 (
        .din(new_Jinkela_wire_2453),
        .dout(new_Jinkela_wire_2454)
    );

    bfr new_Jinkela_buffer_426 (
        .din(new_Jinkela_wire_462),
        .dout(new_Jinkela_wire_463)
    );

    bfr new_Jinkela_buffer_5233 (
        .din(new_Jinkela_wire_6267),
        .dout(new_Jinkela_wire_6268)
    );

    bfr new_Jinkela_buffer_384 (
        .din(new_Jinkela_wire_415),
        .dout(new_Jinkela_wire_416)
    );

    bfr new_Jinkela_buffer_1926 (
        .din(new_Jinkela_wire_2286),
        .dout(new_Jinkela_wire_2287)
    );

    bfr new_Jinkela_buffer_5200 (
        .din(new_Jinkela_wire_6221),
        .dout(new_Jinkela_wire_6222)
    );

    bfr new_Jinkela_buffer_1967 (
        .din(new_Jinkela_wire_2331),
        .dout(new_Jinkela_wire_2332)
    );

    bfr new_Jinkela_buffer_553 (
        .din(N97),
        .dout(new_Jinkela_wire_595)
    );

    bfr new_Jinkela_buffer_5234 (
        .din(new_Jinkela_wire_6268),
        .dout(new_Jinkela_wire_6269)
    );

    bfr new_Jinkela_buffer_385 (
        .din(new_Jinkela_wire_416),
        .dout(new_Jinkela_wire_417)
    );

    bfr new_Jinkela_buffer_1927 (
        .din(new_Jinkela_wire_2287),
        .dout(new_Jinkela_wire_2288)
    );

    bfr new_Jinkela_buffer_5201 (
        .din(new_Jinkela_wire_6222),
        .dout(new_Jinkela_wire_6223)
    );

    bfr new_Jinkela_buffer_2021 (
        .din(new_Jinkela_wire_2390),
        .dout(new_Jinkela_wire_2391)
    );

    bfr new_Jinkela_buffer_427 (
        .din(new_Jinkela_wire_463),
        .dout(new_Jinkela_wire_464)
    );

    spl3L new_Jinkela_splitter_400 (
        .a(n_1206_),
        .d(new_Jinkela_wire_6312),
        .b(new_Jinkela_wire_6313),
        .c(new_Jinkela_wire_6314)
    );

    bfr new_Jinkela_buffer_386 (
        .din(new_Jinkela_wire_417),
        .dout(new_Jinkela_wire_418)
    );

    bfr new_Jinkela_buffer_1928 (
        .din(new_Jinkela_wire_2288),
        .dout(new_Jinkela_wire_2289)
    );

    bfr new_Jinkela_buffer_5202 (
        .din(new_Jinkela_wire_6223),
        .dout(new_Jinkela_wire_6224)
    );

    bfr new_Jinkela_buffer_1968 (
        .din(new_Jinkela_wire_2332),
        .dout(new_Jinkela_wire_2333)
    );

    bfr new_Jinkela_buffer_482 (
        .din(new_Jinkela_wire_523),
        .dout(new_Jinkela_wire_524)
    );

    bfr new_Jinkela_buffer_5235 (
        .din(new_Jinkela_wire_6269),
        .dout(new_Jinkela_wire_6270)
    );

    bfr new_Jinkela_buffer_387 (
        .din(new_Jinkela_wire_418),
        .dout(new_Jinkela_wire_419)
    );

    bfr new_Jinkela_buffer_1929 (
        .din(new_Jinkela_wire_2289),
        .dout(new_Jinkela_wire_2290)
    );

    bfr new_Jinkela_buffer_5203 (
        .din(new_Jinkela_wire_6224),
        .dout(new_Jinkela_wire_6225)
    );

    bfr new_Jinkela_buffer_2093 (
        .din(N153),
        .dout(new_Jinkela_wire_2463)
    );

    bfr new_Jinkela_buffer_428 (
        .din(new_Jinkela_wire_464),
        .dout(new_Jinkela_wire_465)
    );

    spl2 new_Jinkela_splitter_402 (
        .a(n_0719_),
        .b(new_Jinkela_wire_6317),
        .c(new_Jinkela_wire_6318)
    );

    bfr new_Jinkela_buffer_388 (
        .din(new_Jinkela_wire_419),
        .dout(new_Jinkela_wire_420)
    );

    bfr new_Jinkela_buffer_1930 (
        .din(new_Jinkela_wire_2290),
        .dout(new_Jinkela_wire_2291)
    );

    bfr new_Jinkela_buffer_5204 (
        .din(new_Jinkela_wire_6225),
        .dout(new_Jinkela_wire_6226)
    );

    bfr new_Jinkela_buffer_1969 (
        .din(new_Jinkela_wire_2333),
        .dout(new_Jinkela_wire_2334)
    );

    bfr new_Jinkela_buffer_547 (
        .din(new_Jinkela_wire_588),
        .dout(new_Jinkela_wire_589)
    );

    bfr new_Jinkela_buffer_5236 (
        .din(new_Jinkela_wire_6270),
        .dout(new_Jinkela_wire_6271)
    );

    bfr new_Jinkela_buffer_389 (
        .din(new_Jinkela_wire_420),
        .dout(new_Jinkela_wire_421)
    );

    bfr new_Jinkela_buffer_1931 (
        .din(new_Jinkela_wire_2291),
        .dout(new_Jinkela_wire_2292)
    );

    bfr new_Jinkela_buffer_5205 (
        .din(new_Jinkela_wire_6226),
        .dout(new_Jinkela_wire_6227)
    );

    bfr new_Jinkela_buffer_2022 (
        .din(new_Jinkela_wire_2391),
        .dout(new_Jinkela_wire_2392)
    );

    bfr new_Jinkela_buffer_429 (
        .din(new_Jinkela_wire_465),
        .dout(new_Jinkela_wire_466)
    );

    bfr new_Jinkela_buffer_390 (
        .din(new_Jinkela_wire_421),
        .dout(new_Jinkela_wire_422)
    );

    bfr new_Jinkela_buffer_1932 (
        .din(new_Jinkela_wire_2292),
        .dout(new_Jinkela_wire_2293)
    );

    bfr new_Jinkela_buffer_5206 (
        .din(new_Jinkela_wire_6227),
        .dout(new_Jinkela_wire_6228)
    );

    bfr new_Jinkela_buffer_1970 (
        .din(new_Jinkela_wire_2334),
        .dout(new_Jinkela_wire_2335)
    );

    bfr new_Jinkela_buffer_483 (
        .din(new_Jinkela_wire_524),
        .dout(new_Jinkela_wire_525)
    );

    bfr new_Jinkela_buffer_5237 (
        .din(new_Jinkela_wire_6271),
        .dout(new_Jinkela_wire_6272)
    );

    bfr new_Jinkela_buffer_391 (
        .din(new_Jinkela_wire_422),
        .dout(new_Jinkela_wire_423)
    );

    bfr new_Jinkela_buffer_1933 (
        .din(new_Jinkela_wire_2293),
        .dout(new_Jinkela_wire_2294)
    );

    bfr new_Jinkela_buffer_5207 (
        .din(new_Jinkela_wire_6228),
        .dout(new_Jinkela_wire_6229)
    );

    bfr new_Jinkela_buffer_2087 (
        .din(new_Jinkela_wire_2456),
        .dout(new_Jinkela_wire_2457)
    );

    bfr new_Jinkela_buffer_430 (
        .din(new_Jinkela_wire_466),
        .dout(new_Jinkela_wire_467)
    );

    bfr new_Jinkela_buffer_392 (
        .din(new_Jinkela_wire_423),
        .dout(new_Jinkela_wire_424)
    );

    bfr new_Jinkela_buffer_1934 (
        .din(new_Jinkela_wire_2294),
        .dout(new_Jinkela_wire_2295)
    );

    bfr new_Jinkela_buffer_5208 (
        .din(new_Jinkela_wire_6229),
        .dout(new_Jinkela_wire_6230)
    );

    bfr new_Jinkela_buffer_1971 (
        .din(new_Jinkela_wire_2335),
        .dout(new_Jinkela_wire_2336)
    );

    bfr new_Jinkela_buffer_550 (
        .din(new_Jinkela_wire_591),
        .dout(new_Jinkela_wire_592)
    );

    bfr new_Jinkela_buffer_5238 (
        .din(new_Jinkela_wire_6272),
        .dout(new_Jinkela_wire_6273)
    );

    bfr new_Jinkela_buffer_393 (
        .din(new_Jinkela_wire_424),
        .dout(new_Jinkela_wire_425)
    );

    bfr new_Jinkela_buffer_1935 (
        .din(new_Jinkela_wire_2295),
        .dout(new_Jinkela_wire_2296)
    );

    bfr new_Jinkela_buffer_5209 (
        .din(new_Jinkela_wire_6230),
        .dout(new_Jinkela_wire_6231)
    );

    bfr new_Jinkela_buffer_2023 (
        .din(new_Jinkela_wire_2392),
        .dout(new_Jinkela_wire_2393)
    );

    bfr new_Jinkela_buffer_431 (
        .din(new_Jinkela_wire_467),
        .dout(new_Jinkela_wire_468)
    );

    spl2 new_Jinkela_splitter_403 (
        .a(n_0639_),
        .b(new_Jinkela_wire_6321),
        .c(new_Jinkela_wire_6322)
    );

    bfr new_Jinkela_buffer_394 (
        .din(new_Jinkela_wire_425),
        .dout(new_Jinkela_wire_426)
    );

    bfr new_Jinkela_buffer_1936 (
        .din(new_Jinkela_wire_2296),
        .dout(new_Jinkela_wire_2297)
    );

    bfr new_Jinkela_buffer_5210 (
        .din(new_Jinkela_wire_6231),
        .dout(new_Jinkela_wire_6232)
    );

    bfr new_Jinkela_buffer_5275 (
        .din(new_Jinkela_wire_6318),
        .dout(new_Jinkela_wire_6319)
    );

    bfr new_Jinkela_buffer_1972 (
        .din(new_Jinkela_wire_2336),
        .dout(new_Jinkela_wire_2337)
    );

    bfr new_Jinkela_buffer_484 (
        .din(new_Jinkela_wire_525),
        .dout(new_Jinkela_wire_526)
    );

    bfr new_Jinkela_buffer_5239 (
        .din(new_Jinkela_wire_6273),
        .dout(new_Jinkela_wire_6274)
    );

    bfr new_Jinkela_buffer_1937 (
        .din(new_Jinkela_wire_2297),
        .dout(new_Jinkela_wire_2298)
    );

    bfr new_Jinkela_buffer_5211 (
        .din(new_Jinkela_wire_6232),
        .dout(new_Jinkela_wire_6233)
    );

    bfr new_Jinkela_buffer_432 (
        .din(new_Jinkela_wire_468),
        .dout(new_Jinkela_wire_469)
    );

    bfr new_Jinkela_buffer_2090 (
        .din(new_Jinkela_wire_2459),
        .dout(new_Jinkela_wire_2460)
    );

    bfr new_Jinkela_buffer_548 (
        .din(new_Jinkela_wire_589),
        .dout(new_Jinkela_wire_590)
    );

    bfr new_Jinkela_buffer_5277 (
        .din(n_0831_),
        .dout(new_Jinkela_wire_6323)
    );

    bfr new_Jinkela_buffer_1938 (
        .din(new_Jinkela_wire_2298),
        .dout(new_Jinkela_wire_2299)
    );

    bfr new_Jinkela_buffer_5212 (
        .din(new_Jinkela_wire_6233),
        .dout(new_Jinkela_wire_6234)
    );

    bfr new_Jinkela_buffer_433 (
        .din(new_Jinkela_wire_469),
        .dout(new_Jinkela_wire_470)
    );

    spl2 new_Jinkela_splitter_640 (
        .a(new_Jinkela_wire_8434),
        .b(new_Jinkela_wire_8435),
        .c(new_Jinkela_wire_8436)
    );

    spl3L new_Jinkela_splitter_650 (
        .a(n_1353_),
        .d(new_Jinkela_wire_8514),
        .b(new_Jinkela_wire_8515),
        .c(new_Jinkela_wire_8516)
    );

    bfr new_Jinkela_buffer_6843 (
        .din(new_Jinkela_wire_8458),
        .dout(new_Jinkela_wire_8459)
    );

    bfr new_Jinkela_buffer_6862 (
        .din(new_Jinkela_wire_8485),
        .dout(new_Jinkela_wire_8486)
    );

    bfr new_Jinkela_buffer_6844 (
        .din(new_Jinkela_wire_8459),
        .dout(new_Jinkela_wire_8460)
    );

    bfr new_Jinkela_buffer_6886 (
        .din(new_Jinkela_wire_8516),
        .dout(new_Jinkela_wire_8517)
    );

    bfr new_Jinkela_buffer_6845 (
        .din(new_Jinkela_wire_8460),
        .dout(new_Jinkela_wire_8461)
    );

    bfr new_Jinkela_buffer_6863 (
        .din(new_Jinkela_wire_8486),
        .dout(new_Jinkela_wire_8487)
    );

    bfr new_Jinkela_buffer_6846 (
        .din(new_Jinkela_wire_8461),
        .dout(new_Jinkela_wire_8462)
    );

    bfr new_Jinkela_buffer_6909 (
        .din(n_0448_),
        .dout(new_Jinkela_wire_8540)
    );

    bfr new_Jinkela_buffer_6847 (
        .din(new_Jinkela_wire_8462),
        .dout(new_Jinkela_wire_8463)
    );

    bfr new_Jinkela_buffer_6902 (
        .din(n_0483_),
        .dout(new_Jinkela_wire_8533)
    );

    bfr new_Jinkela_buffer_6864 (
        .din(new_Jinkela_wire_8487),
        .dout(new_Jinkela_wire_8488)
    );

    bfr new_Jinkela_buffer_6848 (
        .din(new_Jinkela_wire_8463),
        .dout(new_Jinkela_wire_8464)
    );

    bfr new_Jinkela_buffer_6849 (
        .din(new_Jinkela_wire_8464),
        .dout(new_Jinkela_wire_8465)
    );

    bfr new_Jinkela_buffer_6903 (
        .din(new_Jinkela_wire_8533),
        .dout(new_Jinkela_wire_8534)
    );

    bfr new_Jinkela_buffer_6865 (
        .din(new_Jinkela_wire_8488),
        .dout(new_Jinkela_wire_8489)
    );

    bfr new_Jinkela_buffer_6850 (
        .din(new_Jinkela_wire_8465),
        .dout(new_Jinkela_wire_8466)
    );

    bfr new_Jinkela_buffer_6851 (
        .din(new_Jinkela_wire_8466),
        .dout(new_Jinkela_wire_8467)
    );

    bfr new_Jinkela_buffer_6866 (
        .din(new_Jinkela_wire_8489),
        .dout(new_Jinkela_wire_8490)
    );

    bfr new_Jinkela_buffer_6852 (
        .din(new_Jinkela_wire_8467),
        .dout(new_Jinkela_wire_8468)
    );

    bfr new_Jinkela_buffer_6887 (
        .din(new_Jinkela_wire_8517),
        .dout(new_Jinkela_wire_8518)
    );

    bfr new_Jinkela_buffer_6853 (
        .din(new_Jinkela_wire_8468),
        .dout(new_Jinkela_wire_8469)
    );

    bfr new_Jinkela_buffer_6867 (
        .din(new_Jinkela_wire_8490),
        .dout(new_Jinkela_wire_8491)
    );

    bfr new_Jinkela_buffer_6854 (
        .din(new_Jinkela_wire_8469),
        .dout(new_Jinkela_wire_8470)
    );

    bfr new_Jinkela_buffer_6855 (
        .din(new_Jinkela_wire_8470),
        .dout(new_Jinkela_wire_8471)
    );

    spl2 new_Jinkela_splitter_651 (
        .a(n_0035_),
        .b(new_Jinkela_wire_8567),
        .c(new_Jinkela_wire_8568)
    );

    bfr new_Jinkela_buffer_6868 (
        .din(new_Jinkela_wire_8491),
        .dout(new_Jinkela_wire_8492)
    );

    bfr new_Jinkela_buffer_6856 (
        .din(new_Jinkela_wire_8471),
        .dout(new_Jinkela_wire_8472)
    );

    bfr new_Jinkela_buffer_6888 (
        .din(new_Jinkela_wire_8518),
        .dout(new_Jinkela_wire_8519)
    );

    bfr new_Jinkela_buffer_6857 (
        .din(new_Jinkela_wire_8472),
        .dout(new_Jinkela_wire_8473)
    );

    bfr new_Jinkela_buffer_6869 (
        .din(new_Jinkela_wire_8492),
        .dout(new_Jinkela_wire_8493)
    );

    bfr new_Jinkela_buffer_6858 (
        .din(new_Jinkela_wire_8473),
        .dout(new_Jinkela_wire_8474)
    );

    bfr new_Jinkela_buffer_6936 (
        .din(n_0236_),
        .dout(new_Jinkela_wire_8569)
    );

    bfr new_Jinkela_buffer_6859 (
        .din(new_Jinkela_wire_8474),
        .dout(new_Jinkela_wire_8475)
    );

    bfr new_Jinkela_buffer_6904 (
        .din(new_Jinkela_wire_8534),
        .dout(new_Jinkela_wire_8535)
    );

    bfr new_Jinkela_buffer_6870 (
        .din(new_Jinkela_wire_8493),
        .dout(new_Jinkela_wire_8494)
    );

    bfr new_Jinkela_buffer_6889 (
        .din(new_Jinkela_wire_8519),
        .dout(new_Jinkela_wire_8520)
    );

    bfr new_Jinkela_buffer_6871 (
        .din(new_Jinkela_wire_8494),
        .dout(new_Jinkela_wire_8495)
    );

    bfr new_Jinkela_buffer_6910 (
        .din(new_Jinkela_wire_8540),
        .dout(new_Jinkela_wire_8541)
    );

    bfr new_Jinkela_buffer_6872 (
        .din(new_Jinkela_wire_8495),
        .dout(new_Jinkela_wire_8496)
    );

    bfr new_Jinkela_buffer_6890 (
        .din(new_Jinkela_wire_8520),
        .dout(new_Jinkela_wire_8521)
    );

    bfr new_Jinkela_buffer_2669 (
        .din(new_Jinkela_wire_3078),
        .dout(new_Jinkela_wire_3079)
    );

    bfr new_Jinkela_buffer_2634 (
        .din(new_Jinkela_wire_3039),
        .dout(new_Jinkela_wire_3040)
    );

    bfr new_Jinkela_buffer_2721 (
        .din(new_Jinkela_wire_3135),
        .dout(new_Jinkela_wire_3136)
    );

    bfr new_Jinkela_buffer_2635 (
        .din(new_Jinkela_wire_3040),
        .dout(new_Jinkela_wire_3041)
    );

    bfr new_Jinkela_buffer_2670 (
        .din(new_Jinkela_wire_3079),
        .dout(new_Jinkela_wire_3080)
    );

    bfr new_Jinkela_buffer_2636 (
        .din(new_Jinkela_wire_3041),
        .dout(new_Jinkela_wire_3042)
    );

    bfr new_Jinkela_buffer_2851 (
        .din(new_Jinkela_wire_3272),
        .dout(new_Jinkela_wire_3273)
    );

    bfr new_Jinkela_buffer_2637 (
        .din(new_Jinkela_wire_3042),
        .dout(new_Jinkela_wire_3043)
    );

    bfr new_Jinkela_buffer_2915 (
        .din(N138),
        .dout(new_Jinkela_wire_3339)
    );

    bfr new_Jinkela_buffer_2671 (
        .din(new_Jinkela_wire_3080),
        .dout(new_Jinkela_wire_3081)
    );

    bfr new_Jinkela_buffer_2638 (
        .din(new_Jinkela_wire_3043),
        .dout(new_Jinkela_wire_3044)
    );

    bfr new_Jinkela_buffer_2722 (
        .din(new_Jinkela_wire_3136),
        .dout(new_Jinkela_wire_3137)
    );

    bfr new_Jinkela_buffer_2672 (
        .din(new_Jinkela_wire_3081),
        .dout(new_Jinkela_wire_3082)
    );

    bfr new_Jinkela_buffer_2786 (
        .din(new_Jinkela_wire_3200),
        .dout(new_Jinkela_wire_3201)
    );

    bfr new_Jinkela_buffer_2673 (
        .din(new_Jinkela_wire_3082),
        .dout(new_Jinkela_wire_3083)
    );

    bfr new_Jinkela_buffer_2723 (
        .din(new_Jinkela_wire_3137),
        .dout(new_Jinkela_wire_3138)
    );

    bfr new_Jinkela_buffer_2674 (
        .din(new_Jinkela_wire_3083),
        .dout(new_Jinkela_wire_3084)
    );

    bfr new_Jinkela_buffer_2675 (
        .din(new_Jinkela_wire_3084),
        .dout(new_Jinkela_wire_3085)
    );

    bfr new_Jinkela_buffer_2724 (
        .din(new_Jinkela_wire_3138),
        .dout(new_Jinkela_wire_3139)
    );

    bfr new_Jinkela_buffer_2676 (
        .din(new_Jinkela_wire_3085),
        .dout(new_Jinkela_wire_3086)
    );

    bfr new_Jinkela_buffer_2789 (
        .din(new_Jinkela_wire_3203),
        .dout(new_Jinkela_wire_3204)
    );

    bfr new_Jinkela_buffer_2677 (
        .din(new_Jinkela_wire_3086),
        .dout(new_Jinkela_wire_3087)
    );

    bfr new_Jinkela_buffer_2725 (
        .din(new_Jinkela_wire_3139),
        .dout(new_Jinkela_wire_3140)
    );

    bfr new_Jinkela_buffer_2678 (
        .din(new_Jinkela_wire_3087),
        .dout(new_Jinkela_wire_3088)
    );

    bfr new_Jinkela_buffer_2788 (
        .din(new_Jinkela_wire_3202),
        .dout(new_Jinkela_wire_3203)
    );

    bfr new_Jinkela_buffer_2679 (
        .din(new_Jinkela_wire_3088),
        .dout(new_Jinkela_wire_3089)
    );

    bfr new_Jinkela_buffer_2726 (
        .din(new_Jinkela_wire_3140),
        .dout(new_Jinkela_wire_3141)
    );

    bfr new_Jinkela_buffer_2680 (
        .din(new_Jinkela_wire_3089),
        .dout(new_Jinkela_wire_3090)
    );

    spl2 new_Jinkela_splitter_140 (
        .a(new_Jinkela_wire_3204),
        .b(new_Jinkela_wire_3205),
        .c(new_Jinkela_wire_3206)
    );

    bfr new_Jinkela_buffer_2681 (
        .din(new_Jinkela_wire_3090),
        .dout(new_Jinkela_wire_3091)
    );

    bfr new_Jinkela_buffer_2727 (
        .din(new_Jinkela_wire_3141),
        .dout(new_Jinkela_wire_3142)
    );

    bfr new_Jinkela_buffer_2682 (
        .din(new_Jinkela_wire_3091),
        .dout(new_Jinkela_wire_3092)
    );

    bfr new_Jinkela_buffer_2790 (
        .din(new_Jinkela_wire_3206),
        .dout(new_Jinkela_wire_3207)
    );

    bfr new_Jinkela_buffer_2683 (
        .din(new_Jinkela_wire_3092),
        .dout(new_Jinkela_wire_3093)
    );

    bfr new_Jinkela_buffer_2728 (
        .din(new_Jinkela_wire_3142),
        .dout(new_Jinkela_wire_3143)
    );

    bfr new_Jinkela_buffer_2684 (
        .din(new_Jinkela_wire_3093),
        .dout(new_Jinkela_wire_3094)
    );

    bfr new_Jinkela_buffer_2916 (
        .din(new_Jinkela_wire_3339),
        .dout(new_Jinkela_wire_3340)
    );

    bfr new_Jinkela_buffer_2685 (
        .din(new_Jinkela_wire_3094),
        .dout(new_Jinkela_wire_3095)
    );

    bfr new_Jinkela_buffer_2729 (
        .din(new_Jinkela_wire_3143),
        .dout(new_Jinkela_wire_3144)
    );

    bfr new_Jinkela_buffer_2686 (
        .din(new_Jinkela_wire_3095),
        .dout(new_Jinkela_wire_3096)
    );

    bfr new_Jinkela_buffer_2919 (
        .din(N194),
        .dout(new_Jinkela_wire_3343)
    );

    bfr new_Jinkela_buffer_2687 (
        .din(new_Jinkela_wire_3096),
        .dout(new_Jinkela_wire_3097)
    );

    bfr new_Jinkela_buffer_4401 (
        .din(new_Jinkela_wire_5237),
        .dout(new_Jinkela_wire_5238)
    );

    bfr new_Jinkela_buffer_3584 (
        .din(n_0172_),
        .dout(new_Jinkela_wire_4189)
    );

    bfr new_Jinkela_buffer_3518 (
        .din(new_Jinkela_wire_4113),
        .dout(new_Jinkela_wire_4114)
    );

    bfr new_Jinkela_buffer_4382 (
        .din(new_Jinkela_wire_5201),
        .dout(new_Jinkela_wire_5202)
    );

    bfr new_Jinkela_buffer_7963 (
        .din(new_Jinkela_wire_10035),
        .dout(new_Jinkela_wire_10036)
    );

    bfr new_Jinkela_buffer_7909 (
        .din(new_Jinkela_wire_9976),
        .dout(new_Jinkela_wire_9977)
    );

    bfr new_Jinkela_buffer_4361 (
        .din(new_Jinkela_wire_5178),
        .dout(new_Jinkela_wire_5179)
    );

    spl3L new_Jinkela_splitter_221 (
        .a(n_0110_),
        .d(new_Jinkela_wire_4238),
        .b(new_Jinkela_wire_4239),
        .c(new_Jinkela_wire_4240)
    );

    bfr new_Jinkela_buffer_7922 (
        .din(new_Jinkela_wire_9991),
        .dout(new_Jinkela_wire_9992)
    );

    bfr new_Jinkela_buffer_3535 (
        .din(new_Jinkela_wire_4132),
        .dout(new_Jinkela_wire_4133)
    );

    bfr new_Jinkela_buffer_3519 (
        .din(new_Jinkela_wire_4114),
        .dout(new_Jinkela_wire_4115)
    );

    bfr new_Jinkela_buffer_4400 (
        .din(n_0341_),
        .dout(new_Jinkela_wire_5237)
    );

    bfr new_Jinkela_buffer_7910 (
        .din(new_Jinkela_wire_9977),
        .dout(new_Jinkela_wire_9978)
    );

    bfr new_Jinkela_buffer_4362 (
        .din(new_Jinkela_wire_5179),
        .dout(new_Jinkela_wire_5180)
    );

    bfr new_Jinkela_buffer_3520 (
        .din(new_Jinkela_wire_4115),
        .dout(new_Jinkela_wire_4116)
    );

    bfr new_Jinkela_buffer_4412 (
        .din(n_0822_),
        .dout(new_Jinkela_wire_5249)
    );

    bfr new_Jinkela_buffer_7911 (
        .din(new_Jinkela_wire_9978),
        .dout(new_Jinkela_wire_9979)
    );

    bfr new_Jinkela_buffer_4363 (
        .din(new_Jinkela_wire_5180),
        .dout(new_Jinkela_wire_5181)
    );

    bfr new_Jinkela_buffer_3581 (
        .din(new_Jinkela_wire_4183),
        .dout(new_Jinkela_wire_4184)
    );

    bfr new_Jinkela_buffer_7923 (
        .din(new_Jinkela_wire_9992),
        .dout(new_Jinkela_wire_9993)
    );

    bfr new_Jinkela_buffer_3536 (
        .din(new_Jinkela_wire_4133),
        .dout(new_Jinkela_wire_4134)
    );

    bfr new_Jinkela_buffer_3521 (
        .din(new_Jinkela_wire_4116),
        .dout(new_Jinkela_wire_4117)
    );

    bfr new_Jinkela_buffer_4383 (
        .din(new_Jinkela_wire_5202),
        .dout(new_Jinkela_wire_5203)
    );

    bfr new_Jinkela_buffer_7912 (
        .din(new_Jinkela_wire_9979),
        .dout(new_Jinkela_wire_9980)
    );

    bfr new_Jinkela_buffer_4364 (
        .din(new_Jinkela_wire_5181),
        .dout(new_Jinkela_wire_5182)
    );

    bfr new_Jinkela_buffer_3522 (
        .din(new_Jinkela_wire_4117),
        .dout(new_Jinkela_wire_4118)
    );

    spl2 new_Jinkela_splitter_308 (
        .a(new_Jinkela_wire_5203),
        .b(new_Jinkela_wire_5204),
        .c(new_Jinkela_wire_5205)
    );

    bfr new_Jinkela_buffer_7964 (
        .din(new_Jinkela_wire_10036),
        .dout(new_Jinkela_wire_10037)
    );

    bfr new_Jinkela_buffer_7913 (
        .din(new_Jinkela_wire_9980),
        .dout(new_Jinkela_wire_9981)
    );

    bfr new_Jinkela_buffer_4365 (
        .din(new_Jinkela_wire_5182),
        .dout(new_Jinkela_wire_5183)
    );

    bfr new_Jinkela_buffer_7924 (
        .din(new_Jinkela_wire_9993),
        .dout(new_Jinkela_wire_9994)
    );

    bfr new_Jinkela_buffer_4384 (
        .din(new_Jinkela_wire_5205),
        .dout(new_Jinkela_wire_5206)
    );

    bfr new_Jinkela_buffer_3537 (
        .din(new_Jinkela_wire_4134),
        .dout(new_Jinkela_wire_4135)
    );

    spl2 new_Jinkela_splitter_214 (
        .a(new_Jinkela_wire_4118),
        .b(new_Jinkela_wire_4119),
        .c(new_Jinkela_wire_4120)
    );

    bfr new_Jinkela_buffer_7914 (
        .din(new_Jinkela_wire_9981),
        .dout(new_Jinkela_wire_9982)
    );

    bfr new_Jinkela_buffer_4366 (
        .din(new_Jinkela_wire_5183),
        .dout(new_Jinkela_wire_5184)
    );

    bfr new_Jinkela_buffer_3582 (
        .din(new_Jinkela_wire_4184),
        .dout(new_Jinkela_wire_4185)
    );

    bfr new_Jinkela_buffer_3538 (
        .din(new_Jinkela_wire_4135),
        .dout(new_Jinkela_wire_4136)
    );

    spl2 new_Jinkela_splitter_834 (
        .a(n_0036_),
        .b(new_Jinkela_wire_10104),
        .c(new_Jinkela_wire_10105)
    );

    bfr new_Jinkela_buffer_7925 (
        .din(new_Jinkela_wire_9994),
        .dout(new_Jinkela_wire_9995)
    );

    bfr new_Jinkela_buffer_4367 (
        .din(new_Jinkela_wire_5184),
        .dout(new_Jinkela_wire_5185)
    );

    spl3L new_Jinkela_splitter_219 (
        .a(n_1054_),
        .d(new_Jinkela_wire_4233),
        .b(new_Jinkela_wire_4234),
        .c(new_Jinkela_wire_4235)
    );

    spl3L new_Jinkela_splitter_315 (
        .a(n_0161_),
        .d(new_Jinkela_wire_5250),
        .b(new_Jinkela_wire_5251),
        .c(new_Jinkela_wire_5252)
    );

    bfr new_Jinkela_buffer_3585 (
        .din(new_Jinkela_wire_4189),
        .dout(new_Jinkela_wire_4190)
    );

    bfr new_Jinkela_buffer_4413 (
        .din(new_net_2503),
        .dout(new_Jinkela_wire_5253)
    );

    bfr new_Jinkela_buffer_7965 (
        .din(new_Jinkela_wire_10037),
        .dout(new_Jinkela_wire_10038)
    );

    bfr new_Jinkela_buffer_7926 (
        .din(new_Jinkela_wire_9995),
        .dout(new_Jinkela_wire_9996)
    );

    bfr new_Jinkela_buffer_4368 (
        .din(new_Jinkela_wire_5185),
        .dout(new_Jinkela_wire_5186)
    );

    bfr new_Jinkela_buffer_3539 (
        .din(new_Jinkela_wire_4136),
        .dout(new_Jinkela_wire_4137)
    );

    bfr new_Jinkela_buffer_4402 (
        .din(new_Jinkela_wire_5238),
        .dout(new_Jinkela_wire_5239)
    );

    bfr new_Jinkela_buffer_3583 (
        .din(new_Jinkela_wire_4185),
        .dout(new_Jinkela_wire_4186)
    );

    bfr new_Jinkela_buffer_4385 (
        .din(new_Jinkela_wire_5206),
        .dout(new_Jinkela_wire_5207)
    );

    spl2 new_Jinkela_splitter_835 (
        .a(n_0267_),
        .b(new_Jinkela_wire_10135),
        .c(new_Jinkela_wire_10136)
    );

    bfr new_Jinkela_buffer_7927 (
        .din(new_Jinkela_wire_9996),
        .dout(new_Jinkela_wire_9997)
    );

    bfr new_Jinkela_buffer_4369 (
        .din(new_Jinkela_wire_5186),
        .dout(new_Jinkela_wire_5187)
    );

    bfr new_Jinkela_buffer_3540 (
        .din(new_Jinkela_wire_4137),
        .dout(new_Jinkela_wire_4138)
    );

    bfr new_Jinkela_buffer_8025 (
        .din(new_Jinkela_wire_10105),
        .dout(new_Jinkela_wire_10106)
    );

    spl2 new_Jinkela_splitter_220 (
        .a(new_Jinkela_wire_4235),
        .b(new_Jinkela_wire_4236),
        .c(new_Jinkela_wire_4237)
    );

    bfr new_Jinkela_buffer_7966 (
        .din(new_Jinkela_wire_10038),
        .dout(new_Jinkela_wire_10039)
    );

    bfr new_Jinkela_buffer_7928 (
        .din(new_Jinkela_wire_9997),
        .dout(new_Jinkela_wire_9998)
    );

    bfr new_Jinkela_buffer_4370 (
        .din(new_Jinkela_wire_5187),
        .dout(new_Jinkela_wire_5188)
    );

    bfr new_Jinkela_buffer_3541 (
        .din(new_Jinkela_wire_4138),
        .dout(new_Jinkela_wire_4139)
    );

    bfr new_Jinkela_buffer_3586 (
        .din(new_Jinkela_wire_4190),
        .dout(new_Jinkela_wire_4191)
    );

    bfr new_Jinkela_buffer_4386 (
        .din(new_Jinkela_wire_5207),
        .dout(new_Jinkela_wire_5208)
    );

    spl4L new_Jinkela_splitter_836 (
        .a(n_0848_),
        .d(new_Jinkela_wire_10137),
        .b(new_Jinkela_wire_10138),
        .e(new_Jinkela_wire_10139),
        .c(new_Jinkela_wire_10140)
    );

    bfr new_Jinkela_buffer_7929 (
        .din(new_Jinkela_wire_9998),
        .dout(new_Jinkela_wire_9999)
    );

    bfr new_Jinkela_buffer_4371 (
        .din(new_Jinkela_wire_5188),
        .dout(new_Jinkela_wire_5189)
    );

    bfr new_Jinkela_buffer_3542 (
        .din(new_Jinkela_wire_4139),
        .dout(new_Jinkela_wire_4140)
    );

    spl2 new_Jinkela_splitter_839 (
        .a(n_0102_),
        .b(new_Jinkela_wire_10148),
        .c(new_Jinkela_wire_10149)
    );

    spl2 new_Jinkela_splitter_316 (
        .a(n_0128_),
        .b(new_Jinkela_wire_5278),
        .c(new_Jinkela_wire_5279)
    );

    bfr new_Jinkela_buffer_7967 (
        .din(new_Jinkela_wire_10039),
        .dout(new_Jinkela_wire_10040)
    );

    bfr new_Jinkela_buffer_7930 (
        .din(new_Jinkela_wire_9999),
        .dout(new_Jinkela_wire_10000)
    );

    bfr new_Jinkela_buffer_4372 (
        .din(new_Jinkela_wire_5189),
        .dout(new_Jinkela_wire_5190)
    );

    bfr new_Jinkela_buffer_3543 (
        .din(new_Jinkela_wire_4140),
        .dout(new_Jinkela_wire_4141)
    );

    bfr new_Jinkela_buffer_4403 (
        .din(new_Jinkela_wire_5239),
        .dout(new_Jinkela_wire_5240)
    );

    bfr new_Jinkela_buffer_3627 (
        .din(new_Jinkela_wire_4241),
        .dout(new_Jinkela_wire_4242)
    );

    bfr new_Jinkela_buffer_3587 (
        .din(new_Jinkela_wire_4191),
        .dout(new_Jinkela_wire_4192)
    );

    bfr new_Jinkela_buffer_4387 (
        .din(new_Jinkela_wire_5208),
        .dout(new_Jinkela_wire_5209)
    );

    bfr new_Jinkela_buffer_8054 (
        .din(n_0506_),
        .dout(new_Jinkela_wire_10141)
    );

    bfr new_Jinkela_buffer_7931 (
        .din(new_Jinkela_wire_10000),
        .dout(new_Jinkela_wire_10001)
    );

    bfr new_Jinkela_buffer_4373 (
        .din(new_Jinkela_wire_5190),
        .dout(new_Jinkela_wire_5191)
    );

    bfr new_Jinkela_buffer_3544 (
        .din(new_Jinkela_wire_4141),
        .dout(new_Jinkela_wire_4142)
    );

    bfr new_Jinkela_buffer_8026 (
        .din(new_Jinkela_wire_10106),
        .dout(new_Jinkela_wire_10107)
    );

    bfr new_Jinkela_buffer_7968 (
        .din(new_Jinkela_wire_10040),
        .dout(new_Jinkela_wire_10041)
    );

    bfr new_Jinkela_buffer_7932 (
        .din(new_Jinkela_wire_10001),
        .dout(new_Jinkela_wire_10002)
    );

    bfr new_Jinkela_buffer_4374 (
        .din(new_Jinkela_wire_5191),
        .dout(new_Jinkela_wire_5192)
    );

    bfr new_Jinkela_buffer_3545 (
        .din(new_Jinkela_wire_4142),
        .dout(new_Jinkela_wire_4143)
    );

    bfr new_Jinkela_buffer_4438 (
        .din(n_0617_),
        .dout(new_Jinkela_wire_5280)
    );

    bfr new_Jinkela_buffer_3662 (
        .din(new_net_2556),
        .dout(new_Jinkela_wire_4277)
    );

    spl2 new_Jinkela_splitter_218 (
        .a(new_Jinkela_wire_4192),
        .b(new_Jinkela_wire_4193),
        .c(new_Jinkela_wire_4194)
    );

    bfr new_Jinkela_buffer_4388 (
        .din(new_Jinkela_wire_5209),
        .dout(new_Jinkela_wire_5210)
    );

    bfr new_Jinkela_buffer_7933 (
        .din(new_Jinkela_wire_10002),
        .dout(new_Jinkela_wire_10003)
    );

    bfr new_Jinkela_buffer_4375 (
        .din(new_Jinkela_wire_5192),
        .dout(new_Jinkela_wire_5193)
    );

    bfr new_Jinkela_buffer_3546 (
        .din(new_Jinkela_wire_4143),
        .dout(new_Jinkela_wire_4144)
    );

    spl2 new_Jinkela_splitter_838 (
        .a(n_1323_),
        .b(new_Jinkela_wire_10146),
        .c(new_Jinkela_wire_10147)
    );

    bfr new_Jinkela_buffer_3588 (
        .din(new_Jinkela_wire_4194),
        .dout(new_Jinkela_wire_4195)
    );

    bfr new_Jinkela_buffer_7969 (
        .din(new_Jinkela_wire_10041),
        .dout(new_Jinkela_wire_10042)
    );

    bfr new_Jinkela_buffer_7934 (
        .din(new_Jinkela_wire_10003),
        .dout(new_Jinkela_wire_10004)
    );

    bfr new_Jinkela_buffer_4376 (
        .din(new_Jinkela_wire_5193),
        .dout(new_Jinkela_wire_5194)
    );

    bfr new_Jinkela_buffer_3547 (
        .din(new_Jinkela_wire_4144),
        .dout(new_Jinkela_wire_4145)
    );

    bfr new_Jinkela_buffer_4404 (
        .din(new_Jinkela_wire_5240),
        .dout(new_Jinkela_wire_5241)
    );

    bfr new_Jinkela_buffer_4389 (
        .din(new_Jinkela_wire_5210),
        .dout(new_Jinkela_wire_5211)
    );

    bfr new_Jinkela_buffer_7935 (
        .din(new_Jinkela_wire_10004),
        .dout(new_Jinkela_wire_10005)
    );

    spl2 new_Jinkela_splitter_307 (
        .a(new_Jinkela_wire_5194),
        .b(new_Jinkela_wire_5195),
        .c(new_Jinkela_wire_5196)
    );

    bfr new_Jinkela_buffer_3548 (
        .din(new_Jinkela_wire_4145),
        .dout(new_Jinkela_wire_4146)
    );

    bfr new_Jinkela_buffer_8027 (
        .din(new_Jinkela_wire_10107),
        .dout(new_Jinkela_wire_10108)
    );

    bfr new_Jinkela_buffer_4414 (
        .din(new_Jinkela_wire_5253),
        .dout(new_Jinkela_wire_5254)
    );

    bfr new_Jinkela_buffer_3626 (
        .din(new_Jinkela_wire_4240),
        .dout(new_Jinkela_wire_4241)
    );

    bfr new_Jinkela_buffer_4390 (
        .din(new_Jinkela_wire_5211),
        .dout(new_Jinkela_wire_5212)
    );

    bfr new_Jinkela_buffer_7970 (
        .din(new_Jinkela_wire_10042),
        .dout(new_Jinkela_wire_10043)
    );

    bfr new_Jinkela_buffer_7936 (
        .din(new_Jinkela_wire_10005),
        .dout(new_Jinkela_wire_10006)
    );

    bfr new_Jinkela_buffer_3549 (
        .din(new_Jinkela_wire_4146),
        .dout(new_Jinkela_wire_4147)
    );

    bfr new_Jinkela_buffer_3663 (
        .din(new_Jinkela_wire_4277),
        .dout(new_Jinkela_wire_4278)
    );

    bfr new_Jinkela_buffer_3589 (
        .din(new_Jinkela_wire_4195),
        .dout(new_Jinkela_wire_4196)
    );

    bfr new_Jinkela_buffer_7937 (
        .din(new_Jinkela_wire_10006),
        .dout(new_Jinkela_wire_10007)
    );

    bfr new_Jinkela_buffer_4405 (
        .din(new_Jinkela_wire_5241),
        .dout(new_Jinkela_wire_5242)
    );

    bfr new_Jinkela_buffer_3550 (
        .din(new_Jinkela_wire_4147),
        .dout(new_Jinkela_wire_4148)
    );

    bfr new_Jinkela_buffer_4391 (
        .din(new_Jinkela_wire_5212),
        .dout(new_Jinkela_wire_5213)
    );

    bfr new_Jinkela_buffer_3667 (
        .din(new_net_2521),
        .dout(new_Jinkela_wire_4282)
    );

    bfr new_Jinkela_buffer_7971 (
        .din(new_Jinkela_wire_10043),
        .dout(new_Jinkela_wire_10044)
    );

    bfr new_Jinkela_buffer_7938 (
        .din(new_Jinkela_wire_10007),
        .dout(new_Jinkela_wire_10008)
    );

    bfr new_Jinkela_buffer_3551 (
        .din(new_Jinkela_wire_4148),
        .dout(new_Jinkela_wire_4149)
    );

    bfr new_Jinkela_buffer_4392 (
        .din(new_Jinkela_wire_5213),
        .dout(new_Jinkela_wire_5214)
    );

    bfr new_Jinkela_buffer_3590 (
        .din(new_Jinkela_wire_4196),
        .dout(new_Jinkela_wire_4197)
    );

    bfr new_Jinkela_buffer_7939 (
        .din(new_Jinkela_wire_10008),
        .dout(new_Jinkela_wire_10009)
    );

    bfr new_Jinkela_buffer_4406 (
        .din(new_Jinkela_wire_5242),
        .dout(new_Jinkela_wire_5243)
    );

    bfr new_Jinkela_buffer_3552 (
        .din(new_Jinkela_wire_4149),
        .dout(new_Jinkela_wire_4150)
    );

    bfr new_Jinkela_buffer_4393 (
        .din(new_Jinkela_wire_5214),
        .dout(new_Jinkela_wire_5215)
    );

    and_bi n_2790_ (
        .a(new_Jinkela_wire_8812),
        .b(new_Jinkela_wire_9586),
        .c(n_0646_)
    );

    bfr new_Jinkela_buffer_1973 (
        .din(new_Jinkela_wire_2337),
        .dout(new_Jinkela_wire_2338)
    );

    and_bb n_2073_ (
        .a(new_Jinkela_wire_4646),
        .b(new_Jinkela_wire_521),
        .c(n_1338_)
    );

    bfr new_Jinkela_buffer_1939 (
        .din(new_Jinkela_wire_2299),
        .dout(new_Jinkela_wire_2300)
    );

    and_bi n_2791_ (
        .a(n_0645_),
        .b(n_0646_),
        .c(n_0647_)
    );

    or_bb n_2074_ (
        .a(new_Jinkela_wire_6154),
        .b(new_Jinkela_wire_9556),
        .c(n_1339_)
    );

    and_ii n_2792_ (
        .a(new_Jinkela_wire_6355),
        .b(new_Jinkela_wire_9001),
        .c(n_0648_)
    );

    bfr new_Jinkela_buffer_2024 (
        .din(new_Jinkela_wire_2393),
        .dout(new_Jinkela_wire_2394)
    );

    and_ii n_2075_ (
        .a(new_Jinkela_wire_7315),
        .b(new_Jinkela_wire_3677),
        .c(n_1340_)
    );

    bfr new_Jinkela_buffer_1940 (
        .din(new_Jinkela_wire_2300),
        .dout(new_Jinkela_wire_2301)
    );

    and_bb n_2793_ (
        .a(new_Jinkela_wire_6354),
        .b(new_Jinkela_wire_9000),
        .c(n_0649_)
    );

    inv n_2076_ (
        .din(new_Jinkela_wire_691),
        .dout(n_1341_)
    );

    and_ii n_2794_ (
        .a(n_0649_),
        .b(n_0648_),
        .c(n_0650_)
    );

    bfr new_Jinkela_buffer_1974 (
        .din(new_Jinkela_wire_2338),
        .dout(new_Jinkela_wire_2339)
    );

    and_bi n_2077_ (
        .a(new_Jinkela_wire_3937),
        .b(new_Jinkela_wire_6901),
        .c(n_1342_)
    );

    bfr new_Jinkela_buffer_1941 (
        .din(new_Jinkela_wire_2301),
        .dout(new_Jinkela_wire_2302)
    );

    or_bb n_2795_ (
        .a(new_Jinkela_wire_4079),
        .b(new_Jinkela_wire_9835),
        .c(n_0651_)
    );

    and_bi n_2078_ (
        .a(new_Jinkela_wire_6900),
        .b(new_Jinkela_wire_3939),
        .c(n_1343_)
    );

    and_bb n_2796_ (
        .a(new_Jinkela_wire_4078),
        .b(new_Jinkela_wire_9834),
        .c(n_0652_)
    );

    bfr new_Jinkela_buffer_2088 (
        .din(new_Jinkela_wire_2457),
        .dout(new_Jinkela_wire_2458)
    );

    inv n_2079_ (
        .din(new_Jinkela_wire_2165),
        .dout(n_1344_)
    );

    bfr new_Jinkela_buffer_1942 (
        .din(new_Jinkela_wire_2302),
        .dout(new_Jinkela_wire_2303)
    );

    and_bi n_2797_ (
        .a(n_0651_),
        .b(n_0652_),
        .c(new_net_2541)
    );

    and_bi n_2080_ (
        .a(new_Jinkela_wire_9019),
        .b(new_Jinkela_wire_8085),
        .c(n_1345_)
    );

    and_bi n_2798_ (
        .a(new_Jinkela_wire_10625),
        .b(new_Jinkela_wire_4922),
        .c(new_net_2554)
    );

    bfr new_Jinkela_buffer_1975 (
        .din(new_Jinkela_wire_2339),
        .dout(new_Jinkela_wire_2340)
    );

    inv n_2081_ (
        .din(new_Jinkela_wire_7115),
        .dout(n_1346_)
    );

    bfr new_Jinkela_buffer_1943 (
        .din(new_Jinkela_wire_2303),
        .dout(new_Jinkela_wire_2304)
    );

    and_bi n_2799_ (
        .a(new_Jinkela_wire_8435),
        .b(new_Jinkela_wire_3675),
        .c(new_net_2533)
    );

    and_bi n_2082_ (
        .a(new_Jinkela_wire_8084),
        .b(new_Jinkela_wire_9018),
        .c(n_1347_)
    );

    and_bi n_2800_ (
        .a(new_Jinkela_wire_10628),
        .b(new_Jinkela_wire_4921),
        .c(new_net_2552)
    );

    bfr new_Jinkela_buffer_2025 (
        .din(new_Jinkela_wire_2394),
        .dout(new_Jinkela_wire_2395)
    );

    and_bb n_2083_ (
        .a(new_Jinkela_wire_6840),
        .b(new_Jinkela_wire_1480),
        .c(n_1348_)
    );

    bfr new_Jinkela_buffer_1944 (
        .din(new_Jinkela_wire_2304),
        .dout(new_Jinkela_wire_2305)
    );

    and_bi n_2801_ (
        .a(new_Jinkela_wire_10626),
        .b(new_Jinkela_wire_4924),
        .c(new_net_2519)
    );

    or_bb n_2084_ (
        .a(new_Jinkela_wire_6842),
        .b(new_Jinkela_wire_1481),
        .c(n_1349_)
    );

    bfr new_Jinkela_buffer_1976 (
        .din(new_Jinkela_wire_2340),
        .dout(new_Jinkela_wire_2341)
    );

    inv n_2085_ (
        .din(new_Jinkela_wire_3049),
        .dout(n_1350_)
    );

    bfr new_Jinkela_buffer_2097 (
        .din(N178),
        .dout(new_Jinkela_wire_2467)
    );

    and_bi n_2086_ (
        .a(new_Jinkela_wire_4983),
        .b(new_Jinkela_wire_9249),
        .c(n_1351_)
    );

    bfr new_Jinkela_buffer_1977 (
        .din(new_Jinkela_wire_2341),
        .dout(new_Jinkela_wire_2342)
    );

    and_bi n_2087_ (
        .a(new_Jinkela_wire_8846),
        .b(new_Jinkela_wire_6408),
        .c(n_1352_)
    );

    or_bb n_1420_ (
        .a(new_Jinkela_wire_7749),
        .b(new_Jinkela_wire_4510),
        .c(n_0692_)
    );

    bfr new_Jinkela_buffer_2026 (
        .din(new_Jinkela_wire_2395),
        .dout(new_Jinkela_wire_2396)
    );

    and_ii n_2088_ (
        .a(n_1352_),
        .b(new_Jinkela_wire_5091),
        .c(n_1353_)
    );

    bfr new_Jinkela_buffer_1978 (
        .din(new_Jinkela_wire_2342),
        .dout(new_Jinkela_wire_2343)
    );

    and_ii n_2089_ (
        .a(new_Jinkela_wire_8515),
        .b(new_Jinkela_wire_8662),
        .c(n_1354_)
    );

    bfr new_Jinkela_buffer_2091 (
        .din(new_Jinkela_wire_2460),
        .dout(new_Jinkela_wire_2461)
    );

    and_bi n_2090_ (
        .a(new_Jinkela_wire_3790),
        .b(n_1354_),
        .c(n_1355_)
    );

    bfr new_Jinkela_buffer_1979 (
        .din(new_Jinkela_wire_2343),
        .dout(new_Jinkela_wire_2344)
    );

    and_ii n_2091_ (
        .a(new_Jinkela_wire_6139),
        .b(new_Jinkela_wire_4642),
        .c(n_1356_)
    );

    bfr new_Jinkela_buffer_2027 (
        .din(new_Jinkela_wire_2396),
        .dout(new_Jinkela_wire_2397)
    );

    or_bb n_2092_ (
        .a(n_1356_),
        .b(new_Jinkela_wire_7382),
        .c(n_1357_)
    );

    bfr new_Jinkela_buffer_1980 (
        .din(new_Jinkela_wire_2344),
        .dout(new_Jinkela_wire_2345)
    );

    inv n_2093_ (
        .din(new_Jinkela_wire_9250),
        .dout(n_1358_)
    );

    bfr new_Jinkela_buffer_2094 (
        .din(new_Jinkela_wire_2463),
        .dout(new_Jinkela_wire_2464)
    );

    or_bi n_2094_ (
        .a(new_Jinkela_wire_7323),
        .b(new_Jinkela_wire_9741),
        .c(n_1359_)
    );

    bfr new_Jinkela_buffer_1981 (
        .din(new_Jinkela_wire_2345),
        .dout(new_Jinkela_wire_2346)
    );

    and_bi n_2095_ (
        .a(new_Jinkela_wire_9033),
        .b(new_Jinkela_wire_10565),
        .c(n_1360_)
    );

    bfr new_Jinkela_buffer_2028 (
        .din(new_Jinkela_wire_2397),
        .dout(new_Jinkela_wire_2398)
    );

    or_bb n_2096_ (
        .a(n_1360_),
        .b(new_Jinkela_wire_6779),
        .c(n_1361_)
    );

    bfr new_Jinkela_buffer_1982 (
        .din(new_Jinkela_wire_2346),
        .dout(new_Jinkela_wire_2347)
    );

    and_bi n_2097_ (
        .a(new_Jinkela_wire_5218),
        .b(new_Jinkela_wire_5070),
        .c(n_1362_)
    );

    bfr new_Jinkela_buffer_2092 (
        .din(new_Jinkela_wire_2461),
        .dout(new_Jinkela_wire_2462)
    );

    and_bi n_2098_ (
        .a(new_Jinkela_wire_7993),
        .b(new_Jinkela_wire_9591),
        .c(n_1363_)
    );

    bfr new_Jinkela_buffer_1983 (
        .din(new_Jinkela_wire_2347),
        .dout(new_Jinkela_wire_2348)
    );

    and_bi n_2099_ (
        .a(new_Jinkela_wire_10564),
        .b(new_Jinkela_wire_7022),
        .c(n_1364_)
    );

    bfr new_Jinkela_buffer_2029 (
        .din(new_Jinkela_wire_2398),
        .dout(new_Jinkela_wire_2399)
    );

    and_bi n_2100_ (
        .a(new_Jinkela_wire_9036),
        .b(new_Jinkela_wire_8183),
        .c(n_1365_)
    );

    bfr new_Jinkela_buffer_1984 (
        .din(new_Jinkela_wire_2348),
        .dout(new_Jinkela_wire_2349)
    );

    or_bb n_2101_ (
        .a(n_1365_),
        .b(new_Jinkela_wire_6782),
        .c(n_1366_)
    );

    bfr new_Jinkela_buffer_2101 (
        .din(N191),
        .dout(new_Jinkela_wire_2471)
    );

    and_bi n_2102_ (
        .a(new_Jinkela_wire_4918),
        .b(new_Jinkela_wire_4782),
        .c(n_1367_)
    );

    bfr new_Jinkela_buffer_1985 (
        .din(new_Jinkela_wire_2349),
        .dout(new_Jinkela_wire_2350)
    );

    and_bi n_2103_ (
        .a(new_Jinkela_wire_8843),
        .b(new_Jinkela_wire_5087),
        .c(n_1368_)
    );

    bfr new_Jinkela_buffer_2030 (
        .din(new_Jinkela_wire_2399),
        .dout(new_Jinkela_wire_2400)
    );

    and_bi n_2104_ (
        .a(new_Jinkela_wire_9246),
        .b(new_Jinkela_wire_4982),
        .c(n_1369_)
    );

    bfr new_Jinkela_buffer_1986 (
        .din(new_Jinkela_wire_2350),
        .dout(new_Jinkela_wire_2351)
    );

    and_ii n_2105_ (
        .a(new_Jinkela_wire_9347),
        .b(new_Jinkela_wire_6404),
        .c(n_1370_)
    );

    bfr new_Jinkela_buffer_2095 (
        .din(new_Jinkela_wire_2464),
        .dout(new_Jinkela_wire_2465)
    );

    or_ii n_2106_ (
        .a(new_Jinkela_wire_9118),
        .b(new_Jinkela_wire_10504),
        .c(n_1371_)
    );

    bfr new_Jinkela_buffer_1987 (
        .din(new_Jinkela_wire_2351),
        .dout(new_Jinkela_wire_2352)
    );

    and_ii n_2107_ (
        .a(new_Jinkela_wire_8657),
        .b(new_Jinkela_wire_7114),
        .c(n_0000_)
    );

    bfr new_Jinkela_buffer_2031 (
        .din(new_Jinkela_wire_2400),
        .dout(new_Jinkela_wire_2401)
    );

    and_ii n_2108_ (
        .a(new_Jinkela_wire_4633),
        .b(new_Jinkela_wire_7372),
        .c(n_0001_)
    );

    bfr new_Jinkela_buffer_1988 (
        .din(new_Jinkela_wire_2352),
        .dout(new_Jinkela_wire_2353)
    );

    or_ii n_2109_ (
        .a(new_Jinkela_wire_6746),
        .b(new_Jinkela_wire_5881),
        .c(n_0002_)
    );

    bfr new_Jinkela_buffer_2098 (
        .din(new_Jinkela_wire_2467),
        .dout(new_Jinkela_wire_2468)
    );

    or_bb n_2110_ (
        .a(new_Jinkela_wire_4525),
        .b(new_Jinkela_wire_3730),
        .c(n_0003_)
    );

    bfr new_Jinkela_buffer_1989 (
        .din(new_Jinkela_wire_2353),
        .dout(new_Jinkela_wire_2354)
    );

    and_bi n_2111_ (
        .a(new_Jinkela_wire_9709),
        .b(new_Jinkela_wire_4306),
        .c(n_0004_)
    );

    bfr new_Jinkela_buffer_2032 (
        .din(new_Jinkela_wire_2401),
        .dout(new_Jinkela_wire_2402)
    );

    and_bi n_2112_ (
        .a(new_Jinkela_wire_6548),
        .b(n_0004_),
        .c(n_0005_)
    );

    bfr new_Jinkela_buffer_1990 (
        .din(new_Jinkela_wire_2354),
        .dout(new_Jinkela_wire_2355)
    );

    or_bi n_2113_ (
        .a(new_Jinkela_wire_9434),
        .b(new_Jinkela_wire_7819),
        .c(n_0006_)
    );

    bfr new_Jinkela_buffer_2096 (
        .din(new_Jinkela_wire_2465),
        .dout(new_Jinkela_wire_2466)
    );

    and_bi n_2114_ (
        .a(new_Jinkela_wire_9930),
        .b(new_Jinkela_wire_8761),
        .c(n_0007_)
    );

    bfr new_Jinkela_buffer_5240 (
        .din(new_Jinkela_wire_6274),
        .dout(new_Jinkela_wire_6275)
    );

    bfr new_Jinkela_buffer_485 (
        .din(new_Jinkela_wire_526),
        .dout(new_Jinkela_wire_527)
    );

    bfr new_Jinkela_buffer_5213 (
        .din(new_Jinkela_wire_6234),
        .dout(new_Jinkela_wire_6235)
    );

    bfr new_Jinkela_buffer_434 (
        .din(new_Jinkela_wire_470),
        .dout(new_Jinkela_wire_471)
    );

    spl2 new_Jinkela_splitter_18 (
        .a(N271),
        .b(new_Jinkela_wire_599),
        .c(new_Jinkela_wire_600)
    );

    bfr new_Jinkela_buffer_557 (
        .din(N88),
        .dout(new_Jinkela_wire_601)
    );

    bfr new_Jinkela_buffer_5214 (
        .din(new_Jinkela_wire_6235),
        .dout(new_Jinkela_wire_6236)
    );

    bfr new_Jinkela_buffer_435 (
        .din(new_Jinkela_wire_471),
        .dout(new_Jinkela_wire_472)
    );

    bfr new_Jinkela_buffer_5276 (
        .din(new_Jinkela_wire_6319),
        .dout(new_Jinkela_wire_6320)
    );

    bfr new_Jinkela_buffer_5241 (
        .din(new_Jinkela_wire_6275),
        .dout(new_Jinkela_wire_6276)
    );

    bfr new_Jinkela_buffer_486 (
        .din(new_Jinkela_wire_527),
        .dout(new_Jinkela_wire_528)
    );

    bfr new_Jinkela_buffer_5215 (
        .din(new_Jinkela_wire_6236),
        .dout(new_Jinkela_wire_6237)
    );

    bfr new_Jinkela_buffer_436 (
        .din(new_Jinkela_wire_472),
        .dout(new_Jinkela_wire_473)
    );

    bfr new_Jinkela_buffer_551 (
        .din(new_Jinkela_wire_592),
        .dout(new_Jinkela_wire_593)
    );

    bfr new_Jinkela_buffer_5278 (
        .din(n_0616_),
        .dout(new_Jinkela_wire_6324)
    );

    bfr new_Jinkela_buffer_5242 (
        .din(new_Jinkela_wire_6276),
        .dout(new_Jinkela_wire_6277)
    );

    bfr new_Jinkela_buffer_437 (
        .din(new_Jinkela_wire_473),
        .dout(new_Jinkela_wire_474)
    );

    spl2 new_Jinkela_splitter_405 (
        .a(n_0732_),
        .b(new_Jinkela_wire_6331),
        .c(new_Jinkela_wire_6332)
    );

    bfr new_Jinkela_buffer_487 (
        .din(new_Jinkela_wire_528),
        .dout(new_Jinkela_wire_529)
    );

    spl2 new_Jinkela_splitter_406 (
        .a(n_1117_),
        .b(new_Jinkela_wire_6333),
        .c(new_Jinkela_wire_6334)
    );

    bfr new_Jinkela_buffer_5243 (
        .din(new_Jinkela_wire_6277),
        .dout(new_Jinkela_wire_6278)
    );

    bfr new_Jinkela_buffer_438 (
        .din(new_Jinkela_wire_474),
        .dout(new_Jinkela_wire_475)
    );

    bfr new_Jinkela_buffer_554 (
        .din(new_Jinkela_wire_595),
        .dout(new_Jinkela_wire_596)
    );

    bfr new_Jinkela_buffer_5279 (
        .din(new_Jinkela_wire_6324),
        .dout(new_Jinkela_wire_6325)
    );

    bfr new_Jinkela_buffer_5244 (
        .din(new_Jinkela_wire_6278),
        .dout(new_Jinkela_wire_6279)
    );

    bfr new_Jinkela_buffer_439 (
        .din(new_Jinkela_wire_475),
        .dout(new_Jinkela_wire_476)
    );

    bfr new_Jinkela_buffer_488 (
        .din(new_Jinkela_wire_529),
        .dout(new_Jinkela_wire_530)
    );

    bfr new_Jinkela_buffer_5245 (
        .din(new_Jinkela_wire_6279),
        .dout(new_Jinkela_wire_6280)
    );

    bfr new_Jinkela_buffer_440 (
        .din(new_Jinkela_wire_476),
        .dout(new_Jinkela_wire_477)
    );

    bfr new_Jinkela_buffer_5280 (
        .din(new_Jinkela_wire_6325),
        .dout(new_Jinkela_wire_6326)
    );

    bfr new_Jinkela_buffer_552 (
        .din(new_Jinkela_wire_593),
        .dout(new_Jinkela_wire_594)
    );

    bfr new_Jinkela_buffer_5246 (
        .din(new_Jinkela_wire_6280),
        .dout(new_Jinkela_wire_6281)
    );

    bfr new_Jinkela_buffer_441 (
        .din(new_Jinkela_wire_477),
        .dout(new_Jinkela_wire_478)
    );

    bfr new_Jinkela_buffer_489 (
        .din(new_Jinkela_wire_530),
        .dout(new_Jinkela_wire_531)
    );

    bfr new_Jinkela_buffer_5247 (
        .din(new_Jinkela_wire_6281),
        .dout(new_Jinkela_wire_6282)
    );

    bfr new_Jinkela_buffer_442 (
        .din(new_Jinkela_wire_478),
        .dout(new_Jinkela_wire_479)
    );

    spl3L new_Jinkela_splitter_407 (
        .a(n_1033_),
        .d(new_Jinkela_wire_6335),
        .b(new_Jinkela_wire_6336),
        .c(new_Jinkela_wire_6337)
    );

    bfr new_Jinkela_buffer_558 (
        .din(new_Jinkela_wire_601),
        .dout(new_Jinkela_wire_602)
    );

    bfr new_Jinkela_buffer_5281 (
        .din(new_Jinkela_wire_6326),
        .dout(new_Jinkela_wire_6327)
    );

    bfr new_Jinkela_buffer_5248 (
        .din(new_Jinkela_wire_6282),
        .dout(new_Jinkela_wire_6283)
    );

    bfr new_Jinkela_buffer_443 (
        .din(new_Jinkela_wire_479),
        .dout(new_Jinkela_wire_480)
    );

    bfr new_Jinkela_buffer_490 (
        .din(new_Jinkela_wire_531),
        .dout(new_Jinkela_wire_532)
    );

    spl2 new_Jinkela_splitter_408 (
        .a(new_Jinkela_wire_6337),
        .b(new_Jinkela_wire_6338),
        .c(new_Jinkela_wire_6339)
    );

    bfr new_Jinkela_buffer_5249 (
        .din(new_Jinkela_wire_6283),
        .dout(new_Jinkela_wire_6284)
    );

    bfr new_Jinkela_buffer_444 (
        .din(new_Jinkela_wire_480),
        .dout(new_Jinkela_wire_481)
    );

    bfr new_Jinkela_buffer_5283 (
        .din(n_0647_),
        .dout(new_Jinkela_wire_6340)
    );

    bfr new_Jinkela_buffer_555 (
        .din(new_Jinkela_wire_596),
        .dout(new_Jinkela_wire_597)
    );

    bfr new_Jinkela_buffer_5282 (
        .din(new_Jinkela_wire_6327),
        .dout(new_Jinkela_wire_6328)
    );

    bfr new_Jinkela_buffer_5250 (
        .din(new_Jinkela_wire_6284),
        .dout(new_Jinkela_wire_6285)
    );

    bfr new_Jinkela_buffer_445 (
        .din(new_Jinkela_wire_481),
        .dout(new_Jinkela_wire_482)
    );

    bfr new_Jinkela_buffer_491 (
        .din(new_Jinkela_wire_532),
        .dout(new_Jinkela_wire_533)
    );

    bfr new_Jinkela_buffer_5251 (
        .din(new_Jinkela_wire_6285),
        .dout(new_Jinkela_wire_6286)
    );

    bfr new_Jinkela_buffer_446 (
        .din(new_Jinkela_wire_482),
        .dout(new_Jinkela_wire_483)
    );

    bfr new_Jinkela_buffer_5331 (
        .din(n_0791_),
        .dout(new_Jinkela_wire_6394)
    );

    spl2 new_Jinkela_splitter_404 (
        .a(new_Jinkela_wire_6328),
        .b(new_Jinkela_wire_6329),
        .c(new_Jinkela_wire_6330)
    );

    bfr new_Jinkela_buffer_5252 (
        .din(new_Jinkela_wire_6286),
        .dout(new_Jinkela_wire_6287)
    );

    bfr new_Jinkela_buffer_447 (
        .din(new_Jinkela_wire_483),
        .dout(new_Jinkela_wire_484)
    );

    bfr new_Jinkela_buffer_492 (
        .din(new_Jinkela_wire_533),
        .dout(new_Jinkela_wire_534)
    );

    bfr new_Jinkela_buffer_5253 (
        .din(new_Jinkela_wire_6287),
        .dout(new_Jinkela_wire_6288)
    );

    bfr new_Jinkela_buffer_448 (
        .din(new_Jinkela_wire_484),
        .dout(new_Jinkela_wire_485)
    );

    spl4L new_Jinkela_splitter_410 (
        .a(n_1187_),
        .d(new_Jinkela_wire_6390),
        .b(new_Jinkela_wire_6391),
        .e(new_Jinkela_wire_6392),
        .c(new_Jinkela_wire_6393)
    );

    bfr new_Jinkela_buffer_556 (
        .din(new_Jinkela_wire_597),
        .dout(new_Jinkela_wire_598)
    );

    bfr new_Jinkela_buffer_5254 (
        .din(new_Jinkela_wire_6288),
        .dout(new_Jinkela_wire_6289)
    );

    bfr new_Jinkela_buffer_449 (
        .din(new_Jinkela_wire_485),
        .dout(new_Jinkela_wire_486)
    );

    bfr new_Jinkela_buffer_5297 (
        .din(new_net_2501),
        .dout(new_Jinkela_wire_6356)
    );

    bfr new_Jinkela_buffer_493 (
        .din(new_Jinkela_wire_534),
        .dout(new_Jinkela_wire_535)
    );

    bfr new_Jinkela_buffer_5284 (
        .din(new_Jinkela_wire_6340),
        .dout(new_Jinkela_wire_6341)
    );

    bfr new_Jinkela_buffer_5255 (
        .din(new_Jinkela_wire_6289),
        .dout(new_Jinkela_wire_6290)
    );

    bfr new_Jinkela_buffer_450 (
        .din(new_Jinkela_wire_486),
        .dout(new_Jinkela_wire_487)
    );

    bfr new_Jinkela_buffer_5298 (
        .din(new_Jinkela_wire_6356),
        .dout(new_Jinkela_wire_6357)
    );

    bfr new_Jinkela_buffer_561 (
        .din(N86),
        .dout(new_Jinkela_wire_605)
    );

    bfr new_Jinkela_buffer_5285 (
        .din(new_Jinkela_wire_6341),
        .dout(new_Jinkela_wire_6342)
    );

    bfr new_Jinkela_buffer_5256 (
        .din(new_Jinkela_wire_6290),
        .dout(new_Jinkela_wire_6291)
    );

    bfr new_Jinkela_buffer_451 (
        .din(new_Jinkela_wire_487),
        .dout(new_Jinkela_wire_488)
    );

    bfr new_Jinkela_buffer_494 (
        .din(new_Jinkela_wire_535),
        .dout(new_Jinkela_wire_536)
    );

    bfr new_Jinkela_buffer_5257 (
        .din(new_Jinkela_wire_6291),
        .dout(new_Jinkela_wire_6292)
    );

    bfr new_Jinkela_buffer_452 (
        .din(new_Jinkela_wire_488),
        .dout(new_Jinkela_wire_489)
    );

    bfr new_Jinkela_buffer_565 (
        .din(N242),
        .dout(new_Jinkela_wire_609)
    );

    bfr new_Jinkela_buffer_5286 (
        .din(new_Jinkela_wire_6342),
        .dout(new_Jinkela_wire_6343)
    );

    bfr new_Jinkela_buffer_5258 (
        .din(new_Jinkela_wire_6292),
        .dout(new_Jinkela_wire_6293)
    );

    bfr new_Jinkela_buffer_453 (
        .din(new_Jinkela_wire_489),
        .dout(new_Jinkela_wire_490)
    );

    bfr new_Jinkela_buffer_495 (
        .din(new_Jinkela_wire_536),
        .dout(new_Jinkela_wire_537)
    );

    bfr new_Jinkela_buffer_5259 (
        .din(new_Jinkela_wire_6293),
        .dout(new_Jinkela_wire_6294)
    );

    bfr new_Jinkela_buffer_454 (
        .din(new_Jinkela_wire_490),
        .dout(new_Jinkela_wire_491)
    );

    bfr new_Jinkela_buffer_8028 (
        .din(new_Jinkela_wire_10108),
        .dout(new_Jinkela_wire_10109)
    );

    spl2 new_Jinkela_splitter_525 (
        .a(n_0439_),
        .b(new_Jinkela_wire_7406),
        .c(new_Jinkela_wire_7407)
    );

    bfr new_Jinkela_buffer_7972 (
        .din(new_Jinkela_wire_10044),
        .dout(new_Jinkela_wire_10045)
    );

    bfr new_Jinkela_buffer_7940 (
        .din(new_Jinkela_wire_10009),
        .dout(new_Jinkela_wire_10010)
    );

    bfr new_Jinkela_buffer_6057 (
        .din(new_Jinkela_wire_7390),
        .dout(new_Jinkela_wire_7391)
    );

    bfr new_Jinkela_buffer_6044 (
        .din(new_Jinkela_wire_7375),
        .dout(new_Jinkela_wire_7376)
    );

    bfr new_Jinkela_buffer_6070 (
        .din(n_0681_),
        .dout(new_Jinkela_wire_7408)
    );

    bfr new_Jinkela_buffer_7941 (
        .din(new_Jinkela_wire_10010),
        .dout(new_Jinkela_wire_10011)
    );

    bfr new_Jinkela_buffer_6045 (
        .din(new_Jinkela_wire_7376),
        .dout(new_Jinkela_wire_7377)
    );

    bfr new_Jinkela_buffer_6053 (
        .din(new_Jinkela_wire_7386),
        .dout(new_Jinkela_wire_7387)
    );

    bfr new_Jinkela_buffer_7973 (
        .din(new_Jinkela_wire_10045),
        .dout(new_Jinkela_wire_10046)
    );

    bfr new_Jinkela_buffer_7942 (
        .din(new_Jinkela_wire_10011),
        .dout(new_Jinkela_wire_10012)
    );

    bfr new_Jinkela_buffer_6046 (
        .din(new_Jinkela_wire_7377),
        .dout(new_Jinkela_wire_7378)
    );

    spl2 new_Jinkela_splitter_526 (
        .a(n_0520_),
        .b(new_Jinkela_wire_7412),
        .c(new_Jinkela_wire_7413)
    );

    bfr new_Jinkela_buffer_8055 (
        .din(new_Jinkela_wire_10141),
        .dout(new_Jinkela_wire_10142)
    );

    bfr new_Jinkela_buffer_7943 (
        .din(new_Jinkela_wire_10012),
        .dout(new_Jinkela_wire_10013)
    );

    bfr new_Jinkela_buffer_6047 (
        .din(new_Jinkela_wire_7378),
        .dout(new_Jinkela_wire_7379)
    );

    bfr new_Jinkela_buffer_8029 (
        .din(new_Jinkela_wire_10109),
        .dout(new_Jinkela_wire_10110)
    );

    bfr new_Jinkela_buffer_6054 (
        .din(new_Jinkela_wire_7387),
        .dout(new_Jinkela_wire_7388)
    );

    bfr new_Jinkela_buffer_7974 (
        .din(new_Jinkela_wire_10046),
        .dout(new_Jinkela_wire_10047)
    );

    bfr new_Jinkela_buffer_7944 (
        .din(new_Jinkela_wire_10013),
        .dout(new_Jinkela_wire_10014)
    );

    bfr new_Jinkela_buffer_6048 (
        .din(new_Jinkela_wire_7379),
        .dout(new_Jinkela_wire_7380)
    );

    bfr new_Jinkela_buffer_7945 (
        .din(new_Jinkela_wire_10014),
        .dout(new_Jinkela_wire_10015)
    );

    bfr new_Jinkela_buffer_6071 (
        .din(n_0042_),
        .dout(new_Jinkela_wire_7409)
    );

    bfr new_Jinkela_buffer_6049 (
        .din(new_Jinkela_wire_7380),
        .dout(new_Jinkela_wire_7381)
    );

    bfr new_Jinkela_buffer_6055 (
        .din(new_Jinkela_wire_7388),
        .dout(new_Jinkela_wire_7389)
    );

    bfr new_Jinkela_buffer_7975 (
        .din(new_Jinkela_wire_10047),
        .dout(new_Jinkela_wire_10048)
    );

    bfr new_Jinkela_buffer_7946 (
        .din(new_Jinkela_wire_10015),
        .dout(new_Jinkela_wire_10016)
    );

    bfr new_Jinkela_buffer_6050 (
        .din(new_Jinkela_wire_7381),
        .dout(new_Jinkela_wire_7382)
    );

    spl4L new_Jinkela_splitter_527 (
        .a(n_0062_),
        .d(new_Jinkela_wire_7414),
        .b(new_Jinkela_wire_7415),
        .e(new_Jinkela_wire_7416),
        .c(new_Jinkela_wire_7417)
    );

    bfr new_Jinkela_buffer_8057 (
        .din(new_Jinkela_wire_10149),
        .dout(new_Jinkela_wire_10150)
    );

    bfr new_Jinkela_buffer_7947 (
        .din(new_Jinkela_wire_10016),
        .dout(new_Jinkela_wire_10017)
    );

    bfr new_Jinkela_buffer_6072 (
        .din(new_Jinkela_wire_7409),
        .dout(new_Jinkela_wire_7410)
    );

    bfr new_Jinkela_buffer_6056 (
        .din(new_Jinkela_wire_7389),
        .dout(new_Jinkela_wire_7390)
    );

    bfr new_Jinkela_buffer_8030 (
        .din(new_Jinkela_wire_10110),
        .dout(new_Jinkela_wire_10111)
    );

    bfr new_Jinkela_buffer_7976 (
        .din(new_Jinkela_wire_10048),
        .dout(new_Jinkela_wire_10049)
    );

    bfr new_Jinkela_buffer_7948 (
        .din(new_Jinkela_wire_10017),
        .dout(new_Jinkela_wire_10018)
    );

    spl4L new_Jinkela_splitter_529 (
        .a(n_0679_),
        .d(new_Jinkela_wire_7449),
        .b(new_Jinkela_wire_7450),
        .e(new_Jinkela_wire_7451),
        .c(new_Jinkela_wire_7452)
    );

    bfr new_Jinkela_buffer_7949 (
        .din(new_Jinkela_wire_10018),
        .dout(new_Jinkela_wire_10019)
    );

    bfr new_Jinkela_buffer_6073 (
        .din(new_Jinkela_wire_7410),
        .dout(new_Jinkela_wire_7411)
    );

    bfr new_Jinkela_buffer_6058 (
        .din(new_Jinkela_wire_7391),
        .dout(new_Jinkela_wire_7392)
    );

    bfr new_Jinkela_buffer_8056 (
        .din(new_Jinkela_wire_10142),
        .dout(new_Jinkela_wire_10143)
    );

    bfr new_Jinkela_buffer_7977 (
        .din(new_Jinkela_wire_10049),
        .dout(new_Jinkela_wire_10050)
    );

    bfr new_Jinkela_buffer_7950 (
        .din(new_Jinkela_wire_10019),
        .dout(new_Jinkela_wire_10020)
    );

    bfr new_Jinkela_buffer_6059 (
        .din(new_Jinkela_wire_7392),
        .dout(new_Jinkela_wire_7393)
    );

    bfr new_Jinkela_buffer_7951 (
        .din(new_Jinkela_wire_10020),
        .dout(new_Jinkela_wire_10021)
    );

    spl2 new_Jinkela_splitter_528 (
        .a(n_0092_),
        .b(new_Jinkela_wire_7447),
        .c(new_Jinkela_wire_7448)
    );

    bfr new_Jinkela_buffer_6060 (
        .din(new_Jinkela_wire_7393),
        .dout(new_Jinkela_wire_7394)
    );

    bfr new_Jinkela_buffer_8031 (
        .din(new_Jinkela_wire_10111),
        .dout(new_Jinkela_wire_10112)
    );

    bfr new_Jinkela_buffer_6075 (
        .din(new_Jinkela_wire_7418),
        .dout(new_Jinkela_wire_7419)
    );

    bfr new_Jinkela_buffer_7978 (
        .din(new_Jinkela_wire_10050),
        .dout(new_Jinkela_wire_10051)
    );

    bfr new_Jinkela_buffer_7952 (
        .din(new_Jinkela_wire_10021),
        .dout(new_Jinkela_wire_10022)
    );

    bfr new_Jinkela_buffer_6061 (
        .din(new_Jinkela_wire_7394),
        .dout(new_Jinkela_wire_7395)
    );

    bfr new_Jinkela_buffer_6074 (
        .din(new_Jinkela_wire_7417),
        .dout(new_Jinkela_wire_7418)
    );

    bfr new_Jinkela_buffer_7953 (
        .din(new_Jinkela_wire_10022),
        .dout(new_Jinkela_wire_10023)
    );

    spl2 new_Jinkela_splitter_532 (
        .a(n_0836_),
        .b(new_Jinkela_wire_7457),
        .c(new_Jinkela_wire_7458)
    );

    bfr new_Jinkela_buffer_6062 (
        .din(new_Jinkela_wire_7395),
        .dout(new_Jinkela_wire_7396)
    );

    spl2 new_Jinkela_splitter_530 (
        .a(n_0065_),
        .b(new_Jinkela_wire_7453),
        .c(new_Jinkela_wire_7454)
    );

    bfr new_Jinkela_buffer_7979 (
        .din(new_Jinkela_wire_10051),
        .dout(new_Jinkela_wire_10052)
    );

    bfr new_Jinkela_buffer_7954 (
        .din(new_Jinkela_wire_10023),
        .dout(new_Jinkela_wire_10024)
    );

    bfr new_Jinkela_buffer_6063 (
        .din(new_Jinkela_wire_7396),
        .dout(new_Jinkela_wire_7397)
    );

    spl2 new_Jinkela_splitter_531 (
        .a(n_0085_),
        .b(new_Jinkela_wire_7455),
        .c(new_Jinkela_wire_7456)
    );

    spl2 new_Jinkela_splitter_840 (
        .a(new_net_3),
        .b(new_Jinkela_wire_10154),
        .c(new_Jinkela_wire_10155)
    );

    bfr new_Jinkela_buffer_7955 (
        .din(new_Jinkela_wire_10024),
        .dout(new_Jinkela_wire_10025)
    );

    bfr new_Jinkela_buffer_6064 (
        .din(new_Jinkela_wire_7397),
        .dout(new_Jinkela_wire_7398)
    );

    bfr new_Jinkela_buffer_8032 (
        .din(new_Jinkela_wire_10112),
        .dout(new_Jinkela_wire_10113)
    );

    bfr new_Jinkela_buffer_6076 (
        .din(new_Jinkela_wire_7419),
        .dout(new_Jinkela_wire_7420)
    );

    bfr new_Jinkela_buffer_7980 (
        .din(new_Jinkela_wire_10052),
        .dout(new_Jinkela_wire_10053)
    );

    bfr new_Jinkela_buffer_7956 (
        .din(new_Jinkela_wire_10025),
        .dout(new_Jinkela_wire_10026)
    );

    bfr new_Jinkela_buffer_6065 (
        .din(new_Jinkela_wire_7398),
        .dout(new_Jinkela_wire_7399)
    );

    bfr new_Jinkela_buffer_7957 (
        .din(new_Jinkela_wire_10026),
        .dout(new_Jinkela_wire_10027)
    );

    bfr new_Jinkela_buffer_6066 (
        .din(new_Jinkela_wire_7399),
        .dout(new_Jinkela_wire_7400)
    );

    spl2 new_Jinkela_splitter_837 (
        .a(new_Jinkela_wire_10143),
        .b(new_Jinkela_wire_10144),
        .c(new_Jinkela_wire_10145)
    );

    bfr new_Jinkela_buffer_6077 (
        .din(new_Jinkela_wire_7420),
        .dout(new_Jinkela_wire_7421)
    );

    bfr new_Jinkela_buffer_7981 (
        .din(new_Jinkela_wire_10053),
        .dout(new_Jinkela_wire_10054)
    );

    bfr new_Jinkela_buffer_7958 (
        .din(new_Jinkela_wire_10027),
        .dout(new_Jinkela_wire_10028)
    );

    bfr new_Jinkela_buffer_6067 (
        .din(new_Jinkela_wire_7400),
        .dout(new_Jinkela_wire_7401)
    );

    spl2 new_Jinkela_splitter_533 (
        .a(n_0999_),
        .b(new_Jinkela_wire_7459),
        .c(new_Jinkela_wire_7460)
    );

    bfr new_Jinkela_buffer_7959 (
        .din(new_Jinkela_wire_10028),
        .dout(new_Jinkela_wire_10029)
    );

    bfr new_Jinkela_buffer_6068 (
        .din(new_Jinkela_wire_7401),
        .dout(new_Jinkela_wire_7402)
    );

    bfr new_Jinkela_buffer_8033 (
        .din(new_Jinkela_wire_10113),
        .dout(new_Jinkela_wire_10114)
    );

    bfr new_Jinkela_buffer_6078 (
        .din(new_Jinkela_wire_7421),
        .dout(new_Jinkela_wire_7422)
    );

    bfr new_Jinkela_buffer_7982 (
        .din(new_Jinkela_wire_10054),
        .dout(new_Jinkela_wire_10055)
    );

    bfr new_Jinkela_buffer_6069 (
        .din(new_Jinkela_wire_7402),
        .dout(new_Jinkela_wire_7403)
    );

    bfr new_Jinkela_buffer_6873 (
        .din(new_Jinkela_wire_8496),
        .dout(new_Jinkela_wire_8497)
    );

    bfr new_Jinkela_buffer_4415 (
        .din(new_Jinkela_wire_5254),
        .dout(new_Jinkela_wire_5255)
    );

    bfr new_Jinkela_buffer_4394 (
        .din(new_Jinkela_wire_5215),
        .dout(new_Jinkela_wire_5216)
    );

    bfr new_Jinkela_buffer_6905 (
        .din(new_Jinkela_wire_8535),
        .dout(new_Jinkela_wire_8536)
    );

    bfr new_Jinkela_buffer_6874 (
        .din(new_Jinkela_wire_8497),
        .dout(new_Jinkela_wire_8498)
    );

    bfr new_Jinkela_buffer_4407 (
        .din(new_Jinkela_wire_5243),
        .dout(new_Jinkela_wire_5244)
    );

    spl3L new_Jinkela_splitter_309 (
        .a(new_Jinkela_wire_5216),
        .d(new_Jinkela_wire_5217),
        .b(new_Jinkela_wire_5218),
        .c(new_Jinkela_wire_5219)
    );

    bfr new_Jinkela_buffer_6891 (
        .din(new_Jinkela_wire_8521),
        .dout(new_Jinkela_wire_8522)
    );

    bfr new_Jinkela_buffer_6875 (
        .din(new_Jinkela_wire_8498),
        .dout(new_Jinkela_wire_8499)
    );

    spl3L new_Jinkela_splitter_317 (
        .a(n_1021_),
        .d(new_Jinkela_wire_5282),
        .b(new_Jinkela_wire_5283),
        .c(new_Jinkela_wire_5284)
    );

    bfr new_Jinkela_buffer_4395 (
        .din(new_Jinkela_wire_5219),
        .dout(new_Jinkela_wire_5220)
    );

    bfr new_Jinkela_buffer_4439 (
        .din(n_0308_),
        .dout(new_Jinkela_wire_5281)
    );

    bfr new_Jinkela_buffer_6876 (
        .din(new_Jinkela_wire_8499),
        .dout(new_Jinkela_wire_8500)
    );

    bfr new_Jinkela_buffer_4408 (
        .din(new_Jinkela_wire_5244),
        .dout(new_Jinkela_wire_5245)
    );

    bfr new_Jinkela_buffer_4396 (
        .din(new_Jinkela_wire_5220),
        .dout(new_Jinkela_wire_5221)
    );

    bfr new_Jinkela_buffer_6892 (
        .din(new_Jinkela_wire_8522),
        .dout(new_Jinkela_wire_8523)
    );

    bfr new_Jinkela_buffer_6877 (
        .din(new_Jinkela_wire_8500),
        .dout(new_Jinkela_wire_8501)
    );

    bfr new_Jinkela_buffer_4416 (
        .din(new_Jinkela_wire_5255),
        .dout(new_Jinkela_wire_5256)
    );

    spl2 new_Jinkela_splitter_310 (
        .a(new_Jinkela_wire_5221),
        .b(new_Jinkela_wire_5222),
        .c(new_Jinkela_wire_5223)
    );

    spl4L new_Jinkela_splitter_653 (
        .a(n_1282_),
        .d(new_Jinkela_wire_8574),
        .b(new_Jinkela_wire_8575),
        .e(new_Jinkela_wire_8576),
        .c(new_Jinkela_wire_8577)
    );

    bfr new_Jinkela_buffer_6906 (
        .din(new_Jinkela_wire_8536),
        .dout(new_Jinkela_wire_8537)
    );

    bfr new_Jinkela_buffer_4397 (
        .din(new_Jinkela_wire_5223),
        .dout(new_Jinkela_wire_5224)
    );

    bfr new_Jinkela_buffer_6878 (
        .din(new_Jinkela_wire_8501),
        .dout(new_Jinkela_wire_8502)
    );

    bfr new_Jinkela_buffer_6893 (
        .din(new_Jinkela_wire_8523),
        .dout(new_Jinkela_wire_8524)
    );

    bfr new_Jinkela_buffer_4409 (
        .din(new_Jinkela_wire_5245),
        .dout(new_Jinkela_wire_5246)
    );

    bfr new_Jinkela_buffer_6879 (
        .din(new_Jinkela_wire_8502),
        .dout(new_Jinkela_wire_8503)
    );

    bfr new_Jinkela_buffer_4440 (
        .din(n_1177_),
        .dout(new_Jinkela_wire_5287)
    );

    bfr new_Jinkela_buffer_6911 (
        .din(new_Jinkela_wire_8541),
        .dout(new_Jinkela_wire_8542)
    );

    bfr new_Jinkela_buffer_4410 (
        .din(new_Jinkela_wire_5246),
        .dout(new_Jinkela_wire_5247)
    );

    bfr new_Jinkela_buffer_6880 (
        .din(new_Jinkela_wire_8503),
        .dout(new_Jinkela_wire_8504)
    );

    bfr new_Jinkela_buffer_4417 (
        .din(new_Jinkela_wire_5256),
        .dout(new_Jinkela_wire_5257)
    );

    bfr new_Jinkela_buffer_6894 (
        .din(new_Jinkela_wire_8524),
        .dout(new_Jinkela_wire_8525)
    );

    bfr new_Jinkela_buffer_4411 (
        .din(new_Jinkela_wire_5247),
        .dout(new_Jinkela_wire_5248)
    );

    bfr new_Jinkela_buffer_6881 (
        .din(new_Jinkela_wire_8504),
        .dout(new_Jinkela_wire_8505)
    );

    spl4L new_Jinkela_splitter_320 (
        .a(n_0881_),
        .d(new_Jinkela_wire_5292),
        .b(new_Jinkela_wire_5293),
        .e(new_Jinkela_wire_5294),
        .c(new_Jinkela_wire_5295)
    );

    bfr new_Jinkela_buffer_6907 (
        .din(new_Jinkela_wire_8537),
        .dout(new_Jinkela_wire_8538)
    );

    bfr new_Jinkela_buffer_4418 (
        .din(new_Jinkela_wire_5257),
        .dout(new_Jinkela_wire_5258)
    );

    bfr new_Jinkela_buffer_6882 (
        .din(new_Jinkela_wire_8505),
        .dout(new_Jinkela_wire_8506)
    );

    bfr new_Jinkela_buffer_6895 (
        .din(new_Jinkela_wire_8525),
        .dout(new_Jinkela_wire_8526)
    );

    bfr new_Jinkela_buffer_4419 (
        .din(new_Jinkela_wire_5258),
        .dout(new_Jinkela_wire_5259)
    );

    bfr new_Jinkela_buffer_6883 (
        .din(new_Jinkela_wire_8506),
        .dout(new_Jinkela_wire_8507)
    );

    spl2 new_Jinkela_splitter_318 (
        .a(new_Jinkela_wire_5284),
        .b(new_Jinkela_wire_5285),
        .c(new_Jinkela_wire_5286)
    );

    spl2 new_Jinkela_splitter_319 (
        .a(n_0781_),
        .b(new_Jinkela_wire_5288),
        .c(new_Jinkela_wire_5289)
    );

    bfr new_Jinkela_buffer_6937 (
        .din(new_Jinkela_wire_8569),
        .dout(new_Jinkela_wire_8570)
    );

    bfr new_Jinkela_buffer_4420 (
        .din(new_Jinkela_wire_5259),
        .dout(new_Jinkela_wire_5260)
    );

    bfr new_Jinkela_buffer_6884 (
        .din(new_Jinkela_wire_8507),
        .dout(new_Jinkela_wire_8508)
    );

    bfr new_Jinkela_buffer_6896 (
        .din(new_Jinkela_wire_8526),
        .dout(new_Jinkela_wire_8527)
    );

    bfr new_Jinkela_buffer_4421 (
        .din(new_Jinkela_wire_5260),
        .dout(new_Jinkela_wire_5261)
    );

    bfr new_Jinkela_buffer_6908 (
        .din(new_Jinkela_wire_8538),
        .dout(new_Jinkela_wire_8539)
    );

    bfr new_Jinkela_buffer_4441 (
        .din(new_Jinkela_wire_5289),
        .dout(new_Jinkela_wire_5290)
    );

    bfr new_Jinkela_buffer_6897 (
        .din(new_Jinkela_wire_8527),
        .dout(new_Jinkela_wire_8528)
    );

    bfr new_Jinkela_buffer_4422 (
        .din(new_Jinkela_wire_5261),
        .dout(new_Jinkela_wire_5262)
    );

    bfr new_Jinkela_buffer_6912 (
        .din(new_Jinkela_wire_8542),
        .dout(new_Jinkela_wire_8543)
    );

    spl2 new_Jinkela_splitter_321 (
        .a(n_0703_),
        .b(new_Jinkela_wire_5296),
        .c(new_Jinkela_wire_5297)
    );

    bfr new_Jinkela_buffer_6898 (
        .din(new_Jinkela_wire_8528),
        .dout(new_Jinkela_wire_8529)
    );

    bfr new_Jinkela_buffer_4423 (
        .din(new_Jinkela_wire_5262),
        .dout(new_Jinkela_wire_5263)
    );

    spl2 new_Jinkela_splitter_652 (
        .a(n_0314_),
        .b(new_Jinkela_wire_8571),
        .c(new_Jinkela_wire_8572)
    );

    bfr new_Jinkela_buffer_4443 (
        .din(n_1281_),
        .dout(new_Jinkela_wire_5298)
    );

    bfr new_Jinkela_buffer_4442 (
        .din(new_Jinkela_wire_5290),
        .dout(new_Jinkela_wire_5291)
    );

    bfr new_Jinkela_buffer_6899 (
        .din(new_Jinkela_wire_8529),
        .dout(new_Jinkela_wire_8530)
    );

    bfr new_Jinkela_buffer_4424 (
        .din(new_Jinkela_wire_5263),
        .dout(new_Jinkela_wire_5264)
    );

    bfr new_Jinkela_buffer_6913 (
        .din(new_Jinkela_wire_8543),
        .dout(new_Jinkela_wire_8544)
    );

    spl4L new_Jinkela_splitter_323 (
        .a(n_1167_),
        .d(new_Jinkela_wire_5364),
        .b(new_Jinkela_wire_5365),
        .e(new_Jinkela_wire_5366),
        .c(new_Jinkela_wire_5367)
    );

    bfr new_Jinkela_buffer_6900 (
        .din(new_Jinkela_wire_8530),
        .dout(new_Jinkela_wire_8531)
    );

    bfr new_Jinkela_buffer_4425 (
        .din(new_Jinkela_wire_5264),
        .dout(new_Jinkela_wire_5265)
    );

    bfr new_Jinkela_buffer_6938 (
        .din(new_Jinkela_wire_8572),
        .dout(new_Jinkela_wire_8573)
    );

    spl2 new_Jinkela_splitter_322 (
        .a(n_1312_),
        .b(new_Jinkela_wire_5343),
        .c(new_Jinkela_wire_5344)
    );

    bfr new_Jinkela_buffer_6901 (
        .din(new_Jinkela_wire_8531),
        .dout(new_Jinkela_wire_8532)
    );

    bfr new_Jinkela_buffer_4426 (
        .din(new_Jinkela_wire_5265),
        .dout(new_Jinkela_wire_5266)
    );

    bfr new_Jinkela_buffer_6914 (
        .din(new_Jinkela_wire_8544),
        .dout(new_Jinkela_wire_8545)
    );

    bfr new_Jinkela_buffer_4444 (
        .din(new_net_2513),
        .dout(new_Jinkela_wire_5299)
    );

    bfr new_Jinkela_buffer_4427 (
        .din(new_Jinkela_wire_5266),
        .dout(new_Jinkela_wire_5267)
    );

    spl2 new_Jinkela_splitter_654 (
        .a(new_net_5),
        .b(new_Jinkela_wire_8578),
        .c(new_Jinkela_wire_8579)
    );

    bfr new_Jinkela_buffer_6915 (
        .din(new_Jinkela_wire_8545),
        .dout(new_Jinkela_wire_8546)
    );

    bfr new_Jinkela_buffer_4445 (
        .din(new_Jinkela_wire_5299),
        .dout(new_Jinkela_wire_5300)
    );

    spl3L new_Jinkela_splitter_655 (
        .a(n_1330_),
        .d(new_Jinkela_wire_8624),
        .b(new_Jinkela_wire_8625),
        .c(new_Jinkela_wire_8626)
    );

    bfr new_Jinkela_buffer_4428 (
        .din(new_Jinkela_wire_5267),
        .dout(new_Jinkela_wire_5268)
    );

    bfr new_Jinkela_buffer_6939 (
        .din(new_Jinkela_wire_8579),
        .dout(new_Jinkela_wire_8580)
    );

    bfr new_Jinkela_buffer_6916 (
        .din(new_Jinkela_wire_8546),
        .dout(new_Jinkela_wire_8547)
    );

    bfr new_Jinkela_buffer_4488 (
        .din(new_Jinkela_wire_5344),
        .dout(new_Jinkela_wire_5345)
    );

    bfr new_Jinkela_buffer_4429 (
        .din(new_Jinkela_wire_5268),
        .dout(new_Jinkela_wire_5269)
    );

    bfr new_Jinkela_buffer_6917 (
        .din(new_Jinkela_wire_8547),
        .dout(new_Jinkela_wire_8548)
    );

    bfr new_Jinkela_buffer_4446 (
        .din(new_Jinkela_wire_5300),
        .dout(new_Jinkela_wire_5301)
    );

    bfr new_Jinkela_buffer_559 (
        .din(new_Jinkela_wire_602),
        .dout(new_Jinkela_wire_603)
    );

    bfr new_Jinkela_buffer_455 (
        .din(new_Jinkela_wire_491),
        .dout(new_Jinkela_wire_492)
    );

    bfr new_Jinkela_buffer_496 (
        .din(new_Jinkela_wire_537),
        .dout(new_Jinkela_wire_538)
    );

    bfr new_Jinkela_buffer_456 (
        .din(new_Jinkela_wire_492),
        .dout(new_Jinkela_wire_493)
    );

    bfr new_Jinkela_buffer_562 (
        .din(new_Jinkela_wire_605),
        .dout(new_Jinkela_wire_606)
    );

    bfr new_Jinkela_buffer_457 (
        .din(new_Jinkela_wire_493),
        .dout(new_Jinkela_wire_494)
    );

    bfr new_Jinkela_buffer_497 (
        .din(new_Jinkela_wire_538),
        .dout(new_Jinkela_wire_539)
    );

    bfr new_Jinkela_buffer_458 (
        .din(new_Jinkela_wire_494),
        .dout(new_Jinkela_wire_495)
    );

    bfr new_Jinkela_buffer_560 (
        .din(new_Jinkela_wire_603),
        .dout(new_Jinkela_wire_604)
    );

    bfr new_Jinkela_buffer_459 (
        .din(new_Jinkela_wire_495),
        .dout(new_Jinkela_wire_496)
    );

    bfr new_Jinkela_buffer_498 (
        .din(new_Jinkela_wire_539),
        .dout(new_Jinkela_wire_540)
    );

    bfr new_Jinkela_buffer_460 (
        .din(new_Jinkela_wire_496),
        .dout(new_Jinkela_wire_497)
    );

    bfr new_Jinkela_buffer_566 (
        .din(N260),
        .dout(new_Jinkela_wire_610)
    );

    bfr new_Jinkela_buffer_461 (
        .din(new_Jinkela_wire_497),
        .dout(new_Jinkela_wire_498)
    );

    bfr new_Jinkela_buffer_499 (
        .din(new_Jinkela_wire_540),
        .dout(new_Jinkela_wire_541)
    );

    bfr new_Jinkela_buffer_462 (
        .din(new_Jinkela_wire_498),
        .dout(new_Jinkela_wire_499)
    );

    bfr new_Jinkela_buffer_563 (
        .din(new_Jinkela_wire_606),
        .dout(new_Jinkela_wire_607)
    );

    bfr new_Jinkela_buffer_463 (
        .din(new_Jinkela_wire_499),
        .dout(new_Jinkela_wire_500)
    );

    bfr new_Jinkela_buffer_500 (
        .din(new_Jinkela_wire_541),
        .dout(new_Jinkela_wire_542)
    );

    bfr new_Jinkela_buffer_464 (
        .din(new_Jinkela_wire_500),
        .dout(new_Jinkela_wire_501)
    );

    bfr new_Jinkela_buffer_465 (
        .din(new_Jinkela_wire_501),
        .dout(new_Jinkela_wire_502)
    );

    bfr new_Jinkela_buffer_501 (
        .din(new_Jinkela_wire_542),
        .dout(new_Jinkela_wire_543)
    );

    bfr new_Jinkela_buffer_466 (
        .din(new_Jinkela_wire_502),
        .dout(new_Jinkela_wire_503)
    );

    bfr new_Jinkela_buffer_564 (
        .din(new_Jinkela_wire_607),
        .dout(new_Jinkela_wire_608)
    );

    bfr new_Jinkela_buffer_467 (
        .din(new_Jinkela_wire_503),
        .dout(new_Jinkela_wire_504)
    );

    bfr new_Jinkela_buffer_502 (
        .din(new_Jinkela_wire_543),
        .dout(new_Jinkela_wire_544)
    );

    bfr new_Jinkela_buffer_468 (
        .din(new_Jinkela_wire_504),
        .dout(new_Jinkela_wire_505)
    );

    bfr new_Jinkela_buffer_567 (
        .din(new_Jinkela_wire_610),
        .dout(new_Jinkela_wire_611)
    );

    bfr new_Jinkela_buffer_469 (
        .din(new_Jinkela_wire_505),
        .dout(new_Jinkela_wire_506)
    );

    bfr new_Jinkela_buffer_503 (
        .din(new_Jinkela_wire_544),
        .dout(new_Jinkela_wire_545)
    );

    bfr new_Jinkela_buffer_470 (
        .din(new_Jinkela_wire_506),
        .dout(new_Jinkela_wire_507)
    );

    bfr new_Jinkela_buffer_638 (
        .din(N198),
        .dout(new_Jinkela_wire_687)
    );

    bfr new_Jinkela_buffer_634 (
        .din(N158),
        .dout(new_Jinkela_wire_683)
    );

    bfr new_Jinkela_buffer_504 (
        .din(new_Jinkela_wire_545),
        .dout(new_Jinkela_wire_546)
    );

    bfr new_Jinkela_buffer_568 (
        .din(new_Jinkela_wire_611),
        .dout(new_Jinkela_wire_612)
    );

    bfr new_Jinkela_buffer_505 (
        .din(new_Jinkela_wire_546),
        .dout(new_Jinkela_wire_547)
    );

    bfr new_Jinkela_buffer_631 (
        .din(new_Jinkela_wire_679),
        .dout(new_Jinkela_wire_680)
    );

    bfr new_Jinkela_buffer_630 (
        .din(N189),
        .dout(new_Jinkela_wire_679)
    );

    bfr new_Jinkela_buffer_506 (
        .din(new_Jinkela_wire_547),
        .dout(new_Jinkela_wire_548)
    );

    bfr new_Jinkela_buffer_507 (
        .din(new_Jinkela_wire_548),
        .dout(new_Jinkela_wire_549)
    );

    spl2 new_Jinkela_splitter_19 (
        .a(new_Jinkela_wire_612),
        .b(new_Jinkela_wire_613),
        .c(new_Jinkela_wire_614)
    );

    bfr new_Jinkela_buffer_508 (
        .din(new_Jinkela_wire_549),
        .dout(new_Jinkela_wire_550)
    );

    bfr new_Jinkela_buffer_1991 (
        .din(new_Jinkela_wire_2355),
        .dout(new_Jinkela_wire_2356)
    );

    bfr new_Jinkela_buffer_1487 (
        .din(new_Jinkela_wire_1819),
        .dout(new_Jinkela_wire_1820)
    );

    bfr new_Jinkela_buffer_2730 (
        .din(new_Jinkela_wire_3144),
        .dout(new_Jinkela_wire_3145)
    );

    bfr new_Jinkela_buffer_2033 (
        .din(new_Jinkela_wire_2402),
        .dout(new_Jinkela_wire_2403)
    );

    bfr new_Jinkela_buffer_1421 (
        .din(new_Jinkela_wire_1753),
        .dout(new_Jinkela_wire_1754)
    );

    bfr new_Jinkela_buffer_2688 (
        .din(new_Jinkela_wire_3097),
        .dout(new_Jinkela_wire_3098)
    );

    bfr new_Jinkela_buffer_3553 (
        .din(new_Jinkela_wire_4150),
        .dout(new_Jinkela_wire_4151)
    );

    bfr new_Jinkela_buffer_1992 (
        .din(new_Jinkela_wire_2356),
        .dout(new_Jinkela_wire_2357)
    );

    bfr new_Jinkela_buffer_1485 (
        .din(new_Jinkela_wire_1817),
        .dout(new_Jinkela_wire_1818)
    );

    bfr new_Jinkela_buffer_2852 (
        .din(new_Jinkela_wire_3273),
        .dout(new_Jinkela_wire_3274)
    );

    bfr new_Jinkela_buffer_3591 (
        .din(new_Jinkela_wire_4197),
        .dout(new_Jinkela_wire_4198)
    );

    bfr new_Jinkela_buffer_3681 (
        .din(n_0003_),
        .dout(new_Jinkela_wire_4296)
    );

    bfr new_Jinkela_buffer_2105 (
        .din(N130),
        .dout(new_Jinkela_wire_2475)
    );

    bfr new_Jinkela_buffer_1422 (
        .din(new_Jinkela_wire_1754),
        .dout(new_Jinkela_wire_1755)
    );

    bfr new_Jinkela_buffer_2689 (
        .din(new_Jinkela_wire_3098),
        .dout(new_Jinkela_wire_3099)
    );

    bfr new_Jinkela_buffer_3554 (
        .din(new_Jinkela_wire_4151),
        .dout(new_Jinkela_wire_4152)
    );

    bfr new_Jinkela_buffer_1993 (
        .din(new_Jinkela_wire_2357),
        .dout(new_Jinkela_wire_2358)
    );

    bfr new_Jinkela_buffer_1494 (
        .din(N223),
        .dout(new_Jinkela_wire_1827)
    );

    bfr new_Jinkela_buffer_2731 (
        .din(new_Jinkela_wire_3145),
        .dout(new_Jinkela_wire_3146)
    );

    bfr new_Jinkela_buffer_3628 (
        .din(new_Jinkela_wire_4242),
        .dout(new_Jinkela_wire_4243)
    );

    bfr new_Jinkela_buffer_2034 (
        .din(new_Jinkela_wire_2403),
        .dout(new_Jinkela_wire_2404)
    );

    bfr new_Jinkela_buffer_1423 (
        .din(new_Jinkela_wire_1755),
        .dout(new_Jinkela_wire_1756)
    );

    bfr new_Jinkela_buffer_2690 (
        .din(new_Jinkela_wire_3099),
        .dout(new_Jinkela_wire_3100)
    );

    bfr new_Jinkela_buffer_3555 (
        .din(new_Jinkela_wire_4152),
        .dout(new_Jinkela_wire_4153)
    );

    bfr new_Jinkela_buffer_1994 (
        .din(new_Jinkela_wire_2358),
        .dout(new_Jinkela_wire_2359)
    );

    bfr new_Jinkela_buffer_1488 (
        .din(new_Jinkela_wire_1820),
        .dout(new_Jinkela_wire_1821)
    );

    bfr new_Jinkela_buffer_2791 (
        .din(new_Jinkela_wire_3207),
        .dout(new_Jinkela_wire_3208)
    );

    bfr new_Jinkela_buffer_3592 (
        .din(new_Jinkela_wire_4198),
        .dout(new_Jinkela_wire_4199)
    );

    bfr new_Jinkela_buffer_2099 (
        .din(new_Jinkela_wire_2468),
        .dout(new_Jinkela_wire_2469)
    );

    bfr new_Jinkela_buffer_1424 (
        .din(new_Jinkela_wire_1756),
        .dout(new_Jinkela_wire_1757)
    );

    bfr new_Jinkela_buffer_2691 (
        .din(new_Jinkela_wire_3100),
        .dout(new_Jinkela_wire_3101)
    );

    bfr new_Jinkela_buffer_3556 (
        .din(new_Jinkela_wire_4153),
        .dout(new_Jinkela_wire_4154)
    );

    bfr new_Jinkela_buffer_1995 (
        .din(new_Jinkela_wire_2359),
        .dout(new_Jinkela_wire_2360)
    );

    bfr new_Jinkela_buffer_1491 (
        .din(new_Jinkela_wire_1823),
        .dout(new_Jinkela_wire_1824)
    );

    bfr new_Jinkela_buffer_2732 (
        .din(new_Jinkela_wire_3146),
        .dout(new_Jinkela_wire_3147)
    );

    bfr new_Jinkela_buffer_2035 (
        .din(new_Jinkela_wire_2404),
        .dout(new_Jinkela_wire_2405)
    );

    bfr new_Jinkela_buffer_1425 (
        .din(new_Jinkela_wire_1757),
        .dout(new_Jinkela_wire_1758)
    );

    bfr new_Jinkela_buffer_2692 (
        .din(new_Jinkela_wire_3101),
        .dout(new_Jinkela_wire_3102)
    );

    bfr new_Jinkela_buffer_3557 (
        .din(new_Jinkela_wire_4154),
        .dout(new_Jinkela_wire_4155)
    );

    bfr new_Jinkela_buffer_1996 (
        .din(new_Jinkela_wire_2360),
        .dout(new_Jinkela_wire_2361)
    );

    bfr new_Jinkela_buffer_1489 (
        .din(new_Jinkela_wire_1821),
        .dout(new_Jinkela_wire_1822)
    );

    bfr new_Jinkela_buffer_2923 (
        .din(N23),
        .dout(new_Jinkela_wire_3347)
    );

    bfr new_Jinkela_buffer_3593 (
        .din(new_Jinkela_wire_4199),
        .dout(new_Jinkela_wire_4200)
    );

    bfr new_Jinkela_buffer_3664 (
        .din(new_Jinkela_wire_4278),
        .dout(new_Jinkela_wire_4279)
    );

    bfr new_Jinkela_buffer_2102 (
        .din(new_Jinkela_wire_2471),
        .dout(new_Jinkela_wire_2472)
    );

    bfr new_Jinkela_buffer_1426 (
        .din(new_Jinkela_wire_1758),
        .dout(new_Jinkela_wire_1759)
    );

    bfr new_Jinkela_buffer_2693 (
        .din(new_Jinkela_wire_3102),
        .dout(new_Jinkela_wire_3103)
    );

    bfr new_Jinkela_buffer_3558 (
        .din(new_Jinkela_wire_4155),
        .dout(new_Jinkela_wire_4156)
    );

    bfr new_Jinkela_buffer_1997 (
        .din(new_Jinkela_wire_2361),
        .dout(new_Jinkela_wire_2362)
    );

    bfr new_Jinkela_buffer_1498 (
        .din(N106),
        .dout(new_Jinkela_wire_1831)
    );

    bfr new_Jinkela_buffer_2733 (
        .din(new_Jinkela_wire_3147),
        .dout(new_Jinkela_wire_3148)
    );

    bfr new_Jinkela_buffer_3629 (
        .din(new_Jinkela_wire_4243),
        .dout(new_Jinkela_wire_4244)
    );

    bfr new_Jinkela_buffer_2036 (
        .din(new_Jinkela_wire_2405),
        .dout(new_Jinkela_wire_2406)
    );

    bfr new_Jinkela_buffer_1427 (
        .din(new_Jinkela_wire_1759),
        .dout(new_Jinkela_wire_1760)
    );

    bfr new_Jinkela_buffer_2694 (
        .din(new_Jinkela_wire_3103),
        .dout(new_Jinkela_wire_3104)
    );

    bfr new_Jinkela_buffer_3559 (
        .din(new_Jinkela_wire_4156),
        .dout(new_Jinkela_wire_4157)
    );

    bfr new_Jinkela_buffer_1998 (
        .din(new_Jinkela_wire_2362),
        .dout(new_Jinkela_wire_2363)
    );

    bfr new_Jinkela_buffer_1492 (
        .din(new_Jinkela_wire_1824),
        .dout(new_Jinkela_wire_1825)
    );

    bfr new_Jinkela_buffer_2792 (
        .din(new_Jinkela_wire_3208),
        .dout(new_Jinkela_wire_3209)
    );

    bfr new_Jinkela_buffer_3594 (
        .din(new_Jinkela_wire_4200),
        .dout(new_Jinkela_wire_4201)
    );

    bfr new_Jinkela_buffer_2100 (
        .din(new_Jinkela_wire_2469),
        .dout(new_Jinkela_wire_2470)
    );

    bfr new_Jinkela_buffer_1428 (
        .din(new_Jinkela_wire_1760),
        .dout(new_Jinkela_wire_1761)
    );

    bfr new_Jinkela_buffer_2695 (
        .din(new_Jinkela_wire_3104),
        .dout(new_Jinkela_wire_3105)
    );

    bfr new_Jinkela_buffer_3560 (
        .din(new_Jinkela_wire_4157),
        .dout(new_Jinkela_wire_4158)
    );

    bfr new_Jinkela_buffer_1999 (
        .din(new_Jinkela_wire_2363),
        .dout(new_Jinkela_wire_2364)
    );

    bfr new_Jinkela_buffer_1495 (
        .din(new_Jinkela_wire_1827),
        .dout(new_Jinkela_wire_1828)
    );

    bfr new_Jinkela_buffer_2734 (
        .din(new_Jinkela_wire_3148),
        .dout(new_Jinkela_wire_3149)
    );

    bfr new_Jinkela_buffer_2037 (
        .din(new_Jinkela_wire_2406),
        .dout(new_Jinkela_wire_2407)
    );

    bfr new_Jinkela_buffer_1429 (
        .din(new_Jinkela_wire_1761),
        .dout(new_Jinkela_wire_1762)
    );

    bfr new_Jinkela_buffer_2696 (
        .din(new_Jinkela_wire_3105),
        .dout(new_Jinkela_wire_3106)
    );

    bfr new_Jinkela_buffer_3561 (
        .din(new_Jinkela_wire_4158),
        .dout(new_Jinkela_wire_4159)
    );

    bfr new_Jinkela_buffer_2000 (
        .din(new_Jinkela_wire_2364),
        .dout(new_Jinkela_wire_2365)
    );

    bfr new_Jinkela_buffer_1493 (
        .din(new_Jinkela_wire_1825),
        .dout(new_Jinkela_wire_1826)
    );

    spl2 new_Jinkela_splitter_143 (
        .a(new_Jinkela_wire_3274),
        .b(new_Jinkela_wire_3275),
        .c(new_Jinkela_wire_3276)
    );

    bfr new_Jinkela_buffer_3595 (
        .din(new_Jinkela_wire_4201),
        .dout(new_Jinkela_wire_4202)
    );

    bfr new_Jinkela_buffer_3668 (
        .din(new_Jinkela_wire_4282),
        .dout(new_Jinkela_wire_4283)
    );

    bfr new_Jinkela_buffer_2109 (
        .din(N257),
        .dout(new_Jinkela_wire_2479)
    );

    bfr new_Jinkela_buffer_1430 (
        .din(new_Jinkela_wire_1762),
        .dout(new_Jinkela_wire_1763)
    );

    bfr new_Jinkela_buffer_2697 (
        .din(new_Jinkela_wire_3106),
        .dout(new_Jinkela_wire_3107)
    );

    bfr new_Jinkela_buffer_3562 (
        .din(new_Jinkela_wire_4159),
        .dout(new_Jinkela_wire_4160)
    );

    bfr new_Jinkela_buffer_2735 (
        .din(new_Jinkela_wire_3149),
        .dout(new_Jinkela_wire_3150)
    );

    bfr new_Jinkela_buffer_2001 (
        .din(new_Jinkela_wire_2365),
        .dout(new_Jinkela_wire_2366)
    );

    bfr new_Jinkela_buffer_1630 (
        .din(N74),
        .dout(new_Jinkela_wire_1974)
    );

    bfr new_Jinkela_buffer_3630 (
        .din(new_Jinkela_wire_4244),
        .dout(new_Jinkela_wire_4245)
    );

    bfr new_Jinkela_buffer_2038 (
        .din(new_Jinkela_wire_2407),
        .dout(new_Jinkela_wire_2408)
    );

    bfr new_Jinkela_buffer_1431 (
        .din(new_Jinkela_wire_1763),
        .dout(new_Jinkela_wire_1764)
    );

    bfr new_Jinkela_buffer_2698 (
        .din(new_Jinkela_wire_3107),
        .dout(new_Jinkela_wire_3108)
    );

    bfr new_Jinkela_buffer_3563 (
        .din(new_Jinkela_wire_4160),
        .dout(new_Jinkela_wire_4161)
    );

    bfr new_Jinkela_buffer_2002 (
        .din(new_Jinkela_wire_2366),
        .dout(new_Jinkela_wire_2367)
    );

    bfr new_Jinkela_buffer_1496 (
        .din(new_Jinkela_wire_1828),
        .dout(new_Jinkela_wire_1829)
    );

    spl3L new_Jinkela_splitter_141 (
        .a(new_Jinkela_wire_3209),
        .d(new_Jinkela_wire_3210),
        .b(new_Jinkela_wire_3211),
        .c(new_Jinkela_wire_3212)
    );

    bfr new_Jinkela_buffer_3596 (
        .din(new_Jinkela_wire_4202),
        .dout(new_Jinkela_wire_4203)
    );

    bfr new_Jinkela_buffer_2103 (
        .din(new_Jinkela_wire_2472),
        .dout(new_Jinkela_wire_2473)
    );

    bfr new_Jinkela_buffer_1432 (
        .din(new_Jinkela_wire_1764),
        .dout(new_Jinkela_wire_1765)
    );

    bfr new_Jinkela_buffer_2699 (
        .din(new_Jinkela_wire_3108),
        .dout(new_Jinkela_wire_3109)
    );

    bfr new_Jinkela_buffer_3564 (
        .din(new_Jinkela_wire_4161),
        .dout(new_Jinkela_wire_4162)
    );

    bfr new_Jinkela_buffer_2003 (
        .din(new_Jinkela_wire_2367),
        .dout(new_Jinkela_wire_2368)
    );

    bfr new_Jinkela_buffer_1499 (
        .din(new_Jinkela_wire_1831),
        .dout(new_Jinkela_wire_1832)
    );

    bfr new_Jinkela_buffer_2736 (
        .din(new_Jinkela_wire_3150),
        .dout(new_Jinkela_wire_3151)
    );

    bfr new_Jinkela_buffer_2039 (
        .din(new_Jinkela_wire_2408),
        .dout(new_Jinkela_wire_2409)
    );

    bfr new_Jinkela_buffer_1433 (
        .din(new_Jinkela_wire_1765),
        .dout(new_Jinkela_wire_1766)
    );

    bfr new_Jinkela_buffer_2700 (
        .din(new_Jinkela_wire_3109),
        .dout(new_Jinkela_wire_3110)
    );

    bfr new_Jinkela_buffer_3565 (
        .din(new_Jinkela_wire_4162),
        .dout(new_Jinkela_wire_4163)
    );

    bfr new_Jinkela_buffer_2004 (
        .din(new_Jinkela_wire_2368),
        .dout(new_Jinkela_wire_2369)
    );

    bfr new_Jinkela_buffer_1497 (
        .din(new_Jinkela_wire_1829),
        .dout(new_Jinkela_wire_1830)
    );

    bfr new_Jinkela_buffer_2853 (
        .din(new_Jinkela_wire_3276),
        .dout(new_Jinkela_wire_3277)
    );

    bfr new_Jinkela_buffer_3597 (
        .din(new_Jinkela_wire_4203),
        .dout(new_Jinkela_wire_4204)
    );

    bfr new_Jinkela_buffer_3665 (
        .din(new_Jinkela_wire_4279),
        .dout(new_Jinkela_wire_4280)
    );

    bfr new_Jinkela_buffer_2106 (
        .din(new_Jinkela_wire_2475),
        .dout(new_Jinkela_wire_2476)
    );

    bfr new_Jinkela_buffer_1434 (
        .din(new_Jinkela_wire_1766),
        .dout(new_Jinkela_wire_1767)
    );

    bfr new_Jinkela_buffer_2701 (
        .din(new_Jinkela_wire_3110),
        .dout(new_Jinkela_wire_3111)
    );

    bfr new_Jinkela_buffer_3566 (
        .din(new_Jinkela_wire_4163),
        .dout(new_Jinkela_wire_4164)
    );

    bfr new_Jinkela_buffer_2737 (
        .din(new_Jinkela_wire_3151),
        .dout(new_Jinkela_wire_3152)
    );

    bfr new_Jinkela_buffer_2005 (
        .din(new_Jinkela_wire_2369),
        .dout(new_Jinkela_wire_2370)
    );

    spl4L new_Jinkela_splitter_107 (
        .a(N263),
        .d(new_Jinkela_wire_1904),
        .b(new_Jinkela_wire_1905),
        .e(new_Jinkela_wire_1906),
        .c(new_Jinkela_wire_1907)
    );

    bfr new_Jinkela_buffer_3631 (
        .din(new_Jinkela_wire_4245),
        .dout(new_Jinkela_wire_4246)
    );

    bfr new_Jinkela_buffer_2040 (
        .din(new_Jinkela_wire_2409),
        .dout(new_Jinkela_wire_2410)
    );

    bfr new_Jinkela_buffer_1435 (
        .din(new_Jinkela_wire_1767),
        .dout(new_Jinkela_wire_1768)
    );

    bfr new_Jinkela_buffer_2702 (
        .din(new_Jinkela_wire_3111),
        .dout(new_Jinkela_wire_3112)
    );

    bfr new_Jinkela_buffer_3567 (
        .din(new_Jinkela_wire_4164),
        .dout(new_Jinkela_wire_4165)
    );

    bfr new_Jinkela_buffer_2006 (
        .din(new_Jinkela_wire_2370),
        .dout(new_Jinkela_wire_2371)
    );

    bfr new_Jinkela_buffer_1500 (
        .din(new_Jinkela_wire_1832),
        .dout(new_Jinkela_wire_1833)
    );

    bfr new_Jinkela_buffer_2793 (
        .din(new_Jinkela_wire_3212),
        .dout(new_Jinkela_wire_3213)
    );

    bfr new_Jinkela_buffer_3598 (
        .din(new_Jinkela_wire_4204),
        .dout(new_Jinkela_wire_4205)
    );

    bfr new_Jinkela_buffer_2104 (
        .din(new_Jinkela_wire_2473),
        .dout(new_Jinkela_wire_2474)
    );

    bfr new_Jinkela_buffer_1436 (
        .din(new_Jinkela_wire_1768),
        .dout(new_Jinkela_wire_1769)
    );

    bfr new_Jinkela_buffer_2703 (
        .din(new_Jinkela_wire_3112),
        .dout(new_Jinkela_wire_3113)
    );

    bfr new_Jinkela_buffer_3568 (
        .din(new_Jinkela_wire_4165),
        .dout(new_Jinkela_wire_4166)
    );

    bfr new_Jinkela_buffer_2007 (
        .din(new_Jinkela_wire_2371),
        .dout(new_Jinkela_wire_2372)
    );

    bfr new_Jinkela_buffer_1563 (
        .din(new_Jinkela_wire_1900),
        .dout(new_Jinkela_wire_1901)
    );

    bfr new_Jinkela_buffer_2738 (
        .din(new_Jinkela_wire_3152),
        .dout(new_Jinkela_wire_3153)
    );

    bfr new_Jinkela_buffer_1562 (
        .din(N73),
        .dout(new_Jinkela_wire_1900)
    );

    bfr new_Jinkela_buffer_2041 (
        .din(new_Jinkela_wire_2410),
        .dout(new_Jinkela_wire_2411)
    );

    bfr new_Jinkela_buffer_1437 (
        .din(new_Jinkela_wire_1769),
        .dout(new_Jinkela_wire_1770)
    );

    bfr new_Jinkela_buffer_2704 (
        .din(new_Jinkela_wire_3113),
        .dout(new_Jinkela_wire_3114)
    );

    bfr new_Jinkela_buffer_3569 (
        .din(new_Jinkela_wire_4166),
        .dout(new_Jinkela_wire_4167)
    );

    bfr new_Jinkela_buffer_2008 (
        .din(new_Jinkela_wire_2372),
        .dout(new_Jinkela_wire_2373)
    );

    spl2 new_Jinkela_splitter_105 (
        .a(new_Jinkela_wire_1833),
        .b(new_Jinkela_wire_1834),
        .c(new_Jinkela_wire_1835)
    );

    bfr new_Jinkela_buffer_2917 (
        .din(new_Jinkela_wire_3340),
        .dout(new_Jinkela_wire_3341)
    );

    bfr new_Jinkela_buffer_3599 (
        .din(new_Jinkela_wire_4205),
        .dout(new_Jinkela_wire_4206)
    );

    spl4L new_Jinkela_splitter_222 (
        .a(n_1308_),
        .d(new_Jinkela_wire_4307),
        .b(new_Jinkela_wire_4308),
        .e(new_Jinkela_wire_4309),
        .c(new_Jinkela_wire_4310)
    );

    bfr new_Jinkela_buffer_2705 (
        .din(new_Jinkela_wire_3114),
        .dout(new_Jinkela_wire_3115)
    );

    bfr new_Jinkela_buffer_1438 (
        .din(new_Jinkela_wire_1770),
        .dout(new_Jinkela_wire_1771)
    );

    bfr new_Jinkela_buffer_3570 (
        .din(new_Jinkela_wire_4167),
        .dout(new_Jinkela_wire_4168)
    );

    bfr new_Jinkela_buffer_2177 (
        .din(N200),
        .dout(new_Jinkela_wire_2552)
    );

    bfr new_Jinkela_buffer_2042 (
        .din(new_Jinkela_wire_2411),
        .dout(new_Jinkela_wire_2412)
    );

    bfr new_Jinkela_buffer_1501 (
        .din(new_Jinkela_wire_1835),
        .dout(new_Jinkela_wire_1836)
    );

    bfr new_Jinkela_buffer_2739 (
        .din(new_Jinkela_wire_3153),
        .dout(new_Jinkela_wire_3154)
    );

    bfr new_Jinkela_buffer_3632 (
        .din(new_Jinkela_wire_4246),
        .dout(new_Jinkela_wire_4247)
    );

    bfr new_Jinkela_buffer_2107 (
        .din(new_Jinkela_wire_2476),
        .dout(new_Jinkela_wire_2477)
    );

    bfr new_Jinkela_buffer_1439 (
        .din(new_Jinkela_wire_1771),
        .dout(new_Jinkela_wire_1772)
    );

    bfr new_Jinkela_buffer_2706 (
        .din(new_Jinkela_wire_3115),
        .dout(new_Jinkela_wire_3116)
    );

    bfr new_Jinkela_buffer_3571 (
        .din(new_Jinkela_wire_4168),
        .dout(new_Jinkela_wire_4169)
    );

    bfr new_Jinkela_buffer_2794 (
        .din(new_Jinkela_wire_3213),
        .dout(new_Jinkela_wire_3214)
    );

    bfr new_Jinkela_buffer_2043 (
        .din(new_Jinkela_wire_2412),
        .dout(new_Jinkela_wire_2413)
    );

    bfr new_Jinkela_buffer_3600 (
        .din(new_Jinkela_wire_4206),
        .dout(new_Jinkela_wire_4207)
    );

    bfr new_Jinkela_buffer_2173 (
        .din(N62),
        .dout(new_Jinkela_wire_2548)
    );

    bfr new_Jinkela_buffer_1440 (
        .din(new_Jinkela_wire_1772),
        .dout(new_Jinkela_wire_1773)
    );

    bfr new_Jinkela_buffer_2740 (
        .din(new_Jinkela_wire_3154),
        .dout(new_Jinkela_wire_3155)
    );

    bfr new_Jinkela_buffer_3572 (
        .din(new_Jinkela_wire_4169),
        .dout(new_Jinkela_wire_4170)
    );

    bfr new_Jinkela_buffer_2044 (
        .din(new_Jinkela_wire_2413),
        .dout(new_Jinkela_wire_2414)
    );

    bfr new_Jinkela_buffer_1564 (
        .din(new_Jinkela_wire_1901),
        .dout(new_Jinkela_wire_1902)
    );

    bfr new_Jinkela_buffer_2920 (
        .din(new_Jinkela_wire_3343),
        .dout(new_Jinkela_wire_3344)
    );

    spl2 new_Jinkela_splitter_223 (
        .a(n_0759_),
        .b(new_Jinkela_wire_4337),
        .c(new_Jinkela_wire_4338)
    );

    bfr new_Jinkela_buffer_2108 (
        .din(new_Jinkela_wire_2477),
        .dout(new_Jinkela_wire_2478)
    );

    bfr new_Jinkela_buffer_1441 (
        .din(new_Jinkela_wire_1773),
        .dout(new_Jinkela_wire_1774)
    );

    bfr new_Jinkela_buffer_2741 (
        .din(new_Jinkela_wire_3155),
        .dout(new_Jinkela_wire_3156)
    );

    bfr new_Jinkela_buffer_3601 (
        .din(new_Jinkela_wire_4207),
        .dout(new_Jinkela_wire_4208)
    );

    bfr new_Jinkela_buffer_3666 (
        .din(new_Jinkela_wire_4280),
        .dout(new_Jinkela_wire_4281)
    );

    bfr new_Jinkela_buffer_6173 (
        .din(n_0760_),
        .dout(new_Jinkela_wire_7541)
    );

    spl2 new_Jinkela_splitter_535 (
        .a(n_0223_),
        .b(new_Jinkela_wire_7500),
        .c(new_Jinkela_wire_7501)
    );

    spl2 new_Jinkela_splitter_524 (
        .a(new_Jinkela_wire_7403),
        .b(new_Jinkela_wire_7404),
        .c(new_Jinkela_wire_7405)
    );

    spl4L new_Jinkela_splitter_534 (
        .a(n_1294_),
        .d(new_Jinkela_wire_7461),
        .b(new_Jinkela_wire_7462),
        .e(new_Jinkela_wire_7463),
        .c(new_Jinkela_wire_7464)
    );

    bfr new_Jinkela_buffer_6079 (
        .din(new_Jinkela_wire_7422),
        .dout(new_Jinkela_wire_7423)
    );

    bfr new_Jinkela_buffer_6080 (
        .din(new_Jinkela_wire_7423),
        .dout(new_Jinkela_wire_7424)
    );

    bfr new_Jinkela_buffer_6103 (
        .din(new_Jinkela_wire_7464),
        .dout(new_Jinkela_wire_7465)
    );

    bfr new_Jinkela_buffer_6081 (
        .din(new_Jinkela_wire_7424),
        .dout(new_Jinkela_wire_7425)
    );

    bfr new_Jinkela_buffer_6082 (
        .din(new_Jinkela_wire_7425),
        .dout(new_Jinkela_wire_7426)
    );

    spl2 new_Jinkela_splitter_536 (
        .a(n_0372_),
        .b(new_Jinkela_wire_7503),
        .c(new_Jinkela_wire_7504)
    );

    bfr new_Jinkela_buffer_6083 (
        .din(new_Jinkela_wire_7426),
        .dout(new_Jinkela_wire_7427)
    );

    bfr new_Jinkela_buffer_6104 (
        .din(new_Jinkela_wire_7465),
        .dout(new_Jinkela_wire_7466)
    );

    bfr new_Jinkela_buffer_6084 (
        .din(new_Jinkela_wire_7427),
        .dout(new_Jinkela_wire_7428)
    );

    bfr new_Jinkela_buffer_6138 (
        .din(new_Jinkela_wire_7501),
        .dout(new_Jinkela_wire_7502)
    );

    bfr new_Jinkela_buffer_6085 (
        .din(new_Jinkela_wire_7428),
        .dout(new_Jinkela_wire_7429)
    );

    bfr new_Jinkela_buffer_6105 (
        .din(new_Jinkela_wire_7466),
        .dout(new_Jinkela_wire_7467)
    );

    bfr new_Jinkela_buffer_6086 (
        .din(new_Jinkela_wire_7429),
        .dout(new_Jinkela_wire_7430)
    );

    bfr new_Jinkela_buffer_6087 (
        .din(new_Jinkela_wire_7430),
        .dout(new_Jinkela_wire_7431)
    );

    bfr new_Jinkela_buffer_6106 (
        .din(new_Jinkela_wire_7467),
        .dout(new_Jinkela_wire_7468)
    );

    bfr new_Jinkela_buffer_6088 (
        .din(new_Jinkela_wire_7431),
        .dout(new_Jinkela_wire_7432)
    );

    bfr new_Jinkela_buffer_6174 (
        .din(n_0305_),
        .dout(new_Jinkela_wire_7542)
    );

    bfr new_Jinkela_buffer_6139 (
        .din(new_Jinkela_wire_7504),
        .dout(new_Jinkela_wire_7505)
    );

    bfr new_Jinkela_buffer_6089 (
        .din(new_Jinkela_wire_7432),
        .dout(new_Jinkela_wire_7433)
    );

    bfr new_Jinkela_buffer_6107 (
        .din(new_Jinkela_wire_7468),
        .dout(new_Jinkela_wire_7469)
    );

    bfr new_Jinkela_buffer_6090 (
        .din(new_Jinkela_wire_7433),
        .dout(new_Jinkela_wire_7434)
    );

    spl2 new_Jinkela_splitter_538 (
        .a(n_0155_),
        .b(new_Jinkela_wire_7543),
        .c(new_Jinkela_wire_7544)
    );

    bfr new_Jinkela_buffer_6091 (
        .din(new_Jinkela_wire_7434),
        .dout(new_Jinkela_wire_7435)
    );

    bfr new_Jinkela_buffer_6108 (
        .din(new_Jinkela_wire_7469),
        .dout(new_Jinkela_wire_7470)
    );

    bfr new_Jinkela_buffer_6092 (
        .din(new_Jinkela_wire_7435),
        .dout(new_Jinkela_wire_7436)
    );

    spl2 new_Jinkela_splitter_539 (
        .a(n_0114_),
        .b(new_Jinkela_wire_7545),
        .c(new_Jinkela_wire_7546)
    );

    bfr new_Jinkela_buffer_6140 (
        .din(new_Jinkela_wire_7505),
        .dout(new_Jinkela_wire_7506)
    );

    bfr new_Jinkela_buffer_6093 (
        .din(new_Jinkela_wire_7436),
        .dout(new_Jinkela_wire_7437)
    );

    bfr new_Jinkela_buffer_6109 (
        .din(new_Jinkela_wire_7470),
        .dout(new_Jinkela_wire_7471)
    );

    bfr new_Jinkela_buffer_6094 (
        .din(new_Jinkela_wire_7437),
        .dout(new_Jinkela_wire_7438)
    );

    bfr new_Jinkela_buffer_6095 (
        .din(new_Jinkela_wire_7438),
        .dout(new_Jinkela_wire_7439)
    );

    bfr new_Jinkela_buffer_6110 (
        .din(new_Jinkela_wire_7471),
        .dout(new_Jinkela_wire_7472)
    );

    bfr new_Jinkela_buffer_6096 (
        .din(new_Jinkela_wire_7439),
        .dout(new_Jinkela_wire_7440)
    );

    bfr new_Jinkela_buffer_6141 (
        .din(new_Jinkela_wire_7506),
        .dout(new_Jinkela_wire_7507)
    );

    bfr new_Jinkela_buffer_6097 (
        .din(new_Jinkela_wire_7440),
        .dout(new_Jinkela_wire_7441)
    );

    bfr new_Jinkela_buffer_6111 (
        .din(new_Jinkela_wire_7472),
        .dout(new_Jinkela_wire_7473)
    );

    bfr new_Jinkela_buffer_6098 (
        .din(new_Jinkela_wire_7441),
        .dout(new_Jinkela_wire_7442)
    );

    bfr new_Jinkela_buffer_5299 (
        .din(new_Jinkela_wire_6357),
        .dout(new_Jinkela_wire_6358)
    );

    bfr new_Jinkela_buffer_5287 (
        .din(new_Jinkela_wire_6343),
        .dout(new_Jinkela_wire_6344)
    );

    bfr new_Jinkela_buffer_7983 (
        .din(new_Jinkela_wire_10055),
        .dout(new_Jinkela_wire_10056)
    );

    bfr new_Jinkela_buffer_5260 (
        .din(new_Jinkela_wire_6294),
        .dout(new_Jinkela_wire_6295)
    );

    bfr new_Jinkela_buffer_8034 (
        .din(new_Jinkela_wire_10114),
        .dout(new_Jinkela_wire_10115)
    );

    bfr new_Jinkela_buffer_7984 (
        .din(new_Jinkela_wire_10056),
        .dout(new_Jinkela_wire_10057)
    );

    bfr new_Jinkela_buffer_5261 (
        .din(new_Jinkela_wire_6295),
        .dout(new_Jinkela_wire_6296)
    );

    bfr new_Jinkela_buffer_5332 (
        .din(new_Jinkela_wire_6394),
        .dout(new_Jinkela_wire_6395)
    );

    bfr new_Jinkela_buffer_5288 (
        .din(new_Jinkela_wire_6344),
        .dout(new_Jinkela_wire_6345)
    );

    bfr new_Jinkela_buffer_7985 (
        .din(new_Jinkela_wire_10057),
        .dout(new_Jinkela_wire_10058)
    );

    bfr new_Jinkela_buffer_5262 (
        .din(new_Jinkela_wire_6296),
        .dout(new_Jinkela_wire_6297)
    );

    bfr new_Jinkela_buffer_8124 (
        .din(n_0948_),
        .dout(new_Jinkela_wire_10219)
    );

    bfr new_Jinkela_buffer_8035 (
        .din(new_Jinkela_wire_10115),
        .dout(new_Jinkela_wire_10116)
    );

    bfr new_Jinkela_buffer_5354 (
        .din(n_0768_),
        .dout(new_Jinkela_wire_6428)
    );

    bfr new_Jinkela_buffer_7986 (
        .din(new_Jinkela_wire_10058),
        .dout(new_Jinkela_wire_10059)
    );

    bfr new_Jinkela_buffer_5263 (
        .din(new_Jinkela_wire_6297),
        .dout(new_Jinkela_wire_6298)
    );

    bfr new_Jinkela_buffer_8058 (
        .din(new_Jinkela_wire_10150),
        .dout(new_Jinkela_wire_10151)
    );

    bfr new_Jinkela_buffer_5300 (
        .din(new_Jinkela_wire_6358),
        .dout(new_Jinkela_wire_6359)
    );

    bfr new_Jinkela_buffer_5289 (
        .din(new_Jinkela_wire_6345),
        .dout(new_Jinkela_wire_6346)
    );

    bfr new_Jinkela_buffer_7987 (
        .din(new_Jinkela_wire_10059),
        .dout(new_Jinkela_wire_10060)
    );

    bfr new_Jinkela_buffer_5264 (
        .din(new_Jinkela_wire_6298),
        .dout(new_Jinkela_wire_6299)
    );

    bfr new_Jinkela_buffer_8036 (
        .din(new_Jinkela_wire_10116),
        .dout(new_Jinkela_wire_10117)
    );

    bfr new_Jinkela_buffer_7988 (
        .din(new_Jinkela_wire_10060),
        .dout(new_Jinkela_wire_10061)
    );

    bfr new_Jinkela_buffer_5265 (
        .din(new_Jinkela_wire_6299),
        .dout(new_Jinkela_wire_6300)
    );

    bfr new_Jinkela_buffer_8061 (
        .din(new_Jinkela_wire_10155),
        .dout(new_Jinkela_wire_10156)
    );

    bfr new_Jinkela_buffer_5290 (
        .din(new_Jinkela_wire_6346),
        .dout(new_Jinkela_wire_6347)
    );

    bfr new_Jinkela_buffer_7989 (
        .din(new_Jinkela_wire_10061),
        .dout(new_Jinkela_wire_10062)
    );

    bfr new_Jinkela_buffer_5266 (
        .din(new_Jinkela_wire_6300),
        .dout(new_Jinkela_wire_6301)
    );

    bfr new_Jinkela_buffer_8127 (
        .din(n_1111_),
        .dout(new_Jinkela_wire_10222)
    );

    bfr new_Jinkela_buffer_8037 (
        .din(new_Jinkela_wire_10117),
        .dout(new_Jinkela_wire_10118)
    );

    spl2 new_Jinkela_splitter_413 (
        .a(n_1351_),
        .b(new_Jinkela_wire_6403),
        .c(new_Jinkela_wire_6405)
    );

    bfr new_Jinkela_buffer_7990 (
        .din(new_Jinkela_wire_10062),
        .dout(new_Jinkela_wire_10063)
    );

    bfr new_Jinkela_buffer_5267 (
        .din(new_Jinkela_wire_6301),
        .dout(new_Jinkela_wire_6302)
    );

    bfr new_Jinkela_buffer_8059 (
        .din(new_Jinkela_wire_10151),
        .dout(new_Jinkela_wire_10152)
    );

    bfr new_Jinkela_buffer_5301 (
        .din(new_Jinkela_wire_6359),
        .dout(new_Jinkela_wire_6360)
    );

    bfr new_Jinkela_buffer_5291 (
        .din(new_Jinkela_wire_6347),
        .dout(new_Jinkela_wire_6348)
    );

    bfr new_Jinkela_buffer_7991 (
        .din(new_Jinkela_wire_10063),
        .dout(new_Jinkela_wire_10064)
    );

    bfr new_Jinkela_buffer_5268 (
        .din(new_Jinkela_wire_6302),
        .dout(new_Jinkela_wire_6303)
    );

    bfr new_Jinkela_buffer_8038 (
        .din(new_Jinkela_wire_10118),
        .dout(new_Jinkela_wire_10119)
    );

    bfr new_Jinkela_buffer_7992 (
        .din(new_Jinkela_wire_10064),
        .dout(new_Jinkela_wire_10065)
    );

    bfr new_Jinkela_buffer_5269 (
        .din(new_Jinkela_wire_6303),
        .dout(new_Jinkela_wire_6304)
    );

    spl2 new_Jinkela_splitter_843 (
        .a(new_net_2),
        .b(new_Jinkela_wire_10229),
        .c(new_Jinkela_wire_10230)
    );

    spl3L new_Jinkela_splitter_411 (
        .a(n_0972_),
        .d(new_Jinkela_wire_6398),
        .b(new_Jinkela_wire_6399),
        .c(new_Jinkela_wire_6400)
    );

    bfr new_Jinkela_buffer_5292 (
        .din(new_Jinkela_wire_6348),
        .dout(new_Jinkela_wire_6349)
    );

    bfr new_Jinkela_buffer_7993 (
        .din(new_Jinkela_wire_10065),
        .dout(new_Jinkela_wire_10066)
    );

    bfr new_Jinkela_buffer_5270 (
        .din(new_Jinkela_wire_6304),
        .dout(new_Jinkela_wire_6305)
    );

    bfr new_Jinkela_buffer_8125 (
        .din(new_Jinkela_wire_10219),
        .dout(new_Jinkela_wire_10220)
    );

    bfr new_Jinkela_buffer_8039 (
        .din(new_Jinkela_wire_10119),
        .dout(new_Jinkela_wire_10120)
    );

    bfr new_Jinkela_buffer_7994 (
        .din(new_Jinkela_wire_10066),
        .dout(new_Jinkela_wire_10067)
    );

    bfr new_Jinkela_buffer_5271 (
        .din(new_Jinkela_wire_6305),
        .dout(new_Jinkela_wire_6306)
    );

    bfr new_Jinkela_buffer_8060 (
        .din(new_Jinkela_wire_10152),
        .dout(new_Jinkela_wire_10153)
    );

    bfr new_Jinkela_buffer_5302 (
        .din(new_Jinkela_wire_6360),
        .dout(new_Jinkela_wire_6361)
    );

    bfr new_Jinkela_buffer_5293 (
        .din(new_Jinkela_wire_6349),
        .dout(new_Jinkela_wire_6350)
    );

    bfr new_Jinkela_buffer_7995 (
        .din(new_Jinkela_wire_10067),
        .dout(new_Jinkela_wire_10068)
    );

    bfr new_Jinkela_buffer_5272 (
        .din(new_Jinkela_wire_6306),
        .dout(new_Jinkela_wire_6307)
    );

    bfr new_Jinkela_buffer_8040 (
        .din(new_Jinkela_wire_10120),
        .dout(new_Jinkela_wire_10121)
    );

    bfr new_Jinkela_buffer_7996 (
        .din(new_Jinkela_wire_10068),
        .dout(new_Jinkela_wire_10069)
    );

    bfr new_Jinkela_buffer_5333 (
        .din(new_Jinkela_wire_6395),
        .dout(new_Jinkela_wire_6396)
    );

    bfr new_Jinkela_buffer_5294 (
        .din(new_Jinkela_wire_6350),
        .dout(new_Jinkela_wire_6351)
    );

    bfr new_Jinkela_buffer_8062 (
        .din(new_Jinkela_wire_10156),
        .dout(new_Jinkela_wire_10157)
    );

    bfr new_Jinkela_buffer_7997 (
        .din(new_Jinkela_wire_10069),
        .dout(new_Jinkela_wire_10070)
    );

    bfr new_Jinkela_buffer_5303 (
        .din(new_Jinkela_wire_6361),
        .dout(new_Jinkela_wire_6362)
    );

    bfr new_Jinkela_buffer_5295 (
        .din(new_Jinkela_wire_6351),
        .dout(new_Jinkela_wire_6352)
    );

    bfr new_Jinkela_buffer_8041 (
        .din(new_Jinkela_wire_10121),
        .dout(new_Jinkela_wire_10122)
    );

    bfr new_Jinkela_buffer_7998 (
        .din(new_Jinkela_wire_10070),
        .dout(new_Jinkela_wire_10071)
    );

    bfr new_Jinkela_buffer_5296 (
        .din(new_Jinkela_wire_6352),
        .dout(new_Jinkela_wire_6353)
    );

    bfr new_Jinkela_buffer_5335 (
        .din(new_Jinkela_wire_6403),
        .dout(new_Jinkela_wire_6404)
    );

    bfr new_Jinkela_buffer_7999 (
        .din(new_Jinkela_wire_10071),
        .dout(new_Jinkela_wire_10072)
    );

    bfr new_Jinkela_buffer_5304 (
        .din(new_Jinkela_wire_6362),
        .dout(new_Jinkela_wire_6363)
    );

    spl2 new_Jinkela_splitter_409 (
        .a(new_Jinkela_wire_6353),
        .b(new_Jinkela_wire_6354),
        .c(new_Jinkela_wire_6355)
    );

    bfr new_Jinkela_buffer_8192 (
        .din(new_net_6),
        .dout(new_Jinkela_wire_10294)
    );

    bfr new_Jinkela_buffer_8042 (
        .din(new_Jinkela_wire_10122),
        .dout(new_Jinkela_wire_10123)
    );

    bfr new_Jinkela_buffer_8000 (
        .din(new_Jinkela_wire_10072),
        .dout(new_Jinkela_wire_10073)
    );

    bfr new_Jinkela_buffer_5305 (
        .din(new_Jinkela_wire_6363),
        .dout(new_Jinkela_wire_6364)
    );

    bfr new_Jinkela_buffer_8063 (
        .din(new_Jinkela_wire_10157),
        .dout(new_Jinkela_wire_10158)
    );

    bfr new_Jinkela_buffer_5334 (
        .din(new_Jinkela_wire_6396),
        .dout(new_Jinkela_wire_6397)
    );

    bfr new_Jinkela_buffer_8001 (
        .din(new_Jinkela_wire_10073),
        .dout(new_Jinkela_wire_10074)
    );

    spl2 new_Jinkela_splitter_412 (
        .a(new_Jinkela_wire_6400),
        .b(new_Jinkela_wire_6401),
        .c(new_Jinkela_wire_6402)
    );

    spl4L new_Jinkela_splitter_414 (
        .a(new_Jinkela_wire_6405),
        .d(new_Jinkela_wire_6406),
        .b(new_Jinkela_wire_6407),
        .e(new_Jinkela_wire_6408),
        .c(new_Jinkela_wire_6409)
    );

    bfr new_Jinkela_buffer_8043 (
        .din(new_Jinkela_wire_10123),
        .dout(new_Jinkela_wire_10124)
    );

    bfr new_Jinkela_buffer_5306 (
        .din(new_Jinkela_wire_6364),
        .dout(new_Jinkela_wire_6365)
    );

    bfr new_Jinkela_buffer_8002 (
        .din(new_Jinkela_wire_10074),
        .dout(new_Jinkela_wire_10075)
    );

    bfr new_Jinkela_buffer_5307 (
        .din(new_Jinkela_wire_6365),
        .dout(new_Jinkela_wire_6366)
    );

    bfr new_Jinkela_buffer_8003 (
        .din(new_Jinkela_wire_10075),
        .dout(new_Jinkela_wire_10076)
    );

    bfr new_Jinkela_buffer_8126 (
        .din(new_Jinkela_wire_10220),
        .dout(new_Jinkela_wire_10221)
    );

    bfr new_Jinkela_buffer_1464 (
        .din(new_Jinkela_wire_1796),
        .dout(new_Jinkela_wire_1797)
    );

    inv n_1398_ (
        .din(new_Jinkela_wire_3271),
        .dout(n_0670_)
    );

    or_bb n_2115_ (
        .a(n_0007_),
        .b(new_Jinkela_wire_4084),
        .c(n_0008_)
    );

    bfr new_Jinkela_buffer_1400 (
        .din(new_Jinkela_wire_1732),
        .dout(new_Jinkela_wire_1733)
    );

    and_bb n_1399_ (
        .a(new_Jinkela_wire_2454),
        .b(new_Jinkela_wire_1250),
        .c(n_0671_)
    );

    and_ii n_2116_ (
        .a(new_Jinkela_wire_5370),
        .b(new_Jinkela_wire_7735),
        .c(n_0009_)
    );

    bfr new_Jinkela_buffer_1467 (
        .din(new_Jinkela_wire_1799),
        .dout(new_Jinkela_wire_1800)
    );

    and_bi n_1400_ (
        .a(new_Jinkela_wire_2889),
        .b(new_Jinkela_wire_1172),
        .c(n_0672_)
    );

    and_ii n_2117_ (
        .a(new_Jinkela_wire_5646),
        .b(new_Jinkela_wire_5926),
        .c(n_0010_)
    );

    bfr new_Jinkela_buffer_1401 (
        .din(new_Jinkela_wire_1733),
        .dout(new_Jinkela_wire_1734)
    );

    and_ii n_1401_ (
        .a(new_Jinkela_wire_4188),
        .b(new_Jinkela_wire_5927),
        .c(n_0673_)
    );

    and_ii n_2118_ (
        .a(new_Jinkela_wire_3594),
        .b(new_Jinkela_wire_6096),
        .c(n_0011_)
    );

    bfr new_Jinkela_buffer_1465 (
        .din(new_Jinkela_wire_1797),
        .dout(new_Jinkela_wire_1798)
    );

    and_bi n_1402_ (
        .a(new_Jinkela_wire_4996),
        .b(new_Jinkela_wire_9747),
        .c(n_0674_)
    );

    and_ii n_2119_ (
        .a(n_0011_),
        .b(new_Jinkela_wire_5587),
        .c(n_0012_)
    );

    bfr new_Jinkela_buffer_1402 (
        .din(new_Jinkela_wire_1734),
        .dout(new_Jinkela_wire_1735)
    );

    and_bi n_1403_ (
        .a(new_Jinkela_wire_9746),
        .b(new_Jinkela_wire_4995),
        .c(n_0675_)
    );

    and_ii n_2120_ (
        .a(new_Jinkela_wire_5163),
        .b(new_Jinkela_wire_6166),
        .c(n_0013_)
    );

    bfr new_Jinkela_buffer_1474 (
        .din(N111),
        .dout(new_Jinkela_wire_1807)
    );

    and_ii n_1404_ (
        .a(new_Jinkela_wire_9251),
        .b(new_Jinkela_wire_6768),
        .c(n_0676_)
    );

    or_bb n_2121_ (
        .a(n_0013_),
        .b(new_Jinkela_wire_9569),
        .c(n_0014_)
    );

    bfr new_Jinkela_buffer_1403 (
        .din(new_Jinkela_wire_1735),
        .dout(new_Jinkela_wire_1736)
    );

    or_ii n_1405_ (
        .a(new_Jinkela_wire_2164),
        .b(new_Jinkela_wire_1227),
        .c(n_0677_)
    );

    or_bi n_2122_ (
        .a(new_Jinkela_wire_9495),
        .b(new_Jinkela_wire_8513),
        .c(n_0015_)
    );

    bfr new_Jinkela_buffer_1468 (
        .din(new_Jinkela_wire_1800),
        .dout(new_Jinkela_wire_1801)
    );

    and_bi n_1406_ (
        .a(new_Jinkela_wire_3350),
        .b(new_Jinkela_wire_1346),
        .c(n_0678_)
    );

    and_bi n_2123_ (
        .a(new_Jinkela_wire_5363),
        .b(new_Jinkela_wire_9425),
        .c(n_0016_)
    );

    bfr new_Jinkela_buffer_1404 (
        .din(new_Jinkela_wire_1736),
        .dout(new_Jinkela_wire_1737)
    );

    and_bi n_1407_ (
        .a(new_Jinkela_wire_4520),
        .b(new_Jinkela_wire_6153),
        .c(n_0679_)
    );

    or_bi n_2124_ (
        .a(n_0016_),
        .b(new_Jinkela_wire_9913),
        .c(n_0017_)
    );

    bfr new_Jinkela_buffer_1471 (
        .din(new_Jinkela_wire_1803),
        .dout(new_Jinkela_wire_1804)
    );

    or_ii n_1408_ (
        .a(new_Jinkela_wire_7451),
        .b(new_Jinkela_wire_281),
        .c(n_0680_)
    );

    and_ii n_2125_ (
        .a(new_Jinkela_wire_8073),
        .b(new_Jinkela_wire_7681),
        .c(n_0018_)
    );

    bfr new_Jinkela_buffer_1405 (
        .din(new_Jinkela_wire_1737),
        .dout(new_Jinkela_wire_1738)
    );

    or_ii n_1409_ (
        .a(new_Jinkela_wire_1818),
        .b(new_Jinkela_wire_1203),
        .c(n_0681_)
    );

    and_ii n_2126_ (
        .a(n_0018_),
        .b(new_Jinkela_wire_6705),
        .c(n_0019_)
    );

    bfr new_Jinkela_buffer_1469 (
        .din(new_Jinkela_wire_1801),
        .dout(new_Jinkela_wire_1802)
    );

    and_bi n_1410_ (
        .a(new_Jinkela_wire_199),
        .b(new_Jinkela_wire_1325),
        .c(n_0682_)
    );

    and_bi n_2127_ (
        .a(new_Jinkela_wire_8697),
        .b(new_Jinkela_wire_8382),
        .c(n_0020_)
    );

    bfr new_Jinkela_buffer_1406 (
        .din(new_Jinkela_wire_1738),
        .dout(new_Jinkela_wire_1739)
    );

    and_bi n_1411_ (
        .a(new_Jinkela_wire_7408),
        .b(new_Jinkela_wire_7371),
        .c(n_0683_)
    );

    or_bi n_2128_ (
        .a(new_Jinkela_wire_8696),
        .b(new_Jinkela_wire_8379),
        .c(n_0021_)
    );

    bfr new_Jinkela_buffer_1478 (
        .din(N167),
        .dout(new_Jinkela_wire_1811)
    );

    or_ii n_1412_ (
        .a(new_Jinkela_wire_9024),
        .b(new_Jinkela_wire_889),
        .c(n_0684_)
    );

    and_bi n_2129_ (
        .a(new_Jinkela_wire_9498),
        .b(new_Jinkela_wire_10383),
        .c(new_net_2578)
    );

    bfr new_Jinkela_buffer_1407 (
        .din(new_Jinkela_wire_1739),
        .dout(new_Jinkela_wire_1740)
    );

    and_ii n_1413_ (
        .a(new_Jinkela_wire_9022),
        .b(new_Jinkela_wire_888),
        .c(n_0685_)
    );

    and_ii n_2130_ (
        .a(new_Jinkela_wire_4527),
        .b(new_Jinkela_wire_9458),
        .c(n_0022_)
    );

    bfr new_Jinkela_buffer_1472 (
        .din(new_Jinkela_wire_1804),
        .dout(new_Jinkela_wire_1805)
    );

    and_bi n_1414_ (
        .a(new_Jinkela_wire_6825),
        .b(new_Jinkela_wire_8755),
        .c(n_0686_)
    );

    and_bi n_2131_ (
        .a(new_Jinkela_wire_7936),
        .b(new_Jinkela_wire_2826),
        .c(n_0023_)
    );

    bfr new_Jinkela_buffer_1408 (
        .din(new_Jinkela_wire_1740),
        .dout(new_Jinkela_wire_1741)
    );

    or_ii n_1415_ (
        .a(new_Jinkela_wire_3527),
        .b(new_Jinkela_wire_1385),
        .c(n_0687_)
    );

    and_bi n_2132_ (
        .a(new_Jinkela_wire_2825),
        .b(new_Jinkela_wire_7935),
        .c(n_0024_)
    );

    bfr new_Jinkela_buffer_1475 (
        .din(new_Jinkela_wire_1807),
        .dout(new_Jinkela_wire_1808)
    );

    and_bi n_1416_ (
        .a(new_Jinkela_wire_1694),
        .b(new_Jinkela_wire_1232),
        .c(n_0688_)
    );

    and_ii n_2133_ (
        .a(new_Jinkela_wire_9584),
        .b(new_Jinkela_wire_6437),
        .c(n_0025_)
    );

    bfr new_Jinkela_buffer_1409 (
        .din(new_Jinkela_wire_1741),
        .dout(new_Jinkela_wire_1742)
    );

    or_bi n_1417_ (
        .a(new_Jinkela_wire_7850),
        .b(new_Jinkela_wire_5417),
        .c(n_0689_)
    );

    and_bi n_2134_ (
        .a(new_Jinkela_wire_3130),
        .b(new_Jinkela_wire_6941),
        .c(n_0026_)
    );

    bfr new_Jinkela_buffer_1473 (
        .din(new_Jinkela_wire_1805),
        .dout(new_Jinkela_wire_1806)
    );

    or_bb n_1421_ (
        .a(new_Jinkela_wire_8937),
        .b(new_Jinkela_wire_6103),
        .c(n_0693_)
    );

    and_bi n_2135_ (
        .a(new_Jinkela_wire_6940),
        .b(new_Jinkela_wire_3129),
        .c(n_0027_)
    );

    bfr new_Jinkela_buffer_1410 (
        .din(new_Jinkela_wire_1742),
        .dout(new_Jinkela_wire_1743)
    );

    and_bi n_1422_ (
        .a(new_Jinkela_wire_8816),
        .b(new_Jinkela_wire_8278),
        .c(n_0694_)
    );

    and_bi n_2136_ (
        .a(new_Jinkela_wire_2672),
        .b(new_Jinkela_wire_10387),
        .c(n_0028_)
    );

    bfr new_Jinkela_buffer_1482 (
        .din(N237),
        .dout(new_Jinkela_wire_1815)
    );

    or_ii n_1423_ (
        .a(new_Jinkela_wire_7994),
        .b(new_Jinkela_wire_2573),
        .c(n_0695_)
    );

    and_bi n_2137_ (
        .a(new_Jinkela_wire_10388),
        .b(new_Jinkela_wire_2671),
        .c(n_0029_)
    );

    bfr new_Jinkela_buffer_1411 (
        .din(new_Jinkela_wire_1743),
        .dout(new_Jinkela_wire_1744)
    );

    and_ii n_1424_ (
        .a(new_Jinkela_wire_7449),
        .b(new_Jinkela_wire_280),
        .c(n_0696_)
    );

    and_bi n_2138_ (
        .a(new_Jinkela_wire_1622),
        .b(new_Jinkela_wire_4966),
        .c(n_0030_)
    );

    bfr new_Jinkela_buffer_1476 (
        .din(new_Jinkela_wire_1808),
        .dout(new_Jinkela_wire_1809)
    );

    or_bb n_1425_ (
        .a(new_Jinkela_wire_4508),
        .b(new_Jinkela_wire_3924),
        .c(n_0697_)
    );

    and_bi n_2139_ (
        .a(new_Jinkela_wire_4965),
        .b(new_Jinkela_wire_1623),
        .c(n_0031_)
    );

    bfr new_Jinkela_buffer_1412 (
        .din(new_Jinkela_wire_1744),
        .dout(new_Jinkela_wire_1745)
    );

    or_bb n_1426_ (
        .a(new_Jinkela_wire_7747),
        .b(new_Jinkela_wire_8754),
        .c(n_0698_)
    );

    and_bi n_2140_ (
        .a(new_Jinkela_wire_6742),
        .b(new_Jinkela_wire_958),
        .c(n_0032_)
    );

    bfr new_Jinkela_buffer_1479 (
        .din(new_Jinkela_wire_1811),
        .dout(new_Jinkela_wire_1812)
    );

    and_bi n_1427_ (
        .a(new_Jinkela_wire_8172),
        .b(new_Jinkela_wire_8935),
        .c(n_0699_)
    );

    and_ii n_2141_ (
        .a(new_Jinkela_wire_5014),
        .b(new_Jinkela_wire_4440),
        .c(n_0033_)
    );

    bfr new_Jinkela_buffer_1413 (
        .din(new_Jinkela_wire_1745),
        .dout(new_Jinkela_wire_1746)
    );

    and_bi n_1428_ (
        .a(new_Jinkela_wire_6829),
        .b(n_0699_),
        .c(n_0700_)
    );

    and_ii n_2142_ (
        .a(new_Jinkela_wire_7300),
        .b(new_Jinkela_wire_6803),
        .c(n_0034_)
    );

    bfr new_Jinkela_buffer_1477 (
        .din(new_Jinkela_wire_1809),
        .dout(new_Jinkela_wire_1810)
    );

    and_ii n_1429_ (
        .a(new_Jinkela_wire_5561),
        .b(new_Jinkela_wire_7358),
        .c(n_0701_)
    );

    and_ii n_2143_ (
        .a(new_Jinkela_wire_5107),
        .b(new_Jinkela_wire_7771),
        .c(n_0035_)
    );

    bfr new_Jinkela_buffer_1414 (
        .din(new_Jinkela_wire_1746),
        .dout(new_Jinkela_wire_1747)
    );

    and_bb n_1430_ (
        .a(new_Jinkela_wire_7325),
        .b(new_Jinkela_wire_6316),
        .c(n_0702_)
    );

    or_bb n_2144_ (
        .a(new_Jinkela_wire_8568),
        .b(new_Jinkela_wire_10431),
        .c(n_0036_)
    );

    bfr new_Jinkela_buffer_1486 (
        .din(N112),
        .dout(new_Jinkela_wire_1819)
    );

    and_bi n_1431_ (
        .a(new_Jinkela_wire_9744),
        .b(n_0702_),
        .c(n_0703_)
    );

    and_bi n_2145_ (
        .a(new_Jinkela_wire_957),
        .b(new_Jinkela_wire_6743),
        .c(n_0037_)
    );

    bfr new_Jinkela_buffer_1415 (
        .din(new_Jinkela_wire_1747),
        .dout(new_Jinkela_wire_1748)
    );

    or_ii n_1432_ (
        .a(new_Jinkela_wire_5297),
        .b(new_Jinkela_wire_7765),
        .c(n_0704_)
    );

    and_ii n_2146_ (
        .a(new_Jinkela_wire_9160),
        .b(new_Jinkela_wire_6800),
        .c(n_0038_)
    );

    bfr new_Jinkela_buffer_1480 (
        .din(new_Jinkela_wire_1812),
        .dout(new_Jinkela_wire_1813)
    );

    and_ii n_1433_ (
        .a(new_Jinkela_wire_5296),
        .b(new_Jinkela_wire_7764),
        .c(n_0705_)
    );

    and_bb n_2147_ (
        .a(new_Jinkela_wire_7299),
        .b(new_Jinkela_wire_6824),
        .c(n_0039_)
    );

    bfr new_Jinkela_buffer_1416 (
        .din(new_Jinkela_wire_1748),
        .dout(new_Jinkela_wire_1749)
    );

    and_bi n_1434_ (
        .a(n_0704_),
        .b(n_0705_),
        .c(new_net_2568)
    );

    and_ii n_2148_ (
        .a(new_Jinkela_wire_7766),
        .b(new_Jinkela_wire_10423),
        .c(n_0040_)
    );

    bfr new_Jinkela_buffer_1483 (
        .din(new_Jinkela_wire_1815),
        .dout(new_Jinkela_wire_1816)
    );

    or_bi n_1435_ (
        .a(new_Jinkela_wire_5566),
        .b(new_Jinkela_wire_6315),
        .c(n_0706_)
    );

    inv n_2149_ (
        .din(new_Jinkela_wire_6793),
        .dout(n_0041_)
    );

    bfr new_Jinkela_buffer_1417 (
        .din(new_Jinkela_wire_1749),
        .dout(new_Jinkela_wire_1750)
    );

    or_bi n_1436_ (
        .a(new_Jinkela_wire_7352),
        .b(new_Jinkela_wire_9732),
        .c(n_0707_)
    );

    and_bi n_2150_ (
        .a(new_Jinkela_wire_6605),
        .b(new_Jinkela_wire_9847),
        .c(n_0042_)
    );

    bfr new_Jinkela_buffer_1481 (
        .din(new_Jinkela_wire_1813),
        .dout(new_Jinkela_wire_1814)
    );

    or_ii n_1437_ (
        .a(new_Jinkela_wire_9597),
        .b(new_Jinkela_wire_9571),
        .c(n_0708_)
    );

    and_bi n_2151_ (
        .a(new_Jinkela_wire_10104),
        .b(new_Jinkela_wire_7411),
        .c(n_0043_)
    );

    bfr new_Jinkela_buffer_1418 (
        .din(new_Jinkela_wire_1750),
        .dout(new_Jinkela_wire_1751)
    );

    or_bb n_1438_ (
        .a(new_Jinkela_wire_9596),
        .b(new_Jinkela_wire_9570),
        .c(n_0709_)
    );

    and_bi n_2152_ (
        .a(new_Jinkela_wire_447),
        .b(new_Jinkela_wire_5097),
        .c(n_0044_)
    );

    bfr new_Jinkela_buffer_1490 (
        .din(N113),
        .dout(new_Jinkela_wire_1823)
    );

    or_ii n_1439_ (
        .a(n_0709_),
        .b(n_0708_),
        .c(new_net_2513)
    );

    and_bi n_2153_ (
        .a(new_Jinkela_wire_5098),
        .b(new_Jinkela_wire_446),
        .c(n_0045_)
    );

    bfr new_Jinkela_buffer_1419 (
        .din(new_Jinkela_wire_1751),
        .dout(new_Jinkela_wire_1752)
    );

    and_bi n_1440_ (
        .a(new_Jinkela_wire_3925),
        .b(new_Jinkela_wire_7748),
        .c(n_0710_)
    );

    and_bi n_2154_ (
        .a(new_Jinkela_wire_2090),
        .b(new_Jinkela_wire_6253),
        .c(n_0046_)
    );

    bfr new_Jinkela_buffer_1484 (
        .din(new_Jinkela_wire_1816),
        .dout(new_Jinkela_wire_1817)
    );

    and_bi n_1441_ (
        .a(new_Jinkela_wire_4662),
        .b(new_Jinkela_wire_7930),
        .c(n_0711_)
    );

    and_bi n_2155_ (
        .a(new_Jinkela_wire_6250),
        .b(new_Jinkela_wire_2089),
        .c(n_0047_)
    );

    bfr new_Jinkela_buffer_1420 (
        .din(new_Jinkela_wire_1752),
        .dout(new_Jinkela_wire_1753)
    );

    and_ii n_1442_ (
        .a(n_0711_),
        .b(new_Jinkela_wire_4514),
        .c(n_0712_)
    );

    inv n_2156_ (
        .din(new_Jinkela_wire_3363),
        .dout(n_0048_)
    );

    bfr new_Jinkela_buffer_4430 (
        .din(new_Jinkela_wire_5269),
        .dout(new_Jinkela_wire_5270)
    );

    bfr new_Jinkela_buffer_569 (
        .din(new_Jinkela_wire_614),
        .dout(new_Jinkela_wire_615)
    );

    bfr new_Jinkela_buffer_7004 (
        .din(n_1307_),
        .dout(new_Jinkela_wire_8650)
    );

    bfr new_Jinkela_buffer_6918 (
        .din(new_Jinkela_wire_8548),
        .dout(new_Jinkela_wire_8549)
    );

    bfr new_Jinkela_buffer_509 (
        .din(new_Jinkela_wire_550),
        .dout(new_Jinkela_wire_551)
    );

    bfr new_Jinkela_buffer_4507 (
        .din(n_0825_),
        .dout(new_Jinkela_wire_5368)
    );

    bfr new_Jinkela_buffer_4431 (
        .din(new_Jinkela_wire_5270),
        .dout(new_Jinkela_wire_5271)
    );

    bfr new_Jinkela_buffer_632 (
        .din(new_Jinkela_wire_680),
        .dout(new_Jinkela_wire_681)
    );

    bfr new_Jinkela_buffer_6983 (
        .din(new_Jinkela_wire_8626),
        .dout(new_Jinkela_wire_8627)
    );

    bfr new_Jinkela_buffer_4447 (
        .din(new_Jinkela_wire_5301),
        .dout(new_Jinkela_wire_5302)
    );

    bfr new_Jinkela_buffer_510 (
        .din(new_Jinkela_wire_551),
        .dout(new_Jinkela_wire_552)
    );

    bfr new_Jinkela_buffer_6919 (
        .din(new_Jinkela_wire_8549),
        .dout(new_Jinkela_wire_8550)
    );

    bfr new_Jinkela_buffer_4432 (
        .din(new_Jinkela_wire_5271),
        .dout(new_Jinkela_wire_5272)
    );

    bfr new_Jinkela_buffer_635 (
        .din(new_Jinkela_wire_683),
        .dout(new_Jinkela_wire_684)
    );

    spl2 new_Jinkela_splitter_658 (
        .a(n_1347_),
        .b(new_Jinkela_wire_8657),
        .c(new_Jinkela_wire_8658)
    );

    bfr new_Jinkela_buffer_6940 (
        .din(new_Jinkela_wire_8580),
        .dout(new_Jinkela_wire_8581)
    );

    bfr new_Jinkela_buffer_4528 (
        .din(n_1036_),
        .dout(new_Jinkela_wire_5392)
    );

    bfr new_Jinkela_buffer_511 (
        .din(new_Jinkela_wire_552),
        .dout(new_Jinkela_wire_553)
    );

    bfr new_Jinkela_buffer_6920 (
        .din(new_Jinkela_wire_8550),
        .dout(new_Jinkela_wire_8551)
    );

    bfr new_Jinkela_buffer_4433 (
        .din(new_Jinkela_wire_5272),
        .dout(new_Jinkela_wire_5273)
    );

    bfr new_Jinkela_buffer_570 (
        .din(new_Jinkela_wire_615),
        .dout(new_Jinkela_wire_616)
    );

    bfr new_Jinkela_buffer_7009 (
        .din(new_Jinkela_wire_8658),
        .dout(new_Jinkela_wire_8659)
    );

    bfr new_Jinkela_buffer_4448 (
        .din(new_Jinkela_wire_5302),
        .dout(new_Jinkela_wire_5303)
    );

    bfr new_Jinkela_buffer_512 (
        .din(new_Jinkela_wire_553),
        .dout(new_Jinkela_wire_554)
    );

    bfr new_Jinkela_buffer_6921 (
        .din(new_Jinkela_wire_8551),
        .dout(new_Jinkela_wire_8552)
    );

    bfr new_Jinkela_buffer_4434 (
        .din(new_Jinkela_wire_5273),
        .dout(new_Jinkela_wire_5274)
    );

    bfr new_Jinkela_buffer_633 (
        .din(new_Jinkela_wire_681),
        .dout(new_Jinkela_wire_682)
    );

    spl3L new_Jinkela_splitter_659 (
        .a(n_1296_),
        .d(new_Jinkela_wire_8663),
        .b(new_Jinkela_wire_8664),
        .c(new_Jinkela_wire_8665)
    );

    bfr new_Jinkela_buffer_6941 (
        .din(new_Jinkela_wire_8581),
        .dout(new_Jinkela_wire_8582)
    );

    bfr new_Jinkela_buffer_4508 (
        .din(new_Jinkela_wire_5371),
        .dout(new_Jinkela_wire_5372)
    );

    bfr new_Jinkela_buffer_513 (
        .din(new_Jinkela_wire_554),
        .dout(new_Jinkela_wire_555)
    );

    bfr new_Jinkela_buffer_6922 (
        .din(new_Jinkela_wire_8552),
        .dout(new_Jinkela_wire_8553)
    );

    bfr new_Jinkela_buffer_4489 (
        .din(new_Jinkela_wire_5345),
        .dout(new_Jinkela_wire_5346)
    );

    bfr new_Jinkela_buffer_4435 (
        .din(new_Jinkela_wire_5274),
        .dout(new_Jinkela_wire_5275)
    );

    bfr new_Jinkela_buffer_571 (
        .din(new_Jinkela_wire_616),
        .dout(new_Jinkela_wire_617)
    );

    bfr new_Jinkela_buffer_4449 (
        .din(new_Jinkela_wire_5303),
        .dout(new_Jinkela_wire_5304)
    );

    bfr new_Jinkela_buffer_514 (
        .din(new_Jinkela_wire_555),
        .dout(new_Jinkela_wire_556)
    );

    bfr new_Jinkela_buffer_6923 (
        .din(new_Jinkela_wire_8553),
        .dout(new_Jinkela_wire_8554)
    );

    bfr new_Jinkela_buffer_4436 (
        .din(new_Jinkela_wire_5275),
        .dout(new_Jinkela_wire_5276)
    );

    spl2 new_Jinkela_splitter_21 (
        .a(N334),
        .b(new_Jinkela_wire_691),
        .c(new_Jinkela_wire_692)
    );

    bfr new_Jinkela_buffer_706 (
        .din(N118),
        .dout(new_Jinkela_wire_759)
    );

    bfr new_Jinkela_buffer_6942 (
        .din(new_Jinkela_wire_8582),
        .dout(new_Jinkela_wire_8583)
    );

    bfr new_Jinkela_buffer_6924 (
        .din(new_Jinkela_wire_8554),
        .dout(new_Jinkela_wire_8555)
    );

    bfr new_Jinkela_buffer_515 (
        .din(new_Jinkela_wire_556),
        .dout(new_Jinkela_wire_557)
    );

    spl2 new_Jinkela_splitter_326 (
        .a(n_1125_),
        .b(new_Jinkela_wire_5397),
        .c(new_Jinkela_wire_5398)
    );

    bfr new_Jinkela_buffer_4437 (
        .din(new_Jinkela_wire_5276),
        .dout(new_Jinkela_wire_5277)
    );

    spl3L new_Jinkela_splitter_20 (
        .a(new_Jinkela_wire_617),
        .d(new_Jinkela_wire_618),
        .b(new_Jinkela_wire_619),
        .c(new_Jinkela_wire_620)
    );

    bfr new_Jinkela_buffer_7005 (
        .din(new_Jinkela_wire_8650),
        .dout(new_Jinkela_wire_8651)
    );

    bfr new_Jinkela_buffer_4450 (
        .din(new_Jinkela_wire_5304),
        .dout(new_Jinkela_wire_5305)
    );

    bfr new_Jinkela_buffer_516 (
        .din(new_Jinkela_wire_557),
        .dout(new_Jinkela_wire_558)
    );

    bfr new_Jinkela_buffer_6925 (
        .din(new_Jinkela_wire_8555),
        .dout(new_Jinkela_wire_8556)
    );

    bfr new_Jinkela_buffer_6984 (
        .din(new_Jinkela_wire_8627),
        .dout(new_Jinkela_wire_8628)
    );

    bfr new_Jinkela_buffer_636 (
        .din(new_Jinkela_wire_684),
        .dout(new_Jinkela_wire_685)
    );

    bfr new_Jinkela_buffer_4490 (
        .din(new_Jinkela_wire_5346),
        .dout(new_Jinkela_wire_5347)
    );

    bfr new_Jinkela_buffer_6943 (
        .din(new_Jinkela_wire_8583),
        .dout(new_Jinkela_wire_8584)
    );

    bfr new_Jinkela_buffer_4451 (
        .din(new_Jinkela_wire_5305),
        .dout(new_Jinkela_wire_5306)
    );

    bfr new_Jinkela_buffer_517 (
        .din(new_Jinkela_wire_558),
        .dout(new_Jinkela_wire_559)
    );

    bfr new_Jinkela_buffer_6926 (
        .din(new_Jinkela_wire_8556),
        .dout(new_Jinkela_wire_8557)
    );

    bfr new_Jinkela_buffer_572 (
        .din(new_Jinkela_wire_620),
        .dout(new_Jinkela_wire_621)
    );

    spl3L new_Jinkela_splitter_324 (
        .a(n_0008_),
        .d(new_Jinkela_wire_5369),
        .b(new_Jinkela_wire_5370),
        .c(new_Jinkela_wire_5371)
    );

    bfr new_Jinkela_buffer_4452 (
        .din(new_Jinkela_wire_5306),
        .dout(new_Jinkela_wire_5307)
    );

    bfr new_Jinkela_buffer_518 (
        .din(new_Jinkela_wire_559),
        .dout(new_Jinkela_wire_560)
    );

    bfr new_Jinkela_buffer_6927 (
        .din(new_Jinkela_wire_8557),
        .dout(new_Jinkela_wire_8558)
    );

    bfr new_Jinkela_buffer_639 (
        .din(new_Jinkela_wire_687),
        .dout(new_Jinkela_wire_688)
    );

    bfr new_Jinkela_buffer_4491 (
        .din(new_Jinkela_wire_5347),
        .dout(new_Jinkela_wire_5348)
    );

    bfr new_Jinkela_buffer_6944 (
        .din(new_Jinkela_wire_8584),
        .dout(new_Jinkela_wire_8585)
    );

    bfr new_Jinkela_buffer_4453 (
        .din(new_Jinkela_wire_5307),
        .dout(new_Jinkela_wire_5308)
    );

    bfr new_Jinkela_buffer_519 (
        .din(new_Jinkela_wire_560),
        .dout(new_Jinkela_wire_561)
    );

    bfr new_Jinkela_buffer_6928 (
        .din(new_Jinkela_wire_8558),
        .dout(new_Jinkela_wire_8559)
    );

    bfr new_Jinkela_buffer_573 (
        .din(new_Jinkela_wire_621),
        .dout(new_Jinkela_wire_622)
    );

    bfr new_Jinkela_buffer_4533 (
        .din(n_0306_),
        .dout(new_Jinkela_wire_5401)
    );

    bfr new_Jinkela_buffer_4454 (
        .din(new_Jinkela_wire_5308),
        .dout(new_Jinkela_wire_5309)
    );

    bfr new_Jinkela_buffer_520 (
        .din(new_Jinkela_wire_561),
        .dout(new_Jinkela_wire_562)
    );

    bfr new_Jinkela_buffer_6929 (
        .din(new_Jinkela_wire_8559),
        .dout(new_Jinkela_wire_8560)
    );

    bfr new_Jinkela_buffer_6985 (
        .din(new_Jinkela_wire_8628),
        .dout(new_Jinkela_wire_8629)
    );

    bfr new_Jinkela_buffer_637 (
        .din(new_Jinkela_wire_685),
        .dout(new_Jinkela_wire_686)
    );

    bfr new_Jinkela_buffer_4492 (
        .din(new_Jinkela_wire_5348),
        .dout(new_Jinkela_wire_5349)
    );

    bfr new_Jinkela_buffer_6945 (
        .din(new_Jinkela_wire_8585),
        .dout(new_Jinkela_wire_8586)
    );

    bfr new_Jinkela_buffer_4455 (
        .din(new_Jinkela_wire_5309),
        .dout(new_Jinkela_wire_5310)
    );

    bfr new_Jinkela_buffer_521 (
        .din(new_Jinkela_wire_562),
        .dout(new_Jinkela_wire_563)
    );

    bfr new_Jinkela_buffer_6930 (
        .din(new_Jinkela_wire_8560),
        .dout(new_Jinkela_wire_8561)
    );

    bfr new_Jinkela_buffer_574 (
        .din(new_Jinkela_wire_622),
        .dout(new_Jinkela_wire_623)
    );

    bfr new_Jinkela_buffer_4456 (
        .din(new_Jinkela_wire_5310),
        .dout(new_Jinkela_wire_5311)
    );

    bfr new_Jinkela_buffer_522 (
        .din(new_Jinkela_wire_563),
        .dout(new_Jinkela_wire_564)
    );

    bfr new_Jinkela_buffer_6931 (
        .din(new_Jinkela_wire_8561),
        .dout(new_Jinkela_wire_8562)
    );

    bfr new_Jinkela_buffer_7006 (
        .din(new_Jinkela_wire_8651),
        .dout(new_Jinkela_wire_8652)
    );

    bfr new_Jinkela_buffer_642 (
        .din(new_Jinkela_wire_692),
        .dout(new_Jinkela_wire_693)
    );

    bfr new_Jinkela_buffer_4493 (
        .din(new_Jinkela_wire_5349),
        .dout(new_Jinkela_wire_5350)
    );

    bfr new_Jinkela_buffer_6946 (
        .din(new_Jinkela_wire_8586),
        .dout(new_Jinkela_wire_8587)
    );

    bfr new_Jinkela_buffer_4457 (
        .din(new_Jinkela_wire_5311),
        .dout(new_Jinkela_wire_5312)
    );

    bfr new_Jinkela_buffer_523 (
        .din(new_Jinkela_wire_564),
        .dout(new_Jinkela_wire_565)
    );

    bfr new_Jinkela_buffer_6932 (
        .din(new_Jinkela_wire_8562),
        .dout(new_Jinkela_wire_8563)
    );

    bfr new_Jinkela_buffer_575 (
        .din(new_Jinkela_wire_623),
        .dout(new_Jinkela_wire_624)
    );

    bfr new_Jinkela_buffer_4509 (
        .din(new_Jinkela_wire_5372),
        .dout(new_Jinkela_wire_5373)
    );

    bfr new_Jinkela_buffer_4458 (
        .din(new_Jinkela_wire_5312),
        .dout(new_Jinkela_wire_5313)
    );

    bfr new_Jinkela_buffer_524 (
        .din(new_Jinkela_wire_565),
        .dout(new_Jinkela_wire_566)
    );

    bfr new_Jinkela_buffer_6933 (
        .din(new_Jinkela_wire_8563),
        .dout(new_Jinkela_wire_8564)
    );

    bfr new_Jinkela_buffer_6986 (
        .din(new_Jinkela_wire_8629),
        .dout(new_Jinkela_wire_8630)
    );

    bfr new_Jinkela_buffer_640 (
        .din(new_Jinkela_wire_688),
        .dout(new_Jinkela_wire_689)
    );

    bfr new_Jinkela_buffer_4494 (
        .din(new_Jinkela_wire_5350),
        .dout(new_Jinkela_wire_5351)
    );

    bfr new_Jinkela_buffer_6947 (
        .din(new_Jinkela_wire_8587),
        .dout(new_Jinkela_wire_8588)
    );

    bfr new_Jinkela_buffer_4459 (
        .din(new_Jinkela_wire_5313),
        .dout(new_Jinkela_wire_5314)
    );

    bfr new_Jinkela_buffer_525 (
        .din(new_Jinkela_wire_566),
        .dout(new_Jinkela_wire_567)
    );

    bfr new_Jinkela_buffer_6934 (
        .din(new_Jinkela_wire_8564),
        .dout(new_Jinkela_wire_8565)
    );

    bfr new_Jinkela_buffer_576 (
        .din(new_Jinkela_wire_624),
        .dout(new_Jinkela_wire_625)
    );

    bfr new_Jinkela_buffer_4529 (
        .din(new_Jinkela_wire_5392),
        .dout(new_Jinkela_wire_5393)
    );

    bfr new_Jinkela_buffer_4460 (
        .din(new_Jinkela_wire_5314),
        .dout(new_Jinkela_wire_5315)
    );

    bfr new_Jinkela_buffer_526 (
        .din(new_Jinkela_wire_567),
        .dout(new_Jinkela_wire_568)
    );

    bfr new_Jinkela_buffer_6935 (
        .din(new_Jinkela_wire_8565),
        .dout(new_Jinkela_wire_8566)
    );

    bfr new_Jinkela_buffer_4495 (
        .din(new_Jinkela_wire_5351),
        .dout(new_Jinkela_wire_5352)
    );

    bfr new_Jinkela_buffer_6948 (
        .din(new_Jinkela_wire_8588),
        .dout(new_Jinkela_wire_8589)
    );

    bfr new_Jinkela_buffer_4461 (
        .din(new_Jinkela_wire_5315),
        .dout(new_Jinkela_wire_5316)
    );

    bfr new_Jinkela_buffer_527 (
        .din(new_Jinkela_wire_568),
        .dout(new_Jinkela_wire_569)
    );

    bfr new_Jinkela_buffer_6987 (
        .din(new_Jinkela_wire_8630),
        .dout(new_Jinkela_wire_8631)
    );

    bfr new_Jinkela_buffer_577 (
        .din(new_Jinkela_wire_625),
        .dout(new_Jinkela_wire_626)
    );

    bfr new_Jinkela_buffer_4510 (
        .din(new_Jinkela_wire_5373),
        .dout(new_Jinkela_wire_5374)
    );

    bfr new_Jinkela_buffer_6949 (
        .din(new_Jinkela_wire_8589),
        .dout(new_Jinkela_wire_8590)
    );

    bfr new_Jinkela_buffer_4462 (
        .din(new_Jinkela_wire_5316),
        .dout(new_Jinkela_wire_5317)
    );

    bfr new_Jinkela_buffer_528 (
        .din(new_Jinkela_wire_569),
        .dout(new_Jinkela_wire_570)
    );

    bfr new_Jinkela_buffer_7043 (
        .din(n_1293_),
        .dout(new_Jinkela_wire_8698)
    );

    bfr new_Jinkela_buffer_641 (
        .din(new_Jinkela_wire_689),
        .dout(new_Jinkela_wire_690)
    );

    bfr new_Jinkela_buffer_4496 (
        .din(new_Jinkela_wire_5352),
        .dout(new_Jinkela_wire_5353)
    );

    bfr new_Jinkela_buffer_6950 (
        .din(new_Jinkela_wire_8590),
        .dout(new_Jinkela_wire_8591)
    );

    bfr new_Jinkela_buffer_4463 (
        .din(new_Jinkela_wire_5317),
        .dout(new_Jinkela_wire_5318)
    );

    bfr new_Jinkela_buffer_529 (
        .din(new_Jinkela_wire_570),
        .dout(new_Jinkela_wire_571)
    );

    bfr new_Jinkela_buffer_7007 (
        .din(new_Jinkela_wire_8652),
        .dout(new_Jinkela_wire_8653)
    );

    bfr new_Jinkela_buffer_6275 (
        .din(new_Jinkela_wire_7652),
        .dout(new_Jinkela_wire_7653)
    );

    bfr new_Jinkela_buffer_8044 (
        .din(new_Jinkela_wire_10124),
        .dout(new_Jinkela_wire_10125)
    );

    bfr new_Jinkela_buffer_6099 (
        .din(new_Jinkela_wire_7442),
        .dout(new_Jinkela_wire_7443)
    );

    bfr new_Jinkela_buffer_8004 (
        .din(new_Jinkela_wire_10076),
        .dout(new_Jinkela_wire_10077)
    );

    bfr new_Jinkela_buffer_6112 (
        .din(new_Jinkela_wire_7473),
        .dout(new_Jinkela_wire_7474)
    );

    bfr new_Jinkela_buffer_8064 (
        .din(new_Jinkela_wire_10158),
        .dout(new_Jinkela_wire_10159)
    );

    bfr new_Jinkela_buffer_6100 (
        .din(new_Jinkela_wire_7443),
        .dout(new_Jinkela_wire_7444)
    );

    bfr new_Jinkela_buffer_8005 (
        .din(new_Jinkela_wire_10077),
        .dout(new_Jinkela_wire_10078)
    );

    bfr new_Jinkela_buffer_6212 (
        .din(new_net_10),
        .dout(new_Jinkela_wire_7586)
    );

    bfr new_Jinkela_buffer_6142 (
        .din(new_Jinkela_wire_7507),
        .dout(new_Jinkela_wire_7508)
    );

    bfr new_Jinkela_buffer_8045 (
        .din(new_Jinkela_wire_10125),
        .dout(new_Jinkela_wire_10126)
    );

    bfr new_Jinkela_buffer_6101 (
        .din(new_Jinkela_wire_7444),
        .dout(new_Jinkela_wire_7445)
    );

    bfr new_Jinkela_buffer_8006 (
        .din(new_Jinkela_wire_10078),
        .dout(new_Jinkela_wire_10079)
    );

    bfr new_Jinkela_buffer_6113 (
        .din(new_Jinkela_wire_7474),
        .dout(new_Jinkela_wire_7475)
    );

    bfr new_Jinkela_buffer_6102 (
        .din(new_Jinkela_wire_7445),
        .dout(new_Jinkela_wire_7446)
    );

    bfr new_Jinkela_buffer_8007 (
        .din(new_Jinkela_wire_10079),
        .dout(new_Jinkela_wire_10080)
    );

    spl3L new_Jinkela_splitter_841 (
        .a(new_Jinkela_wire_10222),
        .d(new_Jinkela_wire_10223),
        .b(new_Jinkela_wire_10224),
        .c(new_Jinkela_wire_10225)
    );

    bfr new_Jinkela_buffer_8046 (
        .din(new_Jinkela_wire_10126),
        .dout(new_Jinkela_wire_10127)
    );

    bfr new_Jinkela_buffer_6114 (
        .din(new_Jinkela_wire_7475),
        .dout(new_Jinkela_wire_7476)
    );

    bfr new_Jinkela_buffer_8008 (
        .din(new_Jinkela_wire_10080),
        .dout(new_Jinkela_wire_10081)
    );

    bfr new_Jinkela_buffer_6175 (
        .din(new_Jinkela_wire_7546),
        .dout(new_Jinkela_wire_7547)
    );

    bfr new_Jinkela_buffer_6143 (
        .din(new_Jinkela_wire_7508),
        .dout(new_Jinkela_wire_7509)
    );

    bfr new_Jinkela_buffer_8065 (
        .din(new_Jinkela_wire_10159),
        .dout(new_Jinkela_wire_10160)
    );

    bfr new_Jinkela_buffer_6115 (
        .din(new_Jinkela_wire_7476),
        .dout(new_Jinkela_wire_7477)
    );

    bfr new_Jinkela_buffer_8009 (
        .din(new_Jinkela_wire_10081),
        .dout(new_Jinkela_wire_10082)
    );

    spl2 new_Jinkela_splitter_542 (
        .a(n_1299_),
        .b(new_Jinkela_wire_7651),
        .c(new_Jinkela_wire_7652)
    );

    bfr new_Jinkela_buffer_8047 (
        .din(new_Jinkela_wire_10127),
        .dout(new_Jinkela_wire_10128)
    );

    bfr new_Jinkela_buffer_6116 (
        .din(new_Jinkela_wire_7477),
        .dout(new_Jinkela_wire_7478)
    );

    bfr new_Jinkela_buffer_8010 (
        .din(new_Jinkela_wire_10082),
        .dout(new_Jinkela_wire_10083)
    );

    bfr new_Jinkela_buffer_6144 (
        .din(new_Jinkela_wire_7509),
        .dout(new_Jinkela_wire_7510)
    );

    bfr new_Jinkela_buffer_6117 (
        .din(new_Jinkela_wire_7478),
        .dout(new_Jinkela_wire_7479)
    );

    bfr new_Jinkela_buffer_8011 (
        .din(new_Jinkela_wire_10083),
        .dout(new_Jinkela_wire_10084)
    );

    bfr new_Jinkela_buffer_6213 (
        .din(new_Jinkela_wire_7586),
        .dout(new_Jinkela_wire_7587)
    );

    bfr new_Jinkela_buffer_8048 (
        .din(new_Jinkela_wire_10128),
        .dout(new_Jinkela_wire_10129)
    );

    bfr new_Jinkela_buffer_6118 (
        .din(new_Jinkela_wire_7479),
        .dout(new_Jinkela_wire_7480)
    );

    bfr new_Jinkela_buffer_8012 (
        .din(new_Jinkela_wire_10084),
        .dout(new_Jinkela_wire_10085)
    );

    bfr new_Jinkela_buffer_6304 (
        .din(n_0179_),
        .dout(new_Jinkela_wire_7682)
    );

    bfr new_Jinkela_buffer_6145 (
        .din(new_Jinkela_wire_7510),
        .dout(new_Jinkela_wire_7511)
    );

    bfr new_Jinkela_buffer_8066 (
        .din(new_Jinkela_wire_10160),
        .dout(new_Jinkela_wire_10161)
    );

    bfr new_Jinkela_buffer_6119 (
        .din(new_Jinkela_wire_7480),
        .dout(new_Jinkela_wire_7481)
    );

    bfr new_Jinkela_buffer_8013 (
        .din(new_Jinkela_wire_10085),
        .dout(new_Jinkela_wire_10086)
    );

    spl2 new_Jinkela_splitter_540 (
        .a(new_Jinkela_wire_7547),
        .b(new_Jinkela_wire_7548),
        .c(new_Jinkela_wire_7549)
    );

    bfr new_Jinkela_buffer_8049 (
        .din(new_Jinkela_wire_10129),
        .dout(new_Jinkela_wire_10130)
    );

    bfr new_Jinkela_buffer_6120 (
        .din(new_Jinkela_wire_7481),
        .dout(new_Jinkela_wire_7482)
    );

    bfr new_Jinkela_buffer_8014 (
        .din(new_Jinkela_wire_10086),
        .dout(new_Jinkela_wire_10087)
    );

    bfr new_Jinkela_buffer_6146 (
        .din(new_Jinkela_wire_7511),
        .dout(new_Jinkela_wire_7512)
    );

    bfr new_Jinkela_buffer_8129 (
        .din(new_Jinkela_wire_10230),
        .dout(new_Jinkela_wire_10231)
    );

    bfr new_Jinkela_buffer_6121 (
        .din(new_Jinkela_wire_7482),
        .dout(new_Jinkela_wire_7483)
    );

    bfr new_Jinkela_buffer_8015 (
        .din(new_Jinkela_wire_10087),
        .dout(new_Jinkela_wire_10088)
    );

    bfr new_Jinkela_buffer_8237 (
        .din(n_0586_),
        .dout(new_Jinkela_wire_10341)
    );

    bfr new_Jinkela_buffer_6176 (
        .din(new_Jinkela_wire_7549),
        .dout(new_Jinkela_wire_7550)
    );

    bfr new_Jinkela_buffer_8050 (
        .din(new_Jinkela_wire_10130),
        .dout(new_Jinkela_wire_10131)
    );

    bfr new_Jinkela_buffer_6122 (
        .din(new_Jinkela_wire_7483),
        .dout(new_Jinkela_wire_7484)
    );

    bfr new_Jinkela_buffer_8016 (
        .din(new_Jinkela_wire_10088),
        .dout(new_Jinkela_wire_10089)
    );

    bfr new_Jinkela_buffer_6147 (
        .din(new_Jinkela_wire_7512),
        .dout(new_Jinkela_wire_7513)
    );

    bfr new_Jinkela_buffer_8067 (
        .din(new_Jinkela_wire_10161),
        .dout(new_Jinkela_wire_10162)
    );

    bfr new_Jinkela_buffer_6123 (
        .din(new_Jinkela_wire_7484),
        .dout(new_Jinkela_wire_7485)
    );

    bfr new_Jinkela_buffer_8017 (
        .din(new_Jinkela_wire_10089),
        .dout(new_Jinkela_wire_10090)
    );

    bfr new_Jinkela_buffer_8051 (
        .din(new_Jinkela_wire_10131),
        .dout(new_Jinkela_wire_10132)
    );

    bfr new_Jinkela_buffer_6124 (
        .din(new_Jinkela_wire_7485),
        .dout(new_Jinkela_wire_7486)
    );

    bfr new_Jinkela_buffer_8018 (
        .din(new_Jinkela_wire_10090),
        .dout(new_Jinkela_wire_10091)
    );

    bfr new_Jinkela_buffer_6148 (
        .din(new_Jinkela_wire_7513),
        .dout(new_Jinkela_wire_7514)
    );

    bfr new_Jinkela_buffer_8128 (
        .din(new_Jinkela_wire_10225),
        .dout(new_Jinkela_wire_10226)
    );

    bfr new_Jinkela_buffer_6125 (
        .din(new_Jinkela_wire_7486),
        .dout(new_Jinkela_wire_7487)
    );

    bfr new_Jinkela_buffer_8019 (
        .din(new_Jinkela_wire_10091),
        .dout(new_Jinkela_wire_10092)
    );

    bfr new_Jinkela_buffer_8052 (
        .din(new_Jinkela_wire_10132),
        .dout(new_Jinkela_wire_10133)
    );

    bfr new_Jinkela_buffer_6126 (
        .din(new_Jinkela_wire_7487),
        .dout(new_Jinkela_wire_7488)
    );

    bfr new_Jinkela_buffer_8020 (
        .din(new_Jinkela_wire_10092),
        .dout(new_Jinkela_wire_10093)
    );

    bfr new_Jinkela_buffer_6214 (
        .din(new_Jinkela_wire_7587),
        .dout(new_Jinkela_wire_7588)
    );

    bfr new_Jinkela_buffer_6149 (
        .din(new_Jinkela_wire_7514),
        .dout(new_Jinkela_wire_7515)
    );

    bfr new_Jinkela_buffer_8068 (
        .din(new_Jinkela_wire_10162),
        .dout(new_Jinkela_wire_10163)
    );

    bfr new_Jinkela_buffer_6127 (
        .din(new_Jinkela_wire_7488),
        .dout(new_Jinkela_wire_7489)
    );

    bfr new_Jinkela_buffer_8021 (
        .din(new_Jinkela_wire_10093),
        .dout(new_Jinkela_wire_10094)
    );

    bfr new_Jinkela_buffer_6177 (
        .din(new_Jinkela_wire_7550),
        .dout(new_Jinkela_wire_7551)
    );

    bfr new_Jinkela_buffer_8053 (
        .din(new_Jinkela_wire_10133),
        .dout(new_Jinkela_wire_10134)
    );

    bfr new_Jinkela_buffer_6128 (
        .din(new_Jinkela_wire_7489),
        .dout(new_Jinkela_wire_7490)
    );

    bfr new_Jinkela_buffer_8022 (
        .din(new_Jinkela_wire_10094),
        .dout(new_Jinkela_wire_10095)
    );

    bfr new_Jinkela_buffer_6150 (
        .din(new_Jinkela_wire_7515),
        .dout(new_Jinkela_wire_7516)
    );

    bfr new_Jinkela_buffer_6129 (
        .din(new_Jinkela_wire_7490),
        .dout(new_Jinkela_wire_7491)
    );

    bfr new_Jinkela_buffer_8023 (
        .din(new_Jinkela_wire_10095),
        .dout(new_Jinkela_wire_10096)
    );

    bfr new_Jinkela_buffer_8069 (
        .din(new_Jinkela_wire_10163),
        .dout(new_Jinkela_wire_10164)
    );

    bfr new_Jinkela_buffer_6130 (
        .din(new_Jinkela_wire_7491),
        .dout(new_Jinkela_wire_7492)
    );

    spl2 new_Jinkela_splitter_842 (
        .a(new_Jinkela_wire_10226),
        .b(new_Jinkela_wire_10227),
        .c(new_Jinkela_wire_10228)
    );

    bfr new_Jinkela_buffer_3633 (
        .din(new_Jinkela_wire_4247),
        .dout(new_Jinkela_wire_4248)
    );

    bfr new_Jinkela_buffer_3602 (
        .din(new_Jinkela_wire_4208),
        .dout(new_Jinkela_wire_4209)
    );

    bfr new_Jinkela_buffer_3669 (
        .din(new_Jinkela_wire_4283),
        .dout(new_Jinkela_wire_4284)
    );

    bfr new_Jinkela_buffer_3603 (
        .din(new_Jinkela_wire_4209),
        .dout(new_Jinkela_wire_4210)
    );

    bfr new_Jinkela_buffer_3634 (
        .din(new_Jinkela_wire_4248),
        .dout(new_Jinkela_wire_4249)
    );

    bfr new_Jinkela_buffer_3604 (
        .din(new_Jinkela_wire_4210),
        .dout(new_Jinkela_wire_4211)
    );

    bfr new_Jinkela_buffer_3682 (
        .din(new_Jinkela_wire_4296),
        .dout(new_Jinkela_wire_4297)
    );

    bfr new_Jinkela_buffer_3605 (
        .din(new_Jinkela_wire_4211),
        .dout(new_Jinkela_wire_4212)
    );

    bfr new_Jinkela_buffer_3635 (
        .din(new_Jinkela_wire_4249),
        .dout(new_Jinkela_wire_4250)
    );

    bfr new_Jinkela_buffer_3606 (
        .din(new_Jinkela_wire_4212),
        .dout(new_Jinkela_wire_4213)
    );

    bfr new_Jinkela_buffer_3670 (
        .din(new_Jinkela_wire_4284),
        .dout(new_Jinkela_wire_4285)
    );

    bfr new_Jinkela_buffer_3607 (
        .din(new_Jinkela_wire_4213),
        .dout(new_Jinkela_wire_4214)
    );

    bfr new_Jinkela_buffer_3636 (
        .din(new_Jinkela_wire_4250),
        .dout(new_Jinkela_wire_4251)
    );

    bfr new_Jinkela_buffer_3608 (
        .din(new_Jinkela_wire_4214),
        .dout(new_Jinkela_wire_4215)
    );

    bfr new_Jinkela_buffer_3609 (
        .din(new_Jinkela_wire_4215),
        .dout(new_Jinkela_wire_4216)
    );

    bfr new_Jinkela_buffer_3637 (
        .din(new_Jinkela_wire_4251),
        .dout(new_Jinkela_wire_4252)
    );

    bfr new_Jinkela_buffer_3610 (
        .din(new_Jinkela_wire_4216),
        .dout(new_Jinkela_wire_4217)
    );

    bfr new_Jinkela_buffer_3692 (
        .din(new_Jinkela_wire_4310),
        .dout(new_Jinkela_wire_4311)
    );

    bfr new_Jinkela_buffer_3671 (
        .din(new_Jinkela_wire_4285),
        .dout(new_Jinkela_wire_4286)
    );

    bfr new_Jinkela_buffer_3611 (
        .din(new_Jinkela_wire_4217),
        .dout(new_Jinkela_wire_4218)
    );

    bfr new_Jinkela_buffer_3638 (
        .din(new_Jinkela_wire_4252),
        .dout(new_Jinkela_wire_4253)
    );

    bfr new_Jinkela_buffer_3612 (
        .din(new_Jinkela_wire_4218),
        .dout(new_Jinkela_wire_4219)
    );

    bfr new_Jinkela_buffer_3683 (
        .din(new_Jinkela_wire_4297),
        .dout(new_Jinkela_wire_4298)
    );

    bfr new_Jinkela_buffer_3613 (
        .din(new_Jinkela_wire_4219),
        .dout(new_Jinkela_wire_4220)
    );

    bfr new_Jinkela_buffer_3639 (
        .din(new_Jinkela_wire_4253),
        .dout(new_Jinkela_wire_4254)
    );

    bfr new_Jinkela_buffer_3614 (
        .din(new_Jinkela_wire_4220),
        .dout(new_Jinkela_wire_4221)
    );

    bfr new_Jinkela_buffer_3672 (
        .din(new_Jinkela_wire_4286),
        .dout(new_Jinkela_wire_4287)
    );

    bfr new_Jinkela_buffer_3615 (
        .din(new_Jinkela_wire_4221),
        .dout(new_Jinkela_wire_4222)
    );

    bfr new_Jinkela_buffer_3640 (
        .din(new_Jinkela_wire_4254),
        .dout(new_Jinkela_wire_4255)
    );

    bfr new_Jinkela_buffer_3616 (
        .din(new_Jinkela_wire_4222),
        .dout(new_Jinkela_wire_4223)
    );

    bfr new_Jinkela_buffer_3617 (
        .din(new_Jinkela_wire_4223),
        .dout(new_Jinkela_wire_4224)
    );

    bfr new_Jinkela_buffer_3641 (
        .din(new_Jinkela_wire_4255),
        .dout(new_Jinkela_wire_4256)
    );

    bfr new_Jinkela_buffer_3618 (
        .din(new_Jinkela_wire_4224),
        .dout(new_Jinkela_wire_4225)
    );

    bfr new_Jinkela_buffer_3718 (
        .din(n_0169_),
        .dout(new_Jinkela_wire_4339)
    );

    bfr new_Jinkela_buffer_3673 (
        .din(new_Jinkela_wire_4287),
        .dout(new_Jinkela_wire_4288)
    );

    bfr new_Jinkela_buffer_3619 (
        .din(new_Jinkela_wire_4225),
        .dout(new_Jinkela_wire_4226)
    );

    bfr new_Jinkela_buffer_3642 (
        .din(new_Jinkela_wire_4256),
        .dout(new_Jinkela_wire_4257)
    );

    bfr new_Jinkela_buffer_3620 (
        .din(new_Jinkela_wire_4226),
        .dout(new_Jinkela_wire_4227)
    );

    bfr new_Jinkela_buffer_3684 (
        .din(new_Jinkela_wire_4298),
        .dout(new_Jinkela_wire_4299)
    );

    bfr new_Jinkela_buffer_3621 (
        .din(new_Jinkela_wire_4227),
        .dout(new_Jinkela_wire_4228)
    );

    bfr new_Jinkela_buffer_3643 (
        .din(new_Jinkela_wire_4257),
        .dout(new_Jinkela_wire_4258)
    );

    bfr new_Jinkela_buffer_3622 (
        .din(new_Jinkela_wire_4228),
        .dout(new_Jinkela_wire_4229)
    );

    bfr new_Jinkela_buffer_2795 (
        .din(new_Jinkela_wire_3214),
        .dout(new_Jinkela_wire_3215)
    );

    bfr new_Jinkela_buffer_2742 (
        .din(new_Jinkela_wire_3156),
        .dout(new_Jinkela_wire_3157)
    );

    bfr new_Jinkela_buffer_2854 (
        .din(new_Jinkela_wire_3277),
        .dout(new_Jinkela_wire_3278)
    );

    bfr new_Jinkela_buffer_2743 (
        .din(new_Jinkela_wire_3157),
        .dout(new_Jinkela_wire_3158)
    );

    bfr new_Jinkela_buffer_2796 (
        .din(new_Jinkela_wire_3215),
        .dout(new_Jinkela_wire_3216)
    );

    bfr new_Jinkela_buffer_2744 (
        .din(new_Jinkela_wire_3158),
        .dout(new_Jinkela_wire_3159)
    );

    bfr new_Jinkela_buffer_2918 (
        .din(new_Jinkela_wire_3341),
        .dout(new_Jinkela_wire_3342)
    );

    bfr new_Jinkela_buffer_2745 (
        .din(new_Jinkela_wire_3159),
        .dout(new_Jinkela_wire_3160)
    );

    bfr new_Jinkela_buffer_2797 (
        .din(new_Jinkela_wire_3216),
        .dout(new_Jinkela_wire_3217)
    );

    bfr new_Jinkela_buffer_2746 (
        .din(new_Jinkela_wire_3160),
        .dout(new_Jinkela_wire_3161)
    );

    bfr new_Jinkela_buffer_2855 (
        .din(new_Jinkela_wire_3278),
        .dout(new_Jinkela_wire_3279)
    );

    bfr new_Jinkela_buffer_2747 (
        .din(new_Jinkela_wire_3161),
        .dout(new_Jinkela_wire_3162)
    );

    bfr new_Jinkela_buffer_2798 (
        .din(new_Jinkela_wire_3217),
        .dout(new_Jinkela_wire_3218)
    );

    bfr new_Jinkela_buffer_2748 (
        .din(new_Jinkela_wire_3162),
        .dout(new_Jinkela_wire_3163)
    );

    bfr new_Jinkela_buffer_2927 (
        .din(N161),
        .dout(new_Jinkela_wire_3351)
    );

    bfr new_Jinkela_buffer_2749 (
        .din(new_Jinkela_wire_3163),
        .dout(new_Jinkela_wire_3164)
    );

    bfr new_Jinkela_buffer_2799 (
        .din(new_Jinkela_wire_3218),
        .dout(new_Jinkela_wire_3219)
    );

    bfr new_Jinkela_buffer_2750 (
        .din(new_Jinkela_wire_3164),
        .dout(new_Jinkela_wire_3165)
    );

    bfr new_Jinkela_buffer_2856 (
        .din(new_Jinkela_wire_3279),
        .dout(new_Jinkela_wire_3280)
    );

    bfr new_Jinkela_buffer_2751 (
        .din(new_Jinkela_wire_3165),
        .dout(new_Jinkela_wire_3166)
    );

    bfr new_Jinkela_buffer_2800 (
        .din(new_Jinkela_wire_3219),
        .dout(new_Jinkela_wire_3220)
    );

    bfr new_Jinkela_buffer_2752 (
        .din(new_Jinkela_wire_3166),
        .dout(new_Jinkela_wire_3167)
    );

    bfr new_Jinkela_buffer_2921 (
        .din(new_Jinkela_wire_3344),
        .dout(new_Jinkela_wire_3345)
    );

    bfr new_Jinkela_buffer_2753 (
        .din(new_Jinkela_wire_3167),
        .dout(new_Jinkela_wire_3168)
    );

    bfr new_Jinkela_buffer_2801 (
        .din(new_Jinkela_wire_3220),
        .dout(new_Jinkela_wire_3221)
    );

    bfr new_Jinkela_buffer_2754 (
        .din(new_Jinkela_wire_3168),
        .dout(new_Jinkela_wire_3169)
    );

    bfr new_Jinkela_buffer_2857 (
        .din(new_Jinkela_wire_3280),
        .dout(new_Jinkela_wire_3281)
    );

    bfr new_Jinkela_buffer_2755 (
        .din(new_Jinkela_wire_3169),
        .dout(new_Jinkela_wire_3170)
    );

    bfr new_Jinkela_buffer_2802 (
        .din(new_Jinkela_wire_3221),
        .dout(new_Jinkela_wire_3222)
    );

    bfr new_Jinkela_buffer_2756 (
        .din(new_Jinkela_wire_3170),
        .dout(new_Jinkela_wire_3171)
    );

    bfr new_Jinkela_buffer_2924 (
        .din(new_Jinkela_wire_3347),
        .dout(new_Jinkela_wire_3348)
    );

    bfr new_Jinkela_buffer_2757 (
        .din(new_Jinkela_wire_3171),
        .dout(new_Jinkela_wire_3172)
    );

    bfr new_Jinkela_buffer_2803 (
        .din(new_Jinkela_wire_3222),
        .dout(new_Jinkela_wire_3223)
    );

    bfr new_Jinkela_buffer_2758 (
        .din(new_Jinkela_wire_3172),
        .dout(new_Jinkela_wire_3173)
    );

    bfr new_Jinkela_buffer_2858 (
        .din(new_Jinkela_wire_3281),
        .dout(new_Jinkela_wire_3282)
    );

    bfr new_Jinkela_buffer_2759 (
        .din(new_Jinkela_wire_3173),
        .dout(new_Jinkela_wire_3174)
    );

    bfr new_Jinkela_buffer_2804 (
        .din(new_Jinkela_wire_3223),
        .dout(new_Jinkela_wire_3224)
    );

    bfr new_Jinkela_buffer_2760 (
        .din(new_Jinkela_wire_3174),
        .dout(new_Jinkela_wire_3175)
    );

    bfr new_Jinkela_buffer_2922 (
        .din(new_Jinkela_wire_3345),
        .dout(new_Jinkela_wire_3346)
    );

    bfr new_Jinkela_buffer_2761 (
        .din(new_Jinkela_wire_3175),
        .dout(new_Jinkela_wire_3176)
    );

    bfr new_Jinkela_buffer_2805 (
        .din(new_Jinkela_wire_3224),
        .dout(new_Jinkela_wire_3225)
    );

    bfr new_Jinkela_buffer_2762 (
        .din(new_Jinkela_wire_3176),
        .dout(new_Jinkela_wire_3177)
    );

    bfr new_Jinkela_buffer_1388 (
        .din(new_Jinkela_wire_1720),
        .dout(new_Jinkela_wire_1721)
    );

    bfr new_Jinkela_buffer_578 (
        .din(new_Jinkela_wire_626),
        .dout(new_Jinkela_wire_627)
    );

    bfr new_Jinkela_buffer_1338 (
        .din(new_Jinkela_wire_1663),
        .dout(new_Jinkela_wire_1664)
    );

    bfr new_Jinkela_buffer_530 (
        .din(new_Jinkela_wire_571),
        .dout(new_Jinkela_wire_572)
    );

    bfr new_Jinkela_buffer_1455 (
        .din(new_Jinkela_wire_1787),
        .dout(new_Jinkela_wire_1788)
    );

    spl2 new_Jinkela_splitter_23 (
        .a(N89),
        .b(new_Jinkela_wire_763),
        .c(new_Jinkela_wire_764)
    );

    spl2 new_Jinkela_splitter_24 (
        .a(N212),
        .b(new_Jinkela_wire_770),
        .c(new_Jinkela_wire_771)
    );

    bfr new_Jinkela_buffer_1339 (
        .din(new_Jinkela_wire_1664),
        .dout(new_Jinkela_wire_1665)
    );

    bfr new_Jinkela_buffer_531 (
        .din(new_Jinkela_wire_572),
        .dout(new_Jinkela_wire_573)
    );

    bfr new_Jinkela_buffer_1389 (
        .din(new_Jinkela_wire_1721),
        .dout(new_Jinkela_wire_1722)
    );

    bfr new_Jinkela_buffer_579 (
        .din(new_Jinkela_wire_627),
        .dout(new_Jinkela_wire_628)
    );

    bfr new_Jinkela_buffer_1340 (
        .din(new_Jinkela_wire_1665),
        .dout(new_Jinkela_wire_1666)
    );

    bfr new_Jinkela_buffer_532 (
        .din(new_Jinkela_wire_573),
        .dout(new_Jinkela_wire_574)
    );

    bfr new_Jinkela_buffer_1453 (
        .din(new_Jinkela_wire_1785),
        .dout(new_Jinkela_wire_1786)
    );

    bfr new_Jinkela_buffer_707 (
        .din(new_Jinkela_wire_759),
        .dout(new_Jinkela_wire_760)
    );

    bfr new_Jinkela_buffer_1341 (
        .din(new_Jinkela_wire_1666),
        .dout(new_Jinkela_wire_1667)
    );

    bfr new_Jinkela_buffer_533 (
        .din(new_Jinkela_wire_574),
        .dout(new_Jinkela_wire_575)
    );

    bfr new_Jinkela_buffer_1390 (
        .din(new_Jinkela_wire_1722),
        .dout(new_Jinkela_wire_1723)
    );

    bfr new_Jinkela_buffer_580 (
        .din(new_Jinkela_wire_628),
        .dout(new_Jinkela_wire_629)
    );

    bfr new_Jinkela_buffer_1342 (
        .din(new_Jinkela_wire_1667),
        .dout(new_Jinkela_wire_1668)
    );

    bfr new_Jinkela_buffer_534 (
        .din(new_Jinkela_wire_575),
        .dout(new_Jinkela_wire_576)
    );

    bfr new_Jinkela_buffer_1462 (
        .din(N197),
        .dout(new_Jinkela_wire_1795)
    );

    bfr new_Jinkela_buffer_643 (
        .din(new_Jinkela_wire_693),
        .dout(new_Jinkela_wire_694)
    );

    bfr new_Jinkela_buffer_1343 (
        .din(new_Jinkela_wire_1668),
        .dout(new_Jinkela_wire_1669)
    );

    bfr new_Jinkela_buffer_535 (
        .din(new_Jinkela_wire_576),
        .dout(new_Jinkela_wire_577)
    );

    bfr new_Jinkela_buffer_1391 (
        .din(new_Jinkela_wire_1723),
        .dout(new_Jinkela_wire_1724)
    );

    bfr new_Jinkela_buffer_581 (
        .din(new_Jinkela_wire_629),
        .dout(new_Jinkela_wire_630)
    );

    bfr new_Jinkela_buffer_1344 (
        .din(new_Jinkela_wire_1669),
        .dout(new_Jinkela_wire_1670)
    );

    bfr new_Jinkela_buffer_536 (
        .din(new_Jinkela_wire_577),
        .dout(new_Jinkela_wire_578)
    );

    bfr new_Jinkela_buffer_1456 (
        .din(new_Jinkela_wire_1788),
        .dout(new_Jinkela_wire_1789)
    );

    bfr new_Jinkela_buffer_710 (
        .din(new_Jinkela_wire_764),
        .dout(new_Jinkela_wire_765)
    );

    bfr new_Jinkela_buffer_1345 (
        .din(new_Jinkela_wire_1670),
        .dout(new_Jinkela_wire_1671)
    );

    bfr new_Jinkela_buffer_537 (
        .din(new_Jinkela_wire_578),
        .dout(new_Jinkela_wire_579)
    );

    bfr new_Jinkela_buffer_1392 (
        .din(new_Jinkela_wire_1724),
        .dout(new_Jinkela_wire_1725)
    );

    bfr new_Jinkela_buffer_582 (
        .din(new_Jinkela_wire_630),
        .dout(new_Jinkela_wire_631)
    );

    bfr new_Jinkela_buffer_1346 (
        .din(new_Jinkela_wire_1671),
        .dout(new_Jinkela_wire_1672)
    );

    bfr new_Jinkela_buffer_538 (
        .din(new_Jinkela_wire_579),
        .dout(new_Jinkela_wire_580)
    );

    bfr new_Jinkela_buffer_1459 (
        .din(new_Jinkela_wire_1791),
        .dout(new_Jinkela_wire_1792)
    );

    spl2 new_Jinkela_splitter_22 (
        .a(new_Jinkela_wire_694),
        .b(new_Jinkela_wire_695),
        .c(new_Jinkela_wire_696)
    );

    bfr new_Jinkela_buffer_1347 (
        .din(new_Jinkela_wire_1672),
        .dout(new_Jinkela_wire_1673)
    );

    bfr new_Jinkela_buffer_583 (
        .din(new_Jinkela_wire_631),
        .dout(new_Jinkela_wire_632)
    );

    bfr new_Jinkela_buffer_1393 (
        .din(new_Jinkela_wire_1725),
        .dout(new_Jinkela_wire_1726)
    );

    bfr new_Jinkela_buffer_644 (
        .din(new_Jinkela_wire_696),
        .dout(new_Jinkela_wire_697)
    );

    bfr new_Jinkela_buffer_1348 (
        .din(new_Jinkela_wire_1673),
        .dout(new_Jinkela_wire_1674)
    );

    bfr new_Jinkela_buffer_584 (
        .din(new_Jinkela_wire_632),
        .dout(new_Jinkela_wire_633)
    );

    bfr new_Jinkela_buffer_1457 (
        .din(new_Jinkela_wire_1789),
        .dout(new_Jinkela_wire_1790)
    );

    bfr new_Jinkela_buffer_708 (
        .din(new_Jinkela_wire_760),
        .dout(new_Jinkela_wire_761)
    );

    bfr new_Jinkela_buffer_1349 (
        .din(new_Jinkela_wire_1674),
        .dout(new_Jinkela_wire_1675)
    );

    bfr new_Jinkela_buffer_585 (
        .din(new_Jinkela_wire_633),
        .dout(new_Jinkela_wire_634)
    );

    bfr new_Jinkela_buffer_1394 (
        .din(new_Jinkela_wire_1726),
        .dout(new_Jinkela_wire_1727)
    );

    bfr new_Jinkela_buffer_1350 (
        .din(new_Jinkela_wire_1675),
        .dout(new_Jinkela_wire_1676)
    );

    bfr new_Jinkela_buffer_586 (
        .din(new_Jinkela_wire_634),
        .dout(new_Jinkela_wire_635)
    );

    bfr new_Jinkela_buffer_1466 (
        .din(N181),
        .dout(new_Jinkela_wire_1799)
    );

    bfr new_Jinkela_buffer_645 (
        .din(new_Jinkela_wire_697),
        .dout(new_Jinkela_wire_698)
    );

    bfr new_Jinkela_buffer_1351 (
        .din(new_Jinkela_wire_1676),
        .dout(new_Jinkela_wire_1677)
    );

    bfr new_Jinkela_buffer_587 (
        .din(new_Jinkela_wire_635),
        .dout(new_Jinkela_wire_636)
    );

    bfr new_Jinkela_buffer_1395 (
        .din(new_Jinkela_wire_1727),
        .dout(new_Jinkela_wire_1728)
    );

    bfr new_Jinkela_buffer_709 (
        .din(new_Jinkela_wire_761),
        .dout(new_Jinkela_wire_762)
    );

    bfr new_Jinkela_buffer_1352 (
        .din(new_Jinkela_wire_1677),
        .dout(new_Jinkela_wire_1678)
    );

    bfr new_Jinkela_buffer_588 (
        .din(new_Jinkela_wire_636),
        .dout(new_Jinkela_wire_637)
    );

    bfr new_Jinkela_buffer_1460 (
        .din(new_Jinkela_wire_1792),
        .dout(new_Jinkela_wire_1793)
    );

    bfr new_Jinkela_buffer_646 (
        .din(new_Jinkela_wire_698),
        .dout(new_Jinkela_wire_699)
    );

    bfr new_Jinkela_buffer_1353 (
        .din(new_Jinkela_wire_1678),
        .dout(new_Jinkela_wire_1679)
    );

    bfr new_Jinkela_buffer_589 (
        .din(new_Jinkela_wire_637),
        .dout(new_Jinkela_wire_638)
    );

    bfr new_Jinkela_buffer_1396 (
        .din(new_Jinkela_wire_1728),
        .dout(new_Jinkela_wire_1729)
    );

    bfr new_Jinkela_buffer_715 (
        .din(N168),
        .dout(new_Jinkela_wire_772)
    );

    bfr new_Jinkela_buffer_1354 (
        .din(new_Jinkela_wire_1679),
        .dout(new_Jinkela_wire_1680)
    );

    bfr new_Jinkela_buffer_590 (
        .din(new_Jinkela_wire_638),
        .dout(new_Jinkela_wire_639)
    );

    bfr new_Jinkela_buffer_1463 (
        .din(new_Jinkela_wire_1795),
        .dout(new_Jinkela_wire_1796)
    );

    bfr new_Jinkela_buffer_647 (
        .din(new_Jinkela_wire_699),
        .dout(new_Jinkela_wire_700)
    );

    bfr new_Jinkela_buffer_1355 (
        .din(new_Jinkela_wire_1680),
        .dout(new_Jinkela_wire_1681)
    );

    bfr new_Jinkela_buffer_591 (
        .din(new_Jinkela_wire_639),
        .dout(new_Jinkela_wire_640)
    );

    bfr new_Jinkela_buffer_1397 (
        .din(new_Jinkela_wire_1729),
        .dout(new_Jinkela_wire_1730)
    );

    bfr new_Jinkela_buffer_711 (
        .din(new_Jinkela_wire_765),
        .dout(new_Jinkela_wire_766)
    );

    bfr new_Jinkela_buffer_1356 (
        .din(new_Jinkela_wire_1681),
        .dout(new_Jinkela_wire_1682)
    );

    bfr new_Jinkela_buffer_592 (
        .din(new_Jinkela_wire_640),
        .dout(new_Jinkela_wire_641)
    );

    bfr new_Jinkela_buffer_1461 (
        .din(new_Jinkela_wire_1793),
        .dout(new_Jinkela_wire_1794)
    );

    bfr new_Jinkela_buffer_648 (
        .din(new_Jinkela_wire_700),
        .dout(new_Jinkela_wire_701)
    );

    bfr new_Jinkela_buffer_1398 (
        .din(new_Jinkela_wire_1730),
        .dout(new_Jinkela_wire_1731)
    );

    bfr new_Jinkela_buffer_593 (
        .din(new_Jinkela_wire_641),
        .dout(new_Jinkela_wire_642)
    );

    bfr new_Jinkela_buffer_1470 (
        .din(N196),
        .dout(new_Jinkela_wire_1803)
    );

    bfr new_Jinkela_buffer_719 (
        .din(N205),
        .dout(new_Jinkela_wire_776)
    );

    bfr new_Jinkela_buffer_1399 (
        .din(new_Jinkela_wire_1731),
        .dout(new_Jinkela_wire_1732)
    );

    bfr new_Jinkela_buffer_594 (
        .din(new_Jinkela_wire_642),
        .dout(new_Jinkela_wire_643)
    );

    bfr new_Jinkela_buffer_5308 (
        .din(new_Jinkela_wire_6366),
        .dout(new_Jinkela_wire_6367)
    );

    spl2 new_Jinkela_splitter_415 (
        .a(n_1190_),
        .b(new_Jinkela_wire_6429),
        .c(new_Jinkela_wire_6430)
    );

    bfr new_Jinkela_buffer_5309 (
        .din(new_Jinkela_wire_6367),
        .dout(new_Jinkela_wire_6368)
    );

    bfr new_Jinkela_buffer_5355 (
        .din(n_0213_),
        .dout(new_Jinkela_wire_6431)
    );

    bfr new_Jinkela_buffer_5336 (
        .din(new_Jinkela_wire_6409),
        .dout(new_Jinkela_wire_6410)
    );

    bfr new_Jinkela_buffer_5310 (
        .din(new_Jinkela_wire_6368),
        .dout(new_Jinkela_wire_6369)
    );

    bfr new_Jinkela_buffer_5405 (
        .din(new_net_2576),
        .dout(new_Jinkela_wire_6485)
    );

    bfr new_Jinkela_buffer_5356 (
        .din(new_Jinkela_wire_6431),
        .dout(new_Jinkela_wire_6432)
    );

    bfr new_Jinkela_buffer_5311 (
        .din(new_Jinkela_wire_6369),
        .dout(new_Jinkela_wire_6370)
    );

    bfr new_Jinkela_buffer_5312 (
        .din(new_Jinkela_wire_6370),
        .dout(new_Jinkela_wire_6371)
    );

    bfr new_Jinkela_buffer_5337 (
        .din(new_Jinkela_wire_6410),
        .dout(new_Jinkela_wire_6411)
    );

    bfr new_Jinkela_buffer_5313 (
        .din(new_Jinkela_wire_6371),
        .dout(new_Jinkela_wire_6372)
    );

    spl4L new_Jinkela_splitter_416 (
        .a(n_0023_),
        .d(new_Jinkela_wire_6435),
        .b(new_Jinkela_wire_6436),
        .e(new_Jinkela_wire_6437),
        .c(new_Jinkela_wire_6438)
    );

    bfr new_Jinkela_buffer_5314 (
        .din(new_Jinkela_wire_6372),
        .dout(new_Jinkela_wire_6373)
    );

    bfr new_Jinkela_buffer_5338 (
        .din(new_Jinkela_wire_6411),
        .dout(new_Jinkela_wire_6412)
    );

    bfr new_Jinkela_buffer_5315 (
        .din(new_Jinkela_wire_6373),
        .dout(new_Jinkela_wire_6374)
    );

    bfr new_Jinkela_buffer_5359 (
        .din(new_Jinkela_wire_6438),
        .dout(new_Jinkela_wire_6439)
    );

    bfr new_Jinkela_buffer_5316 (
        .din(new_Jinkela_wire_6374),
        .dout(new_Jinkela_wire_6375)
    );

    bfr new_Jinkela_buffer_5339 (
        .din(new_Jinkela_wire_6412),
        .dout(new_Jinkela_wire_6413)
    );

    bfr new_Jinkela_buffer_5317 (
        .din(new_Jinkela_wire_6375),
        .dout(new_Jinkela_wire_6376)
    );

    bfr new_Jinkela_buffer_5357 (
        .din(new_Jinkela_wire_6432),
        .dout(new_Jinkela_wire_6433)
    );

    bfr new_Jinkela_buffer_5318 (
        .din(new_Jinkela_wire_6376),
        .dout(new_Jinkela_wire_6377)
    );

    bfr new_Jinkela_buffer_5340 (
        .din(new_Jinkela_wire_6413),
        .dout(new_Jinkela_wire_6414)
    );

    bfr new_Jinkela_buffer_5319 (
        .din(new_Jinkela_wire_6377),
        .dout(new_Jinkela_wire_6378)
    );

    bfr new_Jinkela_buffer_5406 (
        .din(new_Jinkela_wire_6485),
        .dout(new_Jinkela_wire_6486)
    );

    bfr new_Jinkela_buffer_5320 (
        .din(new_Jinkela_wire_6378),
        .dout(new_Jinkela_wire_6379)
    );

    bfr new_Jinkela_buffer_5341 (
        .din(new_Jinkela_wire_6414),
        .dout(new_Jinkela_wire_6415)
    );

    bfr new_Jinkela_buffer_5321 (
        .din(new_Jinkela_wire_6379),
        .dout(new_Jinkela_wire_6380)
    );

    bfr new_Jinkela_buffer_5358 (
        .din(new_Jinkela_wire_6433),
        .dout(new_Jinkela_wire_6434)
    );

    bfr new_Jinkela_buffer_5322 (
        .din(new_Jinkela_wire_6380),
        .dout(new_Jinkela_wire_6381)
    );

    bfr new_Jinkela_buffer_5342 (
        .din(new_Jinkela_wire_6415),
        .dout(new_Jinkela_wire_6416)
    );

    bfr new_Jinkela_buffer_5323 (
        .din(new_Jinkela_wire_6381),
        .dout(new_Jinkela_wire_6382)
    );

    spl2 new_Jinkela_splitter_417 (
        .a(n_0957_),
        .b(new_Jinkela_wire_6513),
        .c(new_Jinkela_wire_6514)
    );

    bfr new_Jinkela_buffer_5324 (
        .din(new_Jinkela_wire_6382),
        .dout(new_Jinkela_wire_6383)
    );

    bfr new_Jinkela_buffer_5343 (
        .din(new_Jinkela_wire_6416),
        .dout(new_Jinkela_wire_6417)
    );

    bfr new_Jinkela_buffer_5325 (
        .din(new_Jinkela_wire_6383),
        .dout(new_Jinkela_wire_6384)
    );

    spl2 new_Jinkela_splitter_418 (
        .a(n_0736_),
        .b(new_Jinkela_wire_6515),
        .c(new_Jinkela_wire_6516)
    );

    bfr new_Jinkela_buffer_5360 (
        .din(new_Jinkela_wire_6439),
        .dout(new_Jinkela_wire_6440)
    );

    bfr new_Jinkela_buffer_5326 (
        .din(new_Jinkela_wire_6384),
        .dout(new_Jinkela_wire_6385)
    );

    bfr new_Jinkela_buffer_5344 (
        .din(new_Jinkela_wire_6417),
        .dout(new_Jinkela_wire_6418)
    );

    bfr new_Jinkela_buffer_5327 (
        .din(new_Jinkela_wire_6385),
        .dout(new_Jinkela_wire_6386)
    );

    bfr new_Jinkela_buffer_5328 (
        .din(new_Jinkela_wire_6386),
        .dout(new_Jinkela_wire_6387)
    );

    bfr new_Jinkela_buffer_5345 (
        .din(new_Jinkela_wire_6418),
        .dout(new_Jinkela_wire_6419)
    );

    bfr new_Jinkela_buffer_6988 (
        .din(new_Jinkela_wire_8631),
        .dout(new_Jinkela_wire_8632)
    );

    bfr new_Jinkela_buffer_4531 (
        .din(new_Jinkela_wire_5398),
        .dout(new_Jinkela_wire_5399)
    );

    bfr new_Jinkela_buffer_6951 (
        .din(new_Jinkela_wire_8591),
        .dout(new_Jinkela_wire_8592)
    );

    bfr new_Jinkela_buffer_4464 (
        .din(new_Jinkela_wire_5318),
        .dout(new_Jinkela_wire_5319)
    );

    bfr new_Jinkela_buffer_3674 (
        .din(new_Jinkela_wire_4288),
        .dout(new_Jinkela_wire_4289)
    );

    bfr new_Jinkela_buffer_3623 (
        .din(new_Jinkela_wire_4229),
        .dout(new_Jinkela_wire_4230)
    );

    bfr new_Jinkela_buffer_3644 (
        .din(new_Jinkela_wire_4258),
        .dout(new_Jinkela_wire_4259)
    );

    bfr new_Jinkela_buffer_4497 (
        .din(new_Jinkela_wire_5353),
        .dout(new_Jinkela_wire_5354)
    );

    bfr new_Jinkela_buffer_6952 (
        .din(new_Jinkela_wire_8592),
        .dout(new_Jinkela_wire_8593)
    );

    bfr new_Jinkela_buffer_4465 (
        .din(new_Jinkela_wire_5319),
        .dout(new_Jinkela_wire_5320)
    );

    bfr new_Jinkela_buffer_3624 (
        .din(new_Jinkela_wire_4230),
        .dout(new_Jinkela_wire_4231)
    );

    bfr new_Jinkela_buffer_6989 (
        .din(new_Jinkela_wire_8632),
        .dout(new_Jinkela_wire_8633)
    );

    bfr new_Jinkela_buffer_4511 (
        .din(new_Jinkela_wire_5374),
        .dout(new_Jinkela_wire_5375)
    );

    bfr new_Jinkela_buffer_6953 (
        .din(new_Jinkela_wire_8593),
        .dout(new_Jinkela_wire_8594)
    );

    bfr new_Jinkela_buffer_4466 (
        .din(new_Jinkela_wire_5320),
        .dout(new_Jinkela_wire_5321)
    );

    bfr new_Jinkela_buffer_3788 (
        .din(n_0136_),
        .dout(new_Jinkela_wire_4411)
    );

    bfr new_Jinkela_buffer_3625 (
        .din(new_Jinkela_wire_4231),
        .dout(new_Jinkela_wire_4232)
    );

    bfr new_Jinkela_buffer_3645 (
        .din(new_Jinkela_wire_4259),
        .dout(new_Jinkela_wire_4260)
    );

    bfr new_Jinkela_buffer_4498 (
        .din(new_Jinkela_wire_5354),
        .dout(new_Jinkela_wire_5355)
    );

    bfr new_Jinkela_buffer_6954 (
        .din(new_Jinkela_wire_8594),
        .dout(new_Jinkela_wire_8595)
    );

    bfr new_Jinkela_buffer_7013 (
        .din(new_Jinkela_wire_8665),
        .dout(new_Jinkela_wire_8666)
    );

    bfr new_Jinkela_buffer_4467 (
        .din(new_Jinkela_wire_5321),
        .dout(new_Jinkela_wire_5322)
    );

    bfr new_Jinkela_buffer_7008 (
        .din(new_Jinkela_wire_8653),
        .dout(new_Jinkela_wire_8654)
    );

    bfr new_Jinkela_buffer_3675 (
        .din(new_Jinkela_wire_4289),
        .dout(new_Jinkela_wire_4290)
    );

    bfr new_Jinkela_buffer_3646 (
        .din(new_Jinkela_wire_4260),
        .dout(new_Jinkela_wire_4261)
    );

    bfr new_Jinkela_buffer_4530 (
        .din(new_Jinkela_wire_5393),
        .dout(new_Jinkela_wire_5394)
    );

    bfr new_Jinkela_buffer_6955 (
        .din(new_Jinkela_wire_8595),
        .dout(new_Jinkela_wire_8596)
    );

    bfr new_Jinkela_buffer_6990 (
        .din(new_Jinkela_wire_8633),
        .dout(new_Jinkela_wire_8634)
    );

    bfr new_Jinkela_buffer_4468 (
        .din(new_Jinkela_wire_5322),
        .dout(new_Jinkela_wire_5323)
    );

    bfr new_Jinkela_buffer_3685 (
        .din(new_Jinkela_wire_4299),
        .dout(new_Jinkela_wire_4300)
    );

    bfr new_Jinkela_buffer_3647 (
        .din(new_Jinkela_wire_4261),
        .dout(new_Jinkela_wire_4262)
    );

    bfr new_Jinkela_buffer_4499 (
        .din(new_Jinkela_wire_5355),
        .dout(new_Jinkela_wire_5356)
    );

    bfr new_Jinkela_buffer_6956 (
        .din(new_Jinkela_wire_8596),
        .dout(new_Jinkela_wire_8597)
    );

    bfr new_Jinkela_buffer_4469 (
        .din(new_Jinkela_wire_5323),
        .dout(new_Jinkela_wire_5324)
    );

    bfr new_Jinkela_buffer_7010 (
        .din(new_Jinkela_wire_8659),
        .dout(new_Jinkela_wire_8660)
    );

    bfr new_Jinkela_buffer_3676 (
        .din(new_Jinkela_wire_4290),
        .dout(new_Jinkela_wire_4291)
    );

    bfr new_Jinkela_buffer_3648 (
        .din(new_Jinkela_wire_4262),
        .dout(new_Jinkela_wire_4263)
    );

    bfr new_Jinkela_buffer_4512 (
        .din(new_Jinkela_wire_5375),
        .dout(new_Jinkela_wire_5376)
    );

    bfr new_Jinkela_buffer_6957 (
        .din(new_Jinkela_wire_8597),
        .dout(new_Jinkela_wire_8598)
    );

    bfr new_Jinkela_buffer_6991 (
        .din(new_Jinkela_wire_8634),
        .dout(new_Jinkela_wire_8635)
    );

    bfr new_Jinkela_buffer_4470 (
        .din(new_Jinkela_wire_5324),
        .dout(new_Jinkela_wire_5325)
    );

    bfr new_Jinkela_buffer_3649 (
        .din(new_Jinkela_wire_4263),
        .dout(new_Jinkela_wire_4264)
    );

    bfr new_Jinkela_buffer_4500 (
        .din(new_Jinkela_wire_5356),
        .dout(new_Jinkela_wire_5357)
    );

    bfr new_Jinkela_buffer_6958 (
        .din(new_Jinkela_wire_8598),
        .dout(new_Jinkela_wire_8599)
    );

    bfr new_Jinkela_buffer_4471 (
        .din(new_Jinkela_wire_5325),
        .dout(new_Jinkela_wire_5326)
    );

    bfr new_Jinkela_buffer_3693 (
        .din(new_Jinkela_wire_4311),
        .dout(new_Jinkela_wire_4312)
    );

    spl2 new_Jinkela_splitter_657 (
        .a(new_Jinkela_wire_8654),
        .b(new_Jinkela_wire_8655),
        .c(new_Jinkela_wire_8656)
    );

    bfr new_Jinkela_buffer_6992 (
        .din(new_Jinkela_wire_8635),
        .dout(new_Jinkela_wire_8636)
    );

    bfr new_Jinkela_buffer_3677 (
        .din(new_Jinkela_wire_4291),
        .dout(new_Jinkela_wire_4292)
    );

    bfr new_Jinkela_buffer_3650 (
        .din(new_Jinkela_wire_4264),
        .dout(new_Jinkela_wire_4265)
    );

    bfr new_Jinkela_buffer_6959 (
        .din(new_Jinkela_wire_8599),
        .dout(new_Jinkela_wire_8600)
    );

    bfr new_Jinkela_buffer_4472 (
        .din(new_Jinkela_wire_5326),
        .dout(new_Jinkela_wire_5327)
    );

    bfr new_Jinkela_buffer_4544 (
        .din(n_0494_),
        .dout(new_Jinkela_wire_5412)
    );

    bfr new_Jinkela_buffer_3686 (
        .din(new_Jinkela_wire_4300),
        .dout(new_Jinkela_wire_4301)
    );

    bfr new_Jinkela_buffer_3651 (
        .din(new_Jinkela_wire_4265),
        .dout(new_Jinkela_wire_4266)
    );

    bfr new_Jinkela_buffer_4501 (
        .din(new_Jinkela_wire_5357),
        .dout(new_Jinkela_wire_5358)
    );

    bfr new_Jinkela_buffer_6960 (
        .din(new_Jinkela_wire_8600),
        .dout(new_Jinkela_wire_8601)
    );

    bfr new_Jinkela_buffer_4473 (
        .din(new_Jinkela_wire_5327),
        .dout(new_Jinkela_wire_5328)
    );

    bfr new_Jinkela_buffer_7011 (
        .din(new_Jinkela_wire_8660),
        .dout(new_Jinkela_wire_8661)
    );

    bfr new_Jinkela_buffer_3678 (
        .din(new_Jinkela_wire_4292),
        .dout(new_Jinkela_wire_4293)
    );

    bfr new_Jinkela_buffer_3652 (
        .din(new_Jinkela_wire_4266),
        .dout(new_Jinkela_wire_4267)
    );

    bfr new_Jinkela_buffer_4513 (
        .din(new_Jinkela_wire_5376),
        .dout(new_Jinkela_wire_5377)
    );

    bfr new_Jinkela_buffer_6961 (
        .din(new_Jinkela_wire_8601),
        .dout(new_Jinkela_wire_8602)
    );

    bfr new_Jinkela_buffer_6993 (
        .din(new_Jinkela_wire_8636),
        .dout(new_Jinkela_wire_8637)
    );

    bfr new_Jinkela_buffer_4474 (
        .din(new_Jinkela_wire_5328),
        .dout(new_Jinkela_wire_5329)
    );

    bfr new_Jinkela_buffer_3653 (
        .din(new_Jinkela_wire_4267),
        .dout(new_Jinkela_wire_4268)
    );

    bfr new_Jinkela_buffer_4502 (
        .din(new_Jinkela_wire_5358),
        .dout(new_Jinkela_wire_5359)
    );

    bfr new_Jinkela_buffer_6962 (
        .din(new_Jinkela_wire_8602),
        .dout(new_Jinkela_wire_8603)
    );

    bfr new_Jinkela_buffer_4475 (
        .din(new_Jinkela_wire_5329),
        .dout(new_Jinkela_wire_5330)
    );

    bfr new_Jinkela_buffer_3771 (
        .din(new_net_2549),
        .dout(new_Jinkela_wire_4394)
    );

    spl2 new_Jinkela_splitter_663 (
        .a(n_1309_),
        .b(new_Jinkela_wire_8707),
        .c(new_Jinkela_wire_8708)
    );

    bfr new_Jinkela_buffer_3679 (
        .din(new_Jinkela_wire_4293),
        .dout(new_Jinkela_wire_4294)
    );

    bfr new_Jinkela_buffer_3654 (
        .din(new_Jinkela_wire_4268),
        .dout(new_Jinkela_wire_4269)
    );

    spl2 new_Jinkela_splitter_325 (
        .a(new_Jinkela_wire_5394),
        .b(new_Jinkela_wire_5395),
        .c(new_Jinkela_wire_5396)
    );

    bfr new_Jinkela_buffer_6963 (
        .din(new_Jinkela_wire_8603),
        .dout(new_Jinkela_wire_8604)
    );

    bfr new_Jinkela_buffer_6994 (
        .din(new_Jinkela_wire_8637),
        .dout(new_Jinkela_wire_8638)
    );

    bfr new_Jinkela_buffer_4476 (
        .din(new_Jinkela_wire_5330),
        .dout(new_Jinkela_wire_5331)
    );

    bfr new_Jinkela_buffer_3687 (
        .din(new_Jinkela_wire_4301),
        .dout(new_Jinkela_wire_4302)
    );

    bfr new_Jinkela_buffer_3655 (
        .din(new_Jinkela_wire_4269),
        .dout(new_Jinkela_wire_4270)
    );

    bfr new_Jinkela_buffer_4503 (
        .din(new_Jinkela_wire_5359),
        .dout(new_Jinkela_wire_5360)
    );

    bfr new_Jinkela_buffer_6964 (
        .din(new_Jinkela_wire_8604),
        .dout(new_Jinkela_wire_8605)
    );

    bfr new_Jinkela_buffer_4477 (
        .din(new_Jinkela_wire_5331),
        .dout(new_Jinkela_wire_5332)
    );

    spl2 new_Jinkela_splitter_662 (
        .a(n_0243_),
        .b(new_Jinkela_wire_8705),
        .c(new_Jinkela_wire_8706)
    );

    bfr new_Jinkela_buffer_3680 (
        .din(new_Jinkela_wire_4294),
        .dout(new_Jinkela_wire_4295)
    );

    bfr new_Jinkela_buffer_3656 (
        .din(new_Jinkela_wire_4270),
        .dout(new_Jinkela_wire_4271)
    );

    bfr new_Jinkela_buffer_4514 (
        .din(new_Jinkela_wire_5377),
        .dout(new_Jinkela_wire_5378)
    );

    bfr new_Jinkela_buffer_6965 (
        .din(new_Jinkela_wire_8605),
        .dout(new_Jinkela_wire_8606)
    );

    bfr new_Jinkela_buffer_6995 (
        .din(new_Jinkela_wire_8638),
        .dout(new_Jinkela_wire_8639)
    );

    bfr new_Jinkela_buffer_4478 (
        .din(new_Jinkela_wire_5332),
        .dout(new_Jinkela_wire_5333)
    );

    bfr new_Jinkela_buffer_3657 (
        .din(new_Jinkela_wire_4271),
        .dout(new_Jinkela_wire_4272)
    );

    bfr new_Jinkela_buffer_4504 (
        .din(new_Jinkela_wire_5360),
        .dout(new_Jinkela_wire_5361)
    );

    bfr new_Jinkela_buffer_6966 (
        .din(new_Jinkela_wire_8606),
        .dout(new_Jinkela_wire_8607)
    );

    bfr new_Jinkela_buffer_4479 (
        .din(new_Jinkela_wire_5333),
        .dout(new_Jinkela_wire_5334)
    );

    bfr new_Jinkela_buffer_3694 (
        .din(new_Jinkela_wire_4312),
        .dout(new_Jinkela_wire_4313)
    );

    bfr new_Jinkela_buffer_7012 (
        .din(new_Jinkela_wire_8661),
        .dout(new_Jinkela_wire_8662)
    );

    bfr new_Jinkela_buffer_3688 (
        .din(new_Jinkela_wire_4302),
        .dout(new_Jinkela_wire_4303)
    );

    bfr new_Jinkela_buffer_3658 (
        .din(new_Jinkela_wire_4272),
        .dout(new_Jinkela_wire_4273)
    );

    bfr new_Jinkela_buffer_4534 (
        .din(new_Jinkela_wire_5401),
        .dout(new_Jinkela_wire_5402)
    );

    bfr new_Jinkela_buffer_6967 (
        .din(new_Jinkela_wire_8607),
        .dout(new_Jinkela_wire_8608)
    );

    bfr new_Jinkela_buffer_6996 (
        .din(new_Jinkela_wire_8639),
        .dout(new_Jinkela_wire_8640)
    );

    bfr new_Jinkela_buffer_4480 (
        .din(new_Jinkela_wire_5334),
        .dout(new_Jinkela_wire_5335)
    );

    bfr new_Jinkela_buffer_4532 (
        .din(new_Jinkela_wire_5399),
        .dout(new_Jinkela_wire_5400)
    );

    bfr new_Jinkela_buffer_3659 (
        .din(new_Jinkela_wire_4273),
        .dout(new_Jinkela_wire_4274)
    );

    bfr new_Jinkela_buffer_4505 (
        .din(new_Jinkela_wire_5361),
        .dout(new_Jinkela_wire_5362)
    );

    bfr new_Jinkela_buffer_6968 (
        .din(new_Jinkela_wire_8608),
        .dout(new_Jinkela_wire_8609)
    );

    bfr new_Jinkela_buffer_4481 (
        .din(new_Jinkela_wire_5335),
        .dout(new_Jinkela_wire_5336)
    );

    bfr new_Jinkela_buffer_3719 (
        .din(new_Jinkela_wire_4339),
        .dout(new_Jinkela_wire_4340)
    );

    bfr new_Jinkela_buffer_7044 (
        .din(new_Jinkela_wire_8698),
        .dout(new_Jinkela_wire_8699)
    );

    bfr new_Jinkela_buffer_3689 (
        .din(new_Jinkela_wire_4303),
        .dout(new_Jinkela_wire_4304)
    );

    bfr new_Jinkela_buffer_3660 (
        .din(new_Jinkela_wire_4274),
        .dout(new_Jinkela_wire_4275)
    );

    bfr new_Jinkela_buffer_4515 (
        .din(new_Jinkela_wire_5378),
        .dout(new_Jinkela_wire_5379)
    );

    bfr new_Jinkela_buffer_6969 (
        .din(new_Jinkela_wire_8609),
        .dout(new_Jinkela_wire_8610)
    );

    bfr new_Jinkela_buffer_6997 (
        .din(new_Jinkela_wire_8640),
        .dout(new_Jinkela_wire_8641)
    );

    bfr new_Jinkela_buffer_4482 (
        .din(new_Jinkela_wire_5336),
        .dout(new_Jinkela_wire_5337)
    );

    bfr new_Jinkela_buffer_3661 (
        .din(new_Jinkela_wire_4275),
        .dout(new_Jinkela_wire_4276)
    );

    bfr new_Jinkela_buffer_4506 (
        .din(new_Jinkela_wire_5362),
        .dout(new_Jinkela_wire_5363)
    );

    bfr new_Jinkela_buffer_6970 (
        .din(new_Jinkela_wire_8610),
        .dout(new_Jinkela_wire_8611)
    );

    bfr new_Jinkela_buffer_4483 (
        .din(new_Jinkela_wire_5337),
        .dout(new_Jinkela_wire_5338)
    );

    bfr new_Jinkela_buffer_3695 (
        .din(new_Jinkela_wire_4313),
        .dout(new_Jinkela_wire_4314)
    );

    bfr new_Jinkela_buffer_6998 (
        .din(new_Jinkela_wire_8641),
        .dout(new_Jinkela_wire_8642)
    );

    bfr new_Jinkela_buffer_3690 (
        .din(new_Jinkela_wire_4304),
        .dout(new_Jinkela_wire_4305)
    );

    bfr new_Jinkela_buffer_4547 (
        .din(n_0687_),
        .dout(new_Jinkela_wire_5417)
    );

    bfr new_Jinkela_buffer_6971 (
        .din(new_Jinkela_wire_8611),
        .dout(new_Jinkela_wire_8612)
    );

    bfr new_Jinkela_buffer_4484 (
        .din(new_Jinkela_wire_5338),
        .dout(new_Jinkela_wire_5339)
    );

    bfr new_Jinkela_buffer_6151 (
        .din(new_Jinkela_wire_7516),
        .dout(new_Jinkela_wire_7517)
    );

    bfr new_Jinkela_buffer_2859 (
        .din(new_Jinkela_wire_3282),
        .dout(new_Jinkela_wire_3283)
    );

    bfr new_Jinkela_buffer_8070 (
        .din(new_Jinkela_wire_10164),
        .dout(new_Jinkela_wire_10165)
    );

    and_bi n_1443_ (
        .a(new_Jinkela_wire_6529),
        .b(new_Jinkela_wire_8818),
        .c(n_0713_)
    );

    and_bi n_2157_ (
        .a(new_Jinkela_wire_9920),
        .b(new_Jinkela_wire_3862),
        .c(n_0049_)
    );

    bfr new_Jinkela_buffer_6131 (
        .din(new_Jinkela_wire_7492),
        .dout(new_Jinkela_wire_7493)
    );

    bfr new_Jinkela_buffer_2763 (
        .din(new_Jinkela_wire_3177),
        .dout(new_Jinkela_wire_3178)
    );

    and_bi n_1444_ (
        .a(new_Jinkela_wire_8819),
        .b(new_Jinkela_wire_6528),
        .c(n_0714_)
    );

    inv n_2158_ (
        .din(new_Jinkela_wire_5644),
        .dout(n_0050_)
    );

    bfr new_Jinkela_buffer_6178 (
        .din(new_Jinkela_wire_7551),
        .dout(new_Jinkela_wire_7552)
    );

    bfr new_Jinkela_buffer_2806 (
        .din(new_Jinkela_wire_3225),
        .dout(new_Jinkela_wire_3226)
    );

    bfr new_Jinkela_buffer_8071 (
        .din(new_Jinkela_wire_10165),
        .dout(new_Jinkela_wire_10166)
    );

    or_bb n_1445_ (
        .a(n_0714_),
        .b(n_0713_),
        .c(new_net_2558)
    );

    and_bi n_2159_ (
        .a(new_Jinkela_wire_3865),
        .b(new_Jinkela_wire_9919),
        .c(n_0051_)
    );

    bfr new_Jinkela_buffer_6132 (
        .din(new_Jinkela_wire_7493),
        .dout(new_Jinkela_wire_7494)
    );

    spl2 new_Jinkela_splitter_844 (
        .a(new_Jinkela_wire_10294),
        .b(new_Jinkela_wire_10295),
        .c(new_Jinkela_wire_10296)
    );

    bfr new_Jinkela_buffer_2764 (
        .din(new_Jinkela_wire_3178),
        .dout(new_Jinkela_wire_3179)
    );

    and_bi n_1446_ (
        .a(new_Jinkela_wire_3928),
        .b(new_Jinkela_wire_7929),
        .c(n_0715_)
    );

    and_ii n_2160_ (
        .a(new_Jinkela_wire_5157),
        .b(new_Jinkela_wire_1412),
        .c(n_0052_)
    );

    bfr new_Jinkela_buffer_8238 (
        .din(n_1200_),
        .dout(new_Jinkela_wire_10342)
    );

    bfr new_Jinkela_buffer_6152 (
        .din(new_Jinkela_wire_7517),
        .dout(new_Jinkela_wire_7518)
    );

    bfr new_Jinkela_buffer_2931 (
        .din(N54),
        .dout(new_Jinkela_wire_3355)
    );

    bfr new_Jinkela_buffer_8072 (
        .din(new_Jinkela_wire_10166),
        .dout(new_Jinkela_wire_10167)
    );

    and_bi n_1447_ (
        .a(new_Jinkela_wire_4664),
        .b(new_Jinkela_wire_8941),
        .c(n_0716_)
    );

    and_bb n_2161_ (
        .a(new_Jinkela_wire_5158),
        .b(new_Jinkela_wire_1411),
        .c(n_0053_)
    );

    bfr new_Jinkela_buffer_6133 (
        .din(new_Jinkela_wire_7494),
        .dout(new_Jinkela_wire_7495)
    );

    bfr new_Jinkela_buffer_8130 (
        .din(new_Jinkela_wire_10231),
        .dout(new_Jinkela_wire_10232)
    );

    bfr new_Jinkela_buffer_2765 (
        .din(new_Jinkela_wire_3179),
        .dout(new_Jinkela_wire_3180)
    );

    and_bi n_1448_ (
        .a(new_Jinkela_wire_8940),
        .b(new_Jinkela_wire_4663),
        .c(n_0717_)
    );

    and_bi n_2162_ (
        .a(new_Jinkela_wire_7461),
        .b(new_Jinkela_wire_4538),
        .c(n_0054_)
    );

    spl4L new_Jinkela_splitter_543 (
        .a(n_0890_),
        .d(new_Jinkela_wire_7683),
        .b(new_Jinkela_wire_7684),
        .e(new_Jinkela_wire_7685),
        .c(new_Jinkela_wire_7686)
    );

    bfr new_Jinkela_buffer_2807 (
        .din(new_Jinkela_wire_3226),
        .dout(new_Jinkela_wire_3227)
    );

    bfr new_Jinkela_buffer_8073 (
        .din(new_Jinkela_wire_10167),
        .dout(new_Jinkela_wire_10168)
    );

    or_bb n_1449_ (
        .a(n_0717_),
        .b(n_0716_),
        .c(new_net_2507)
    );

    and_ii n_2163_ (
        .a(new_Jinkela_wire_7235),
        .b(new_Jinkela_wire_7339),
        .c(n_0055_)
    );

    bfr new_Jinkela_buffer_6134 (
        .din(new_Jinkela_wire_7495),
        .dout(new_Jinkela_wire_7496)
    );

    bfr new_Jinkela_buffer_8131 (
        .din(new_Jinkela_wire_10232),
        .dout(new_Jinkela_wire_10233)
    );

    bfr new_Jinkela_buffer_2766 (
        .din(new_Jinkela_wire_3180),
        .dout(new_Jinkela_wire_3181)
    );

    and_bb n_1450_ (
        .a(N9),
        .b(N12),
        .c(n_0718_)
    );

    and_ii n_2164_ (
        .a(new_Jinkela_wire_7772),
        .b(new_Jinkela_wire_4186),
        .c(n_0056_)
    );

    bfr new_Jinkela_buffer_6215 (
        .din(new_Jinkela_wire_7588),
        .dout(new_Jinkela_wire_7589)
    );

    bfr new_Jinkela_buffer_6153 (
        .din(new_Jinkela_wire_7518),
        .dout(new_Jinkela_wire_7519)
    );

    bfr new_Jinkela_buffer_2860 (
        .din(new_Jinkela_wire_3283),
        .dout(new_Jinkela_wire_3284)
    );

    bfr new_Jinkela_buffer_8074 (
        .din(new_Jinkela_wire_10168),
        .dout(new_Jinkela_wire_10169)
    );

    and_bi n_1451_ (
        .a(new_Jinkela_wire_1267),
        .b(new_Jinkela_wire_1794),
        .c(n_0719_)
    );

    and_bi n_2165_ (
        .a(new_Jinkela_wire_8306),
        .b(n_0056_),
        .c(n_0057_)
    );

    bfr new_Jinkela_buffer_6135 (
        .din(new_Jinkela_wire_7496),
        .dout(new_Jinkela_wire_7497)
    );

    bfr new_Jinkela_buffer_8193 (
        .din(new_Jinkela_wire_10296),
        .dout(new_Jinkela_wire_10297)
    );

    bfr new_Jinkela_buffer_2767 (
        .din(new_Jinkela_wire_3181),
        .dout(new_Jinkela_wire_3182)
    );

    and_ii n_1452_ (
        .a(new_Jinkela_wire_6317),
        .b(new_Jinkela_wire_9453),
        .c(n_0720_)
    );

    or_bi n_2166_ (
        .a(new_Jinkela_wire_10442),
        .b(new_Jinkela_wire_7955),
        .c(n_0058_)
    );

    bfr new_Jinkela_buffer_6179 (
        .din(new_Jinkela_wire_7552),
        .dout(new_Jinkela_wire_7553)
    );

    bfr new_Jinkela_buffer_2808 (
        .din(new_Jinkela_wire_3227),
        .dout(new_Jinkela_wire_3228)
    );

    bfr new_Jinkela_buffer_8075 (
        .din(new_Jinkela_wire_10169),
        .dout(new_Jinkela_wire_10170)
    );

    and_bi n_1453_ (
        .a(new_Jinkela_wire_1178),
        .b(new_Jinkela_wire_2466),
        .c(n_0721_)
    );

    and_bi n_2167_ (
        .a(n_0058_),
        .b(new_Jinkela_wire_6939),
        .c(n_0059_)
    );

    bfr new_Jinkela_buffer_6136 (
        .din(new_Jinkela_wire_7497),
        .dout(new_Jinkela_wire_7498)
    );

    bfr new_Jinkela_buffer_8132 (
        .din(new_Jinkela_wire_10233),
        .dout(new_Jinkela_wire_10234)
    );

    bfr new_Jinkela_buffer_2768 (
        .din(new_Jinkela_wire_3182),
        .dout(new_Jinkela_wire_3183)
    );

    or_ii n_1454_ (
        .a(new_Jinkela_wire_4048),
        .b(new_Jinkela_wire_10389),
        .c(n_0722_)
    );

    and_ii n_2168_ (
        .a(new_Jinkela_wire_8482),
        .b(new_Jinkela_wire_3576),
        .c(n_0060_)
    );

    bfr new_Jinkela_buffer_6154 (
        .din(new_Jinkela_wire_7519),
        .dout(new_Jinkela_wire_7520)
    );

    bfr new_Jinkela_buffer_2925 (
        .din(new_Jinkela_wire_3348),
        .dout(new_Jinkela_wire_3349)
    );

    bfr new_Jinkela_buffer_8076 (
        .din(new_Jinkela_wire_10170),
        .dout(new_Jinkela_wire_10171)
    );

    and_ii n_1455_ (
        .a(new_Jinkela_wire_4045),
        .b(new_Jinkela_wire_9448),
        .c(n_0723_)
    );

    and_ii n_2169_ (
        .a(new_Jinkela_wire_4536),
        .b(new_Jinkela_wire_7335),
        .c(n_0061_)
    );

    bfr new_Jinkela_buffer_6137 (
        .din(new_Jinkela_wire_7498),
        .dout(new_Jinkela_wire_7499)
    );

    bfr new_Jinkela_buffer_2769 (
        .din(new_Jinkela_wire_3183),
        .dout(new_Jinkela_wire_3184)
    );

    and_bb n_1456_ (
        .a(new_Jinkela_wire_6942),
        .b(new_Jinkela_wire_6320),
        .c(n_0724_)
    );

    and_bb n_2170_ (
        .a(new_Jinkela_wire_9253),
        .b(new_Jinkela_wire_8664),
        .c(n_0062_)
    );

    bfr new_Jinkela_buffer_8239 (
        .din(new_net_2517),
        .dout(new_Jinkela_wire_10343)
    );

    bfr new_Jinkela_buffer_8077 (
        .din(new_Jinkela_wire_10171),
        .dout(new_Jinkela_wire_10172)
    );

    bfr new_Jinkela_buffer_2809 (
        .din(new_Jinkela_wire_3228),
        .dout(new_Jinkela_wire_3229)
    );

    and_bi n_1457_ (
        .a(n_0722_),
        .b(n_0724_),
        .c(n_0725_)
    );

    and_ii n_2171_ (
        .a(new_Jinkela_wire_10433),
        .b(new_Jinkela_wire_6929),
        .c(n_0063_)
    );

    bfr new_Jinkela_buffer_6305 (
        .din(n_0477_),
        .dout(new_Jinkela_wire_7687)
    );

    bfr new_Jinkela_buffer_6155 (
        .din(new_Jinkela_wire_7520),
        .dout(new_Jinkela_wire_7521)
    );

    bfr new_Jinkela_buffer_2770 (
        .din(new_Jinkela_wire_3184),
        .dout(new_Jinkela_wire_3185)
    );

    bfr new_Jinkela_buffer_8133 (
        .din(new_Jinkela_wire_10234),
        .dout(new_Jinkela_wire_10235)
    );

    and_bi n_1458_ (
        .a(new_Jinkela_wire_1338),
        .b(new_Jinkela_wire_348),
        .c(n_0726_)
    );

    and_ii n_2172_ (
        .a(new_Jinkela_wire_4181),
        .b(new_Jinkela_wire_5643),
        .c(n_0064_)
    );

    bfr new_Jinkela_buffer_6180 (
        .din(new_Jinkela_wire_7553),
        .dout(new_Jinkela_wire_7554)
    );

    bfr new_Jinkela_buffer_2861 (
        .din(new_Jinkela_wire_3284),
        .dout(new_Jinkela_wire_3285)
    );

    bfr new_Jinkela_buffer_8078 (
        .din(new_Jinkela_wire_10172),
        .dout(new_Jinkela_wire_10173)
    );

    and_ii n_1459_ (
        .a(new_Jinkela_wire_5146),
        .b(new_Jinkela_wire_9462),
        .c(n_0727_)
    );

    and_bb n_2173_ (
        .a(new_Jinkela_wire_3721),
        .b(new_Jinkela_wire_9112),
        .c(n_0065_)
    );

    bfr new_Jinkela_buffer_6156 (
        .din(new_Jinkela_wire_7521),
        .dout(new_Jinkela_wire_7522)
    );

    bfr new_Jinkela_buffer_2771 (
        .din(new_Jinkela_wire_3185),
        .dout(new_Jinkela_wire_3186)
    );

    and_bi n_1460_ (
        .a(new_Jinkela_wire_1239),
        .b(new_Jinkela_wire_795),
        .c(n_0728_)
    );

    and_bb n_2174_ (
        .a(new_Jinkela_wire_7454),
        .b(new_Jinkela_wire_7415),
        .c(n_0066_)
    );

    spl2 new_Jinkela_splitter_845 (
        .a(n_0823_),
        .b(new_Jinkela_wire_10360),
        .c(new_Jinkela_wire_10361)
    );

    bfr new_Jinkela_buffer_6344 (
        .din(n_1318_),
        .dout(new_Jinkela_wire_7728)
    );

    bfr new_Jinkela_buffer_2810 (
        .din(new_Jinkela_wire_3229),
        .dout(new_Jinkela_wire_3230)
    );

    bfr new_Jinkela_buffer_8079 (
        .din(new_Jinkela_wire_10173),
        .dout(new_Jinkela_wire_10174)
    );

    and_bb n_1461_ (
        .a(new_Jinkela_wire_10632),
        .b(new_Jinkela_wire_6744),
        .c(n_0729_)
    );

    or_bi n_2175_ (
        .a(new_Jinkela_wire_9408),
        .b(new_Jinkela_wire_9961),
        .c(n_0067_)
    );

    bfr new_Jinkela_buffer_6216 (
        .din(new_Jinkela_wire_7589),
        .dout(new_Jinkela_wire_7590)
    );

    bfr new_Jinkela_buffer_6157 (
        .din(new_Jinkela_wire_7522),
        .dout(new_Jinkela_wire_7523)
    );

    bfr new_Jinkela_buffer_2772 (
        .din(new_Jinkela_wire_3186),
        .dout(new_Jinkela_wire_3187)
    );

    bfr new_Jinkela_buffer_8134 (
        .din(new_Jinkela_wire_10235),
        .dout(new_Jinkela_wire_10236)
    );

    and_ii n_1462_ (
        .a(new_Jinkela_wire_10629),
        .b(new_Jinkela_wire_9460),
        .c(n_0730_)
    );

    and_bi n_2176_ (
        .a(n_0067_),
        .b(new_Jinkela_wire_7113),
        .c(n_0068_)
    );

    bfr new_Jinkela_buffer_6181 (
        .din(new_Jinkela_wire_7554),
        .dout(new_Jinkela_wire_7555)
    );

    bfr new_Jinkela_buffer_2928 (
        .din(new_Jinkela_wire_3351),
        .dout(new_Jinkela_wire_3352)
    );

    bfr new_Jinkela_buffer_8080 (
        .din(new_Jinkela_wire_10174),
        .dout(new_Jinkela_wire_10175)
    );

    and_bb n_1463_ (
        .a(new_Jinkela_wire_4967),
        .b(new_Jinkela_wire_5149),
        .c(n_0731_)
    );

    and_bb n_2177_ (
        .a(new_Jinkela_wire_9982),
        .b(new_Jinkela_wire_8377),
        .c(n_0069_)
    );

    bfr new_Jinkela_buffer_6158 (
        .din(new_Jinkela_wire_7523),
        .dout(new_Jinkela_wire_7524)
    );

    bfr new_Jinkela_buffer_2773 (
        .din(new_Jinkela_wire_3187),
        .dout(new_Jinkela_wire_3188)
    );

    bfr new_Jinkela_buffer_8194 (
        .din(new_Jinkela_wire_10297),
        .dout(new_Jinkela_wire_10298)
    );

    or_bb n_1464_ (
        .a(n_0731_),
        .b(n_0729_),
        .c(n_0732_)
    );

    and_bi n_2178_ (
        .a(new_Jinkela_wire_8842),
        .b(n_0069_),
        .c(n_0070_)
    );

    bfr new_Jinkela_buffer_8081 (
        .din(new_Jinkela_wire_10175),
        .dout(new_Jinkela_wire_10176)
    );

    bfr new_Jinkela_buffer_2811 (
        .din(new_Jinkela_wire_3230),
        .dout(new_Jinkela_wire_3231)
    );

    and_bi n_1465_ (
        .a(new_Jinkela_wire_1402),
        .b(new_Jinkela_wire_1384),
        .c(n_0733_)
    );

    and_bi n_2179_ (
        .a(new_Jinkela_wire_10134),
        .b(new_Jinkela_wire_9580),
        .c(n_0071_)
    );

    bfr new_Jinkela_buffer_6276 (
        .din(new_Jinkela_wire_7653),
        .dout(new_Jinkela_wire_7654)
    );

    bfr new_Jinkela_buffer_6159 (
        .din(new_Jinkela_wire_7524),
        .dout(new_Jinkela_wire_7525)
    );

    bfr new_Jinkela_buffer_2774 (
        .din(new_Jinkela_wire_3188),
        .dout(new_Jinkela_wire_3189)
    );

    bfr new_Jinkela_buffer_8135 (
        .din(new_Jinkela_wire_10236),
        .dout(new_Jinkela_wire_10237)
    );

    and_bb n_1466_ (
        .a(new_Jinkela_wire_3354),
        .b(new_Jinkela_wire_1281),
        .c(n_0734_)
    );

    and_ii n_2180_ (
        .a(n_0071_),
        .b(new_Jinkela_wire_5448),
        .c(n_0072_)
    );

    bfr new_Jinkela_buffer_6182 (
        .din(new_Jinkela_wire_7555),
        .dout(new_Jinkela_wire_7556)
    );

    bfr new_Jinkela_buffer_2862 (
        .din(new_Jinkela_wire_3285),
        .dout(new_Jinkela_wire_3286)
    );

    bfr new_Jinkela_buffer_8082 (
        .din(new_Jinkela_wire_10176),
        .dout(new_Jinkela_wire_10177)
    );

    and_ii n_1467_ (
        .a(new_Jinkela_wire_4505),
        .b(new_Jinkela_wire_7341),
        .c(n_0735_)
    );

    and_ii n_2181_ (
        .a(new_Jinkela_wire_4434),
        .b(new_Jinkela_wire_5499),
        .c(n_0073_)
    );

    bfr new_Jinkela_buffer_6160 (
        .din(new_Jinkela_wire_7525),
        .dout(new_Jinkela_wire_7526)
    );

    bfr new_Jinkela_buffer_2812 (
        .din(new_Jinkela_wire_3231),
        .dout(new_Jinkela_wire_3232)
    );

    spl4L new_Jinkela_splitter_846 (
        .a(n_0857_),
        .d(new_Jinkela_wire_10362),
        .b(new_Jinkela_wire_10363),
        .e(new_Jinkela_wire_10364),
        .c(new_Jinkela_wire_10365)
    );

    and_bi n_1468_ (
        .a(new_Jinkela_wire_3434),
        .b(new_Jinkela_wire_1302),
        .c(n_0736_)
    );

    or_bb n_2182_ (
        .a(new_Jinkela_wire_5636),
        .b(new_Jinkela_wire_8811),
        .c(n_0074_)
    );

    bfr new_Jinkela_buffer_8240 (
        .din(new_Jinkela_wire_10343),
        .dout(new_Jinkela_wire_10344)
    );

    bfr new_Jinkela_buffer_8083 (
        .din(new_Jinkela_wire_10177),
        .dout(new_Jinkela_wire_10178)
    );

    bfr new_Jinkela_buffer_2926 (
        .din(new_Jinkela_wire_3349),
        .dout(new_Jinkela_wire_3350)
    );

    and_bb n_1469_ (
        .a(new_Jinkela_wire_185),
        .b(new_Jinkela_wire_1303),
        .c(n_0737_)
    );

    and_bi n_2183_ (
        .a(new_Jinkela_wire_9245),
        .b(new_Jinkela_wire_4531),
        .c(n_0075_)
    );

    bfr new_Jinkela_buffer_6217 (
        .din(new_Jinkela_wire_7590),
        .dout(new_Jinkela_wire_7591)
    );

    bfr new_Jinkela_buffer_6161 (
        .din(new_Jinkela_wire_7526),
        .dout(new_Jinkela_wire_7527)
    );

    bfr new_Jinkela_buffer_2813 (
        .din(new_Jinkela_wire_3232),
        .dout(new_Jinkela_wire_3233)
    );

    bfr new_Jinkela_buffer_8136 (
        .din(new_Jinkela_wire_10237),
        .dout(new_Jinkela_wire_10238)
    );

    and_ii n_1470_ (
        .a(new_Jinkela_wire_8361),
        .b(new_Jinkela_wire_6516),
        .c(n_0738_)
    );

    and_ii n_2184_ (
        .a(new_Jinkela_wire_5635),
        .b(new_Jinkela_wire_8810),
        .c(n_0076_)
    );

    bfr new_Jinkela_buffer_6183 (
        .din(new_Jinkela_wire_7556),
        .dout(new_Jinkela_wire_7557)
    );

    bfr new_Jinkela_buffer_2863 (
        .din(new_Jinkela_wire_3286),
        .dout(new_Jinkela_wire_3287)
    );

    bfr new_Jinkela_buffer_8084 (
        .din(new_Jinkela_wire_10178),
        .dout(new_Jinkela_wire_10179)
    );

    and_bb n_1471_ (
        .a(new_Jinkela_wire_5057),
        .b(new_Jinkela_wire_9299),
        .c(n_0739_)
    );

    or_bb n_2185_ (
        .a(new_Jinkela_wire_5145),
        .b(new_Jinkela_wire_9244),
        .c(n_0077_)
    );

    bfr new_Jinkela_buffer_6162 (
        .din(new_Jinkela_wire_7527),
        .dout(new_Jinkela_wire_7528)
    );

    bfr new_Jinkela_buffer_2814 (
        .din(new_Jinkela_wire_3233),
        .dout(new_Jinkela_wire_3234)
    );

    bfr new_Jinkela_buffer_8195 (
        .din(new_Jinkela_wire_10298),
        .dout(new_Jinkela_wire_10299)
    );

    and_ii n_1472_ (
        .a(new_Jinkela_wire_5055),
        .b(new_Jinkela_wire_9298),
        .c(n_0740_)
    );

    and_bi n_2186_ (
        .a(new_Jinkela_wire_8357),
        .b(new_Jinkela_wire_4013),
        .c(new_net_2545)
    );

    bfr new_Jinkela_buffer_8085 (
        .din(new_Jinkela_wire_10179),
        .dout(new_Jinkela_wire_10180)
    );

    bfr new_Jinkela_buffer_2935 (
        .din(N225),
        .dout(new_Jinkela_wire_3359)
    );

    and_ii n_1473_ (
        .a(n_0740_),
        .b(n_0739_),
        .c(n_0741_)
    );

    and_ii n_2187_ (
        .a(new_Jinkela_wire_3563),
        .b(new_Jinkela_wire_7097),
        .c(n_0078_)
    );

    bfr new_Jinkela_buffer_6163 (
        .din(new_Jinkela_wire_7528),
        .dout(new_Jinkela_wire_7529)
    );

    bfr new_Jinkela_buffer_2815 (
        .din(new_Jinkela_wire_3234),
        .dout(new_Jinkela_wire_3235)
    );

    bfr new_Jinkela_buffer_8137 (
        .din(new_Jinkela_wire_10238),
        .dout(new_Jinkela_wire_10239)
    );

    or_bb n_1474_ (
        .a(new_Jinkela_wire_9958),
        .b(new_Jinkela_wire_6332),
        .c(n_0742_)
    );

    inv n_2188_ (
        .din(new_Jinkela_wire_9336),
        .dout(n_0079_)
    );

    bfr new_Jinkela_buffer_6184 (
        .din(new_Jinkela_wire_7557),
        .dout(new_Jinkela_wire_7558)
    );

    bfr new_Jinkela_buffer_2864 (
        .din(new_Jinkela_wire_3287),
        .dout(new_Jinkela_wire_3288)
    );

    bfr new_Jinkela_buffer_8086 (
        .din(new_Jinkela_wire_10180),
        .dout(new_Jinkela_wire_10181)
    );

    and_bb n_1475_ (
        .a(new_Jinkela_wire_9957),
        .b(new_Jinkela_wire_6331),
        .c(n_0743_)
    );

    inv n_2189_ (
        .din(new_Jinkela_wire_9110),
        .dout(n_0080_)
    );

    bfr new_Jinkela_buffer_6164 (
        .din(new_Jinkela_wire_7529),
        .dout(new_Jinkela_wire_7530)
    );

    bfr new_Jinkela_buffer_2816 (
        .din(new_Jinkela_wire_3235),
        .dout(new_Jinkela_wire_3236)
    );

    and_bi n_1476_ (
        .a(n_0742_),
        .b(n_0743_),
        .c(n_0744_)
    );

    inv n_2190_ (
        .din(new_Jinkela_wire_3720),
        .dout(n_0081_)
    );

    bfr new_Jinkela_buffer_8087 (
        .din(new_Jinkela_wire_10181),
        .dout(new_Jinkela_wire_10182)
    );

    bfr new_Jinkela_buffer_2929 (
        .din(new_Jinkela_wire_3352),
        .dout(new_Jinkela_wire_3353)
    );

    and_ii n_1477_ (
        .a(new_Jinkela_wire_9555),
        .b(new_Jinkela_wire_6523),
        .c(n_0745_)
    );

    and_bi n_2191_ (
        .a(new_Jinkela_wire_7414),
        .b(new_Jinkela_wire_5935),
        .c(n_0082_)
    );

    bfr new_Jinkela_buffer_6218 (
        .din(new_Jinkela_wire_7591),
        .dout(new_Jinkela_wire_7592)
    );

    bfr new_Jinkela_buffer_6165 (
        .din(new_Jinkela_wire_7530),
        .dout(new_Jinkela_wire_7531)
    );

    bfr new_Jinkela_buffer_2817 (
        .din(new_Jinkela_wire_3236),
        .dout(new_Jinkela_wire_3237)
    );

    bfr new_Jinkela_buffer_8138 (
        .din(new_Jinkela_wire_10239),
        .dout(new_Jinkela_wire_10240)
    );

    and_bb n_1478_ (
        .a(new_Jinkela_wire_9554),
        .b(new_Jinkela_wire_6522),
        .c(n_0746_)
    );

    and_bi n_2192_ (
        .a(new_Jinkela_wire_4044),
        .b(new_Jinkela_wire_8380),
        .c(n_0083_)
    );

    bfr new_Jinkela_buffer_6185 (
        .din(new_Jinkela_wire_7558),
        .dout(new_Jinkela_wire_7559)
    );

    bfr new_Jinkela_buffer_2865 (
        .din(new_Jinkela_wire_3288),
        .dout(new_Jinkela_wire_3289)
    );

    bfr new_Jinkela_buffer_8088 (
        .din(new_Jinkela_wire_10182),
        .dout(new_Jinkela_wire_10183)
    );

    and_ii n_1479_ (
        .a(n_0746_),
        .b(n_0745_),
        .c(n_0747_)
    );

    and_bi n_2193_ (
        .a(new_Jinkela_wire_8284),
        .b(new_Jinkela_wire_3764),
        .c(n_0084_)
    );

    bfr new_Jinkela_buffer_6166 (
        .din(new_Jinkela_wire_7531),
        .dout(new_Jinkela_wire_7532)
    );

    bfr new_Jinkela_buffer_2818 (
        .din(new_Jinkela_wire_3237),
        .dout(new_Jinkela_wire_3238)
    );

    bfr new_Jinkela_buffer_8196 (
        .din(new_Jinkela_wire_10299),
        .dout(new_Jinkela_wire_10300)
    );

    and_bi n_1480_ (
        .a(new_Jinkela_wire_1997),
        .b(new_Jinkela_wire_1340),
        .c(n_0748_)
    );

    and_ii n_2194_ (
        .a(n_0084_),
        .b(new_Jinkela_wire_8508),
        .c(n_0085_)
    );

    bfr new_Jinkela_buffer_8089 (
        .din(new_Jinkela_wire_10183),
        .dout(new_Jinkela_wire_10184)
    );

    bfr new_Jinkela_buffer_2932 (
        .din(new_Jinkela_wire_3355),
        .dout(new_Jinkela_wire_3356)
    );

    and_bb n_1481_ (
        .a(new_Jinkela_wire_686),
        .b(new_Jinkela_wire_1219),
        .c(n_0749_)
    );

    and_bi n_2195_ (
        .a(new_Jinkela_wire_7456),
        .b(new_Jinkela_wire_4913),
        .c(n_0086_)
    );

    bfr new_Jinkela_buffer_6277 (
        .din(new_Jinkela_wire_7654),
        .dout(new_Jinkela_wire_7655)
    );

    bfr new_Jinkela_buffer_6167 (
        .din(new_Jinkela_wire_7532),
        .dout(new_Jinkela_wire_7533)
    );

    bfr new_Jinkela_buffer_2819 (
        .din(new_Jinkela_wire_3238),
        .dout(new_Jinkela_wire_3239)
    );

    bfr new_Jinkela_buffer_8139 (
        .din(new_Jinkela_wire_10240),
        .dout(new_Jinkela_wire_10241)
    );

    or_bb n_1482_ (
        .a(new_Jinkela_wire_9553),
        .b(new_Jinkela_wire_8280),
        .c(n_0750_)
    );

    and_bi n_2196_ (
        .a(new_Jinkela_wire_4912),
        .b(new_Jinkela_wire_7455),
        .c(n_0087_)
    );

    bfr new_Jinkela_buffer_6186 (
        .din(new_Jinkela_wire_7559),
        .dout(new_Jinkela_wire_7560)
    );

    bfr new_Jinkela_buffer_2866 (
        .din(new_Jinkela_wire_3289),
        .dout(new_Jinkela_wire_3290)
    );

    bfr new_Jinkela_buffer_8090 (
        .din(new_Jinkela_wire_10184),
        .dout(new_Jinkela_wire_10185)
    );

    and_bi n_1483_ (
        .a(new_Jinkela_wire_1387),
        .b(new_Jinkela_wire_1790),
        .c(n_0751_)
    );

    or_bb n_2197_ (
        .a(n_0087_),
        .b(n_0086_),
        .c(new_net_2505)
    );

    bfr new_Jinkela_buffer_6168 (
        .din(new_Jinkela_wire_7533),
        .dout(new_Jinkela_wire_7534)
    );

    bfr new_Jinkela_buffer_2820 (
        .din(new_Jinkela_wire_3239),
        .dout(new_Jinkela_wire_3240)
    );

    and_ii n_1484_ (
        .a(n_0751_),
        .b(new_Jinkela_wire_9439),
        .c(n_0752_)
    );

    and_bi n_2198_ (
        .a(new_Jinkela_wire_7984),
        .b(new_Jinkela_wire_8283),
        .c(n_0088_)
    );

    bfr new_Jinkela_buffer_8241 (
        .din(new_Jinkela_wire_10344),
        .dout(new_Jinkela_wire_10345)
    );

    bfr new_Jinkela_buffer_649 (
        .din(new_Jinkela_wire_701),
        .dout(new_Jinkela_wire_702)
    );

    bfr new_Jinkela_buffer_1283 (
        .din(new_Jinkela_wire_1603),
        .dout(new_Jinkela_wire_1604)
    );

    bfr new_Jinkela_buffer_5329 (
        .din(new_Jinkela_wire_6387),
        .dout(new_Jinkela_wire_6388)
    );

    bfr new_Jinkela_buffer_595 (
        .din(new_Jinkela_wire_643),
        .dout(new_Jinkela_wire_644)
    );

    bfr new_Jinkela_buffer_1319 (
        .din(new_Jinkela_wire_1644),
        .dout(new_Jinkela_wire_1645)
    );

    bfr new_Jinkela_buffer_5361 (
        .din(new_Jinkela_wire_6440),
        .dout(new_Jinkela_wire_6441)
    );

    bfr new_Jinkela_buffer_716 (
        .din(new_Jinkela_wire_772),
        .dout(new_Jinkela_wire_773)
    );

    bfr new_Jinkela_buffer_1284 (
        .din(new_Jinkela_wire_1604),
        .dout(new_Jinkela_wire_1605)
    );

    bfr new_Jinkela_buffer_5330 (
        .din(new_Jinkela_wire_6388),
        .dout(new_Jinkela_wire_6389)
    );

    bfr new_Jinkela_buffer_712 (
        .din(new_Jinkela_wire_766),
        .dout(new_Jinkela_wire_767)
    );

    bfr new_Jinkela_buffer_596 (
        .din(new_Jinkela_wire_644),
        .dout(new_Jinkela_wire_645)
    );

    spl2 new_Jinkela_splitter_103 (
        .a(new_Jinkela_wire_1708),
        .b(new_Jinkela_wire_1709),
        .c(new_Jinkela_wire_1710)
    );

    bfr new_Jinkela_buffer_5346 (
        .din(new_Jinkela_wire_6419),
        .dout(new_Jinkela_wire_6420)
    );

    bfr new_Jinkela_buffer_1381 (
        .din(new_Jinkela_wire_1710),
        .dout(new_Jinkela_wire_1711)
    );

    bfr new_Jinkela_buffer_650 (
        .din(new_Jinkela_wire_702),
        .dout(new_Jinkela_wire_703)
    );

    bfr new_Jinkela_buffer_1285 (
        .din(new_Jinkela_wire_1605),
        .dout(new_Jinkela_wire_1606)
    );

    bfr new_Jinkela_buffer_597 (
        .din(new_Jinkela_wire_645),
        .dout(new_Jinkela_wire_646)
    );

    bfr new_Jinkela_buffer_1320 (
        .din(new_Jinkela_wire_1645),
        .dout(new_Jinkela_wire_1646)
    );

    bfr new_Jinkela_buffer_5347 (
        .din(new_Jinkela_wire_6420),
        .dout(new_Jinkela_wire_6421)
    );

    bfr new_Jinkela_buffer_1286 (
        .din(new_Jinkela_wire_1606),
        .dout(new_Jinkela_wire_1607)
    );

    bfr new_Jinkela_buffer_5407 (
        .din(new_Jinkela_wire_6486),
        .dout(new_Jinkela_wire_6487)
    );

    bfr new_Jinkela_buffer_5362 (
        .din(new_Jinkela_wire_6441),
        .dout(new_Jinkela_wire_6442)
    );

    bfr new_Jinkela_buffer_598 (
        .din(new_Jinkela_wire_646),
        .dout(new_Jinkela_wire_647)
    );

    bfr new_Jinkela_buffer_5348 (
        .din(new_Jinkela_wire_6421),
        .dout(new_Jinkela_wire_6422)
    );

    bfr new_Jinkela_buffer_651 (
        .din(new_Jinkela_wire_703),
        .dout(new_Jinkela_wire_704)
    );

    bfr new_Jinkela_buffer_1287 (
        .din(new_Jinkela_wire_1607),
        .dout(new_Jinkela_wire_1608)
    );

    bfr new_Jinkela_buffer_599 (
        .din(new_Jinkela_wire_647),
        .dout(new_Jinkela_wire_648)
    );

    bfr new_Jinkela_buffer_1321 (
        .din(new_Jinkela_wire_1646),
        .dout(new_Jinkela_wire_1647)
    );

    bfr new_Jinkela_buffer_5349 (
        .din(new_Jinkela_wire_6422),
        .dout(new_Jinkela_wire_6423)
    );

    bfr new_Jinkela_buffer_723 (
        .din(N224),
        .dout(new_Jinkela_wire_780)
    );

    bfr new_Jinkela_buffer_1444 (
        .din(new_Jinkela_wire_1776),
        .dout(new_Jinkela_wire_1777)
    );

    bfr new_Jinkela_buffer_713 (
        .din(new_Jinkela_wire_767),
        .dout(new_Jinkela_wire_768)
    );

    bfr new_Jinkela_buffer_5363 (
        .din(new_Jinkela_wire_6442),
        .dout(new_Jinkela_wire_6443)
    );

    bfr new_Jinkela_buffer_600 (
        .din(new_Jinkela_wire_648),
        .dout(new_Jinkela_wire_649)
    );

    bfr new_Jinkela_buffer_1322 (
        .din(new_Jinkela_wire_1647),
        .dout(new_Jinkela_wire_1648)
    );

    bfr new_Jinkela_buffer_5350 (
        .din(new_Jinkela_wire_6423),
        .dout(new_Jinkela_wire_6424)
    );

    bfr new_Jinkela_buffer_652 (
        .din(new_Jinkela_wire_704),
        .dout(new_Jinkela_wire_705)
    );

    bfr new_Jinkela_buffer_1447 (
        .din(new_Jinkela_wire_1779),
        .dout(new_Jinkela_wire_1780)
    );

    spl2 new_Jinkela_splitter_419 (
        .a(n_0850_),
        .b(new_Jinkela_wire_6517),
        .c(new_Jinkela_wire_6518)
    );

    bfr new_Jinkela_buffer_601 (
        .din(new_Jinkela_wire_649),
        .dout(new_Jinkela_wire_650)
    );

    bfr new_Jinkela_buffer_1323 (
        .din(new_Jinkela_wire_1648),
        .dout(new_Jinkela_wire_1649)
    );

    bfr new_Jinkela_buffer_5351 (
        .din(new_Jinkela_wire_6424),
        .dout(new_Jinkela_wire_6425)
    );

    bfr new_Jinkela_buffer_1382 (
        .din(new_Jinkela_wire_1711),
        .dout(new_Jinkela_wire_1712)
    );

    bfr new_Jinkela_buffer_5408 (
        .din(new_Jinkela_wire_6487),
        .dout(new_Jinkela_wire_6488)
    );

    bfr new_Jinkela_buffer_5364 (
        .din(new_Jinkela_wire_6443),
        .dout(new_Jinkela_wire_6444)
    );

    bfr new_Jinkela_buffer_602 (
        .din(new_Jinkela_wire_650),
        .dout(new_Jinkela_wire_651)
    );

    bfr new_Jinkela_buffer_1324 (
        .din(new_Jinkela_wire_1649),
        .dout(new_Jinkela_wire_1650)
    );

    bfr new_Jinkela_buffer_5352 (
        .din(new_Jinkela_wire_6425),
        .dout(new_Jinkela_wire_6426)
    );

    bfr new_Jinkela_buffer_653 (
        .din(new_Jinkela_wire_705),
        .dout(new_Jinkela_wire_706)
    );

    bfr new_Jinkela_buffer_1445 (
        .din(new_Jinkela_wire_1777),
        .dout(new_Jinkela_wire_1778)
    );

    bfr new_Jinkela_buffer_603 (
        .din(new_Jinkela_wire_651),
        .dout(new_Jinkela_wire_652)
    );

    bfr new_Jinkela_buffer_1325 (
        .din(new_Jinkela_wire_1650),
        .dout(new_Jinkela_wire_1651)
    );

    bfr new_Jinkela_buffer_5353 (
        .din(new_Jinkela_wire_6426),
        .dout(new_Jinkela_wire_6427)
    );

    bfr new_Jinkela_buffer_717 (
        .din(new_Jinkela_wire_773),
        .dout(new_Jinkela_wire_774)
    );

    bfr new_Jinkela_buffer_1383 (
        .din(new_Jinkela_wire_1712),
        .dout(new_Jinkela_wire_1713)
    );

    spl2 new_Jinkela_splitter_421 (
        .a(n_0712_),
        .b(new_Jinkela_wire_6528),
        .c(new_Jinkela_wire_6529)
    );

    bfr new_Jinkela_buffer_714 (
        .din(new_Jinkela_wire_768),
        .dout(new_Jinkela_wire_769)
    );

    bfr new_Jinkela_buffer_5365 (
        .din(new_Jinkela_wire_6444),
        .dout(new_Jinkela_wire_6445)
    );

    bfr new_Jinkela_buffer_604 (
        .din(new_Jinkela_wire_652),
        .dout(new_Jinkela_wire_653)
    );

    bfr new_Jinkela_buffer_1326 (
        .din(new_Jinkela_wire_1651),
        .dout(new_Jinkela_wire_1652)
    );

    bfr new_Jinkela_buffer_654 (
        .din(new_Jinkela_wire_706),
        .dout(new_Jinkela_wire_707)
    );

    bfr new_Jinkela_buffer_1454 (
        .din(N157),
        .dout(new_Jinkela_wire_1787)
    );

    bfr new_Jinkela_buffer_5409 (
        .din(new_Jinkela_wire_6488),
        .dout(new_Jinkela_wire_6489)
    );

    bfr new_Jinkela_buffer_5366 (
        .din(new_Jinkela_wire_6445),
        .dout(new_Jinkela_wire_6446)
    );

    bfr new_Jinkela_buffer_605 (
        .din(new_Jinkela_wire_653),
        .dout(new_Jinkela_wire_654)
    );

    bfr new_Jinkela_buffer_1327 (
        .din(new_Jinkela_wire_1652),
        .dout(new_Jinkela_wire_1653)
    );

    spl3L new_Jinkela_splitter_104 (
        .a(new_Jinkela_wire_1713),
        .d(new_Jinkela_wire_1714),
        .b(new_Jinkela_wire_1715),
        .c(new_Jinkela_wire_1716)
    );

    bfr new_Jinkela_buffer_5433 (
        .din(n_0725_),
        .dout(new_Jinkela_wire_6519)
    );

    bfr new_Jinkela_buffer_5367 (
        .din(new_Jinkela_wire_6446),
        .dout(new_Jinkela_wire_6447)
    );

    bfr new_Jinkela_buffer_606 (
        .din(new_Jinkela_wire_654),
        .dout(new_Jinkela_wire_655)
    );

    bfr new_Jinkela_buffer_1328 (
        .din(new_Jinkela_wire_1653),
        .dout(new_Jinkela_wire_1654)
    );

    bfr new_Jinkela_buffer_5440 (
        .din(n_1313_),
        .dout(new_Jinkela_wire_6530)
    );

    bfr new_Jinkela_buffer_655 (
        .din(new_Jinkela_wire_707),
        .dout(new_Jinkela_wire_708)
    );

    bfr new_Jinkela_buffer_1448 (
        .din(new_Jinkela_wire_1780),
        .dout(new_Jinkela_wire_1781)
    );

    bfr new_Jinkela_buffer_5410 (
        .din(new_Jinkela_wire_6489),
        .dout(new_Jinkela_wire_6490)
    );

    bfr new_Jinkela_buffer_5368 (
        .din(new_Jinkela_wire_6447),
        .dout(new_Jinkela_wire_6448)
    );

    bfr new_Jinkela_buffer_607 (
        .din(new_Jinkela_wire_655),
        .dout(new_Jinkela_wire_656)
    );

    bfr new_Jinkela_buffer_1329 (
        .din(new_Jinkela_wire_1654),
        .dout(new_Jinkela_wire_1655)
    );

    bfr new_Jinkela_buffer_720 (
        .din(new_Jinkela_wire_776),
        .dout(new_Jinkela_wire_777)
    );

    bfr new_Jinkela_buffer_1384 (
        .din(new_Jinkela_wire_1716),
        .dout(new_Jinkela_wire_1717)
    );

    bfr new_Jinkela_buffer_5436 (
        .din(n_0182_),
        .dout(new_Jinkela_wire_6524)
    );

    bfr new_Jinkela_buffer_5369 (
        .din(new_Jinkela_wire_6448),
        .dout(new_Jinkela_wire_6449)
    );

    bfr new_Jinkela_buffer_608 (
        .din(new_Jinkela_wire_656),
        .dout(new_Jinkela_wire_657)
    );

    bfr new_Jinkela_buffer_1330 (
        .din(new_Jinkela_wire_1655),
        .dout(new_Jinkela_wire_1656)
    );

    bfr new_Jinkela_buffer_5434 (
        .din(new_Jinkela_wire_6519),
        .dout(new_Jinkela_wire_6520)
    );

    bfr new_Jinkela_buffer_656 (
        .din(new_Jinkela_wire_708),
        .dout(new_Jinkela_wire_709)
    );

    bfr new_Jinkela_buffer_1451 (
        .din(new_Jinkela_wire_1783),
        .dout(new_Jinkela_wire_1784)
    );

    bfr new_Jinkela_buffer_5411 (
        .din(new_Jinkela_wire_6490),
        .dout(new_Jinkela_wire_6491)
    );

    bfr new_Jinkela_buffer_5370 (
        .din(new_Jinkela_wire_6449),
        .dout(new_Jinkela_wire_6450)
    );

    bfr new_Jinkela_buffer_609 (
        .din(new_Jinkela_wire_657),
        .dout(new_Jinkela_wire_658)
    );

    bfr new_Jinkela_buffer_1331 (
        .din(new_Jinkela_wire_1656),
        .dout(new_Jinkela_wire_1657)
    );

    bfr new_Jinkela_buffer_718 (
        .din(new_Jinkela_wire_774),
        .dout(new_Jinkela_wire_775)
    );

    bfr new_Jinkela_buffer_1385 (
        .din(new_Jinkela_wire_1717),
        .dout(new_Jinkela_wire_1718)
    );

    bfr new_Jinkela_buffer_5371 (
        .din(new_Jinkela_wire_6450),
        .dout(new_Jinkela_wire_6451)
    );

    bfr new_Jinkela_buffer_610 (
        .din(new_Jinkela_wire_658),
        .dout(new_Jinkela_wire_659)
    );

    bfr new_Jinkela_buffer_1332 (
        .din(new_Jinkela_wire_1657),
        .dout(new_Jinkela_wire_1658)
    );

    bfr new_Jinkela_buffer_5437 (
        .din(new_Jinkela_wire_6524),
        .dout(new_Jinkela_wire_6525)
    );

    bfr new_Jinkela_buffer_657 (
        .din(new_Jinkela_wire_709),
        .dout(new_Jinkela_wire_710)
    );

    bfr new_Jinkela_buffer_1449 (
        .din(new_Jinkela_wire_1781),
        .dout(new_Jinkela_wire_1782)
    );

    bfr new_Jinkela_buffer_5412 (
        .din(new_Jinkela_wire_6491),
        .dout(new_Jinkela_wire_6492)
    );

    bfr new_Jinkela_buffer_5372 (
        .din(new_Jinkela_wire_6451),
        .dout(new_Jinkela_wire_6452)
    );

    bfr new_Jinkela_buffer_611 (
        .din(new_Jinkela_wire_659),
        .dout(new_Jinkela_wire_660)
    );

    bfr new_Jinkela_buffer_1333 (
        .din(new_Jinkela_wire_1658),
        .dout(new_Jinkela_wire_1659)
    );

    bfr new_Jinkela_buffer_727 (
        .din(N64),
        .dout(new_Jinkela_wire_784)
    );

    bfr new_Jinkela_buffer_1386 (
        .din(new_Jinkela_wire_1718),
        .dout(new_Jinkela_wire_1719)
    );

    bfr new_Jinkela_buffer_5373 (
        .din(new_Jinkela_wire_6452),
        .dout(new_Jinkela_wire_6453)
    );

    bfr new_Jinkela_buffer_612 (
        .din(new_Jinkela_wire_660),
        .dout(new_Jinkela_wire_661)
    );

    bfr new_Jinkela_buffer_1334 (
        .din(new_Jinkela_wire_1659),
        .dout(new_Jinkela_wire_1660)
    );

    bfr new_Jinkela_buffer_5435 (
        .din(new_Jinkela_wire_6520),
        .dout(new_Jinkela_wire_6521)
    );

    bfr new_Jinkela_buffer_658 (
        .din(new_Jinkela_wire_710),
        .dout(new_Jinkela_wire_711)
    );

    bfr new_Jinkela_buffer_1458 (
        .din(N154),
        .dout(new_Jinkela_wire_1791)
    );

    bfr new_Jinkela_buffer_5413 (
        .din(new_Jinkela_wire_6492),
        .dout(new_Jinkela_wire_6493)
    );

    bfr new_Jinkela_buffer_5374 (
        .din(new_Jinkela_wire_6453),
        .dout(new_Jinkela_wire_6454)
    );

    bfr new_Jinkela_buffer_613 (
        .din(new_Jinkela_wire_661),
        .dout(new_Jinkela_wire_662)
    );

    bfr new_Jinkela_buffer_1335 (
        .din(new_Jinkela_wire_1660),
        .dout(new_Jinkela_wire_1661)
    );

    bfr new_Jinkela_buffer_721 (
        .din(new_Jinkela_wire_777),
        .dout(new_Jinkela_wire_778)
    );

    bfr new_Jinkela_buffer_1387 (
        .din(new_Jinkela_wire_1719),
        .dout(new_Jinkela_wire_1720)
    );

    bfr new_Jinkela_buffer_5375 (
        .din(new_Jinkela_wire_6454),
        .dout(new_Jinkela_wire_6455)
    );

    bfr new_Jinkela_buffer_614 (
        .din(new_Jinkela_wire_662),
        .dout(new_Jinkela_wire_663)
    );

    bfr new_Jinkela_buffer_1336 (
        .din(new_Jinkela_wire_1661),
        .dout(new_Jinkela_wire_1662)
    );

    bfr new_Jinkela_buffer_659 (
        .din(new_Jinkela_wire_711),
        .dout(new_Jinkela_wire_712)
    );

    bfr new_Jinkela_buffer_1452 (
        .din(new_Jinkela_wire_1784),
        .dout(new_Jinkela_wire_1785)
    );

    bfr new_Jinkela_buffer_5414 (
        .din(new_Jinkela_wire_6493),
        .dout(new_Jinkela_wire_6494)
    );

    bfr new_Jinkela_buffer_5376 (
        .din(new_Jinkela_wire_6455),
        .dout(new_Jinkela_wire_6456)
    );

    bfr new_Jinkela_buffer_615 (
        .din(new_Jinkela_wire_663),
        .dout(new_Jinkela_wire_664)
    );

    bfr new_Jinkela_buffer_1337 (
        .din(new_Jinkela_wire_1662),
        .dout(new_Jinkela_wire_1663)
    );

    bfr new_Jinkela_buffer_8091 (
        .din(new_Jinkela_wire_10185),
        .dout(new_Jinkela_wire_10186)
    );

    bfr new_Jinkela_buffer_8140 (
        .din(new_Jinkela_wire_10241),
        .dout(new_Jinkela_wire_10242)
    );

    bfr new_Jinkela_buffer_8092 (
        .din(new_Jinkela_wire_10186),
        .dout(new_Jinkela_wire_10187)
    );

    bfr new_Jinkela_buffer_8197 (
        .din(new_Jinkela_wire_10300),
        .dout(new_Jinkela_wire_10301)
    );

    bfr new_Jinkela_buffer_8093 (
        .din(new_Jinkela_wire_10187),
        .dout(new_Jinkela_wire_10188)
    );

    bfr new_Jinkela_buffer_8141 (
        .din(new_Jinkela_wire_10242),
        .dout(new_Jinkela_wire_10243)
    );

    bfr new_Jinkela_buffer_8094 (
        .din(new_Jinkela_wire_10188),
        .dout(new_Jinkela_wire_10189)
    );

    spl2 new_Jinkela_splitter_848 (
        .a(n_1027_),
        .b(new_Jinkela_wire_10378),
        .c(new_Jinkela_wire_10379)
    );

    bfr new_Jinkela_buffer_8095 (
        .din(new_Jinkela_wire_10189),
        .dout(new_Jinkela_wire_10190)
    );

    bfr new_Jinkela_buffer_8142 (
        .din(new_Jinkela_wire_10243),
        .dout(new_Jinkela_wire_10244)
    );

    bfr new_Jinkela_buffer_8096 (
        .din(new_Jinkela_wire_10190),
        .dout(new_Jinkela_wire_10191)
    );

    bfr new_Jinkela_buffer_8198 (
        .din(new_Jinkela_wire_10301),
        .dout(new_Jinkela_wire_10302)
    );

    bfr new_Jinkela_buffer_8097 (
        .din(new_Jinkela_wire_10191),
        .dout(new_Jinkela_wire_10192)
    );

    bfr new_Jinkela_buffer_8143 (
        .din(new_Jinkela_wire_10244),
        .dout(new_Jinkela_wire_10245)
    );

    bfr new_Jinkela_buffer_8098 (
        .din(new_Jinkela_wire_10192),
        .dout(new_Jinkela_wire_10193)
    );

    spl3L new_Jinkela_splitter_847 (
        .a(n_0098_),
        .d(new_Jinkela_wire_10366),
        .b(new_Jinkela_wire_10367),
        .c(new_Jinkela_wire_10368)
    );

    bfr new_Jinkela_buffer_8242 (
        .din(new_Jinkela_wire_10345),
        .dout(new_Jinkela_wire_10346)
    );

    bfr new_Jinkela_buffer_8099 (
        .din(new_Jinkela_wire_10193),
        .dout(new_Jinkela_wire_10194)
    );

    bfr new_Jinkela_buffer_8144 (
        .din(new_Jinkela_wire_10245),
        .dout(new_Jinkela_wire_10246)
    );

    bfr new_Jinkela_buffer_8100 (
        .din(new_Jinkela_wire_10194),
        .dout(new_Jinkela_wire_10195)
    );

    bfr new_Jinkela_buffer_8199 (
        .din(new_Jinkela_wire_10302),
        .dout(new_Jinkela_wire_10303)
    );

    bfr new_Jinkela_buffer_8101 (
        .din(new_Jinkela_wire_10195),
        .dout(new_Jinkela_wire_10196)
    );

    bfr new_Jinkela_buffer_8145 (
        .din(new_Jinkela_wire_10246),
        .dout(new_Jinkela_wire_10247)
    );

    bfr new_Jinkela_buffer_8102 (
        .din(new_Jinkela_wire_10196),
        .dout(new_Jinkela_wire_10197)
    );

    bfr new_Jinkela_buffer_8103 (
        .din(new_Jinkela_wire_10197),
        .dout(new_Jinkela_wire_10198)
    );

    bfr new_Jinkela_buffer_8146 (
        .din(new_Jinkela_wire_10247),
        .dout(new_Jinkela_wire_10248)
    );

    bfr new_Jinkela_buffer_8104 (
        .din(new_Jinkela_wire_10198),
        .dout(new_Jinkela_wire_10199)
    );

    bfr new_Jinkela_buffer_8200 (
        .din(new_Jinkela_wire_10303),
        .dout(new_Jinkela_wire_10304)
    );

    bfr new_Jinkela_buffer_8105 (
        .din(new_Jinkela_wire_10199),
        .dout(new_Jinkela_wire_10200)
    );

    bfr new_Jinkela_buffer_8147 (
        .din(new_Jinkela_wire_10248),
        .dout(new_Jinkela_wire_10249)
    );

    bfr new_Jinkela_buffer_8106 (
        .din(new_Jinkela_wire_10200),
        .dout(new_Jinkela_wire_10201)
    );

    bfr new_Jinkela_buffer_8265 (
        .din(n_0224_),
        .dout(new_Jinkela_wire_10380)
    );

    bfr new_Jinkela_buffer_8243 (
        .din(new_Jinkela_wire_10346),
        .dout(new_Jinkela_wire_10347)
    );

    bfr new_Jinkela_buffer_8107 (
        .din(new_Jinkela_wire_10201),
        .dout(new_Jinkela_wire_10202)
    );

    bfr new_Jinkela_buffer_8148 (
        .din(new_Jinkela_wire_10249),
        .dout(new_Jinkela_wire_10250)
    );

    bfr new_Jinkela_buffer_8108 (
        .din(new_Jinkela_wire_10202),
        .dout(new_Jinkela_wire_10203)
    );

    bfr new_Jinkela_buffer_8201 (
        .din(new_Jinkela_wire_10304),
        .dout(new_Jinkela_wire_10305)
    );

    bfr new_Jinkela_buffer_8109 (
        .din(new_Jinkela_wire_10203),
        .dout(new_Jinkela_wire_10204)
    );

    bfr new_Jinkela_buffer_8149 (
        .din(new_Jinkela_wire_10250),
        .dout(new_Jinkela_wire_10251)
    );

    bfr new_Jinkela_buffer_8110 (
        .din(new_Jinkela_wire_10204),
        .dout(new_Jinkela_wire_10205)
    );

    bfr new_Jinkela_buffer_8111 (
        .din(new_Jinkela_wire_10205),
        .dout(new_Jinkela_wire_10206)
    );

    bfr new_Jinkela_buffer_8150 (
        .din(new_Jinkela_wire_10251),
        .dout(new_Jinkela_wire_10252)
    );

    bfr new_Jinkela_buffer_4516 (
        .din(new_Jinkela_wire_5379),
        .dout(new_Jinkela_wire_5380)
    );

    bfr new_Jinkela_buffer_6972 (
        .din(new_Jinkela_wire_8612),
        .dout(new_Jinkela_wire_8613)
    );

    bfr new_Jinkela_buffer_4485 (
        .din(new_Jinkela_wire_5339),
        .dout(new_Jinkela_wire_5340)
    );

    bfr new_Jinkela_buffer_7049 (
        .din(new_Jinkela_wire_8709),
        .dout(new_Jinkela_wire_8710)
    );

    bfr new_Jinkela_buffer_6999 (
        .din(new_Jinkela_wire_8642),
        .dout(new_Jinkela_wire_8643)
    );

    bfr new_Jinkela_buffer_6973 (
        .din(new_Jinkela_wire_8613),
        .dout(new_Jinkela_wire_8614)
    );

    bfr new_Jinkela_buffer_4486 (
        .din(new_Jinkela_wire_5340),
        .dout(new_Jinkela_wire_5341)
    );

    bfr new_Jinkela_buffer_7015 (
        .din(new_Jinkela_wire_8667),
        .dout(new_Jinkela_wire_8668)
    );

    bfr new_Jinkela_buffer_4517 (
        .din(new_Jinkela_wire_5380),
        .dout(new_Jinkela_wire_5381)
    );

    bfr new_Jinkela_buffer_6974 (
        .din(new_Jinkela_wire_8614),
        .dout(new_Jinkela_wire_8615)
    );

    bfr new_Jinkela_buffer_4487 (
        .din(new_Jinkela_wire_5341),
        .dout(new_Jinkela_wire_5342)
    );

    bfr new_Jinkela_buffer_7000 (
        .din(new_Jinkela_wire_8643),
        .dout(new_Jinkela_wire_8644)
    );

    bfr new_Jinkela_buffer_6975 (
        .din(new_Jinkela_wire_8615),
        .dout(new_Jinkela_wire_8616)
    );

    bfr new_Jinkela_buffer_4535 (
        .din(new_Jinkela_wire_5402),
        .dout(new_Jinkela_wire_5403)
    );

    bfr new_Jinkela_buffer_4518 (
        .din(new_Jinkela_wire_5381),
        .dout(new_Jinkela_wire_5382)
    );

    bfr new_Jinkela_buffer_6976 (
        .din(new_Jinkela_wire_8616),
        .dout(new_Jinkela_wire_8617)
    );

    spl3L new_Jinkela_splitter_328 (
        .a(n_0043_),
        .d(new_Jinkela_wire_5418),
        .b(new_Jinkela_wire_5419),
        .c(new_Jinkela_wire_5420)
    );

    bfr new_Jinkela_buffer_4519 (
        .din(new_Jinkela_wire_5382),
        .dout(new_Jinkela_wire_5383)
    );

    bfr new_Jinkela_buffer_7045 (
        .din(new_Jinkela_wire_8699),
        .dout(new_Jinkela_wire_8700)
    );

    bfr new_Jinkela_buffer_7001 (
        .din(new_Jinkela_wire_8644),
        .dout(new_Jinkela_wire_8645)
    );

    bfr new_Jinkela_buffer_4545 (
        .din(new_Jinkela_wire_5412),
        .dout(new_Jinkela_wire_5413)
    );

    bfr new_Jinkela_buffer_6977 (
        .din(new_Jinkela_wire_8617),
        .dout(new_Jinkela_wire_8618)
    );

    bfr new_Jinkela_buffer_4536 (
        .din(new_Jinkela_wire_5403),
        .dout(new_Jinkela_wire_5404)
    );

    bfr new_Jinkela_buffer_4520 (
        .din(new_Jinkela_wire_5383),
        .dout(new_Jinkela_wire_5384)
    );

    bfr new_Jinkela_buffer_7016 (
        .din(new_Jinkela_wire_8668),
        .dout(new_Jinkela_wire_8669)
    );

    bfr new_Jinkela_buffer_6978 (
        .din(new_Jinkela_wire_8618),
        .dout(new_Jinkela_wire_8619)
    );

    bfr new_Jinkela_buffer_4521 (
        .din(new_Jinkela_wire_5384),
        .dout(new_Jinkela_wire_5385)
    );

    bfr new_Jinkela_buffer_7002 (
        .din(new_Jinkela_wire_8645),
        .dout(new_Jinkela_wire_8646)
    );

    bfr new_Jinkela_buffer_4576 (
        .din(n_0665_),
        .dout(new_Jinkela_wire_5449)
    );

    bfr new_Jinkela_buffer_6979 (
        .din(new_Jinkela_wire_8619),
        .dout(new_Jinkela_wire_8620)
    );

    bfr new_Jinkela_buffer_4537 (
        .din(new_Jinkela_wire_5404),
        .dout(new_Jinkela_wire_5405)
    );

    bfr new_Jinkela_buffer_4522 (
        .din(new_Jinkela_wire_5385),
        .dout(new_Jinkela_wire_5386)
    );

    bfr new_Jinkela_buffer_6980 (
        .din(new_Jinkela_wire_8620),
        .dout(new_Jinkela_wire_8621)
    );

    bfr new_Jinkela_buffer_4523 (
        .din(new_Jinkela_wire_5386),
        .dout(new_Jinkela_wire_5387)
    );

    bfr new_Jinkela_buffer_7003 (
        .din(new_Jinkela_wire_8646),
        .dout(new_Jinkela_wire_8647)
    );

    bfr new_Jinkela_buffer_4546 (
        .din(new_Jinkela_wire_5413),
        .dout(new_Jinkela_wire_5414)
    );

    bfr new_Jinkela_buffer_6981 (
        .din(new_Jinkela_wire_8621),
        .dout(new_Jinkela_wire_8622)
    );

    bfr new_Jinkela_buffer_4538 (
        .din(new_Jinkela_wire_5405),
        .dout(new_Jinkela_wire_5406)
    );

    bfr new_Jinkela_buffer_4524 (
        .din(new_Jinkela_wire_5387),
        .dout(new_Jinkela_wire_5388)
    );

    bfr new_Jinkela_buffer_7017 (
        .din(new_Jinkela_wire_8669),
        .dout(new_Jinkela_wire_8670)
    );

    bfr new_Jinkela_buffer_6982 (
        .din(new_Jinkela_wire_8622),
        .dout(new_Jinkela_wire_8623)
    );

    bfr new_Jinkela_buffer_4525 (
        .din(new_Jinkela_wire_5388),
        .dout(new_Jinkela_wire_5389)
    );

    spl2 new_Jinkela_splitter_656 (
        .a(new_Jinkela_wire_8647),
        .b(new_Jinkela_wire_8648),
        .c(new_Jinkela_wire_8649)
    );

    spl2 new_Jinkela_splitter_331 (
        .a(n_0027_),
        .b(new_Jinkela_wire_5458),
        .c(new_Jinkela_wire_5459)
    );

    bfr new_Jinkela_buffer_4539 (
        .din(new_Jinkela_wire_5406),
        .dout(new_Jinkela_wire_5407)
    );

    bfr new_Jinkela_buffer_7018 (
        .din(new_Jinkela_wire_8670),
        .dout(new_Jinkela_wire_8671)
    );

    bfr new_Jinkela_buffer_4526 (
        .din(new_Jinkela_wire_5389),
        .dout(new_Jinkela_wire_5390)
    );

    bfr new_Jinkela_buffer_7048 (
        .din(n_0263_),
        .dout(new_Jinkela_wire_8709)
    );

    bfr new_Jinkela_buffer_7046 (
        .din(new_Jinkela_wire_8700),
        .dout(new_Jinkela_wire_8701)
    );

    bfr new_Jinkela_buffer_4548 (
        .din(new_Jinkela_wire_5420),
        .dout(new_Jinkela_wire_5421)
    );

    bfr new_Jinkela_buffer_4527 (
        .din(new_Jinkela_wire_5390),
        .dout(new_Jinkela_wire_5391)
    );

    spl2 new_Jinkela_splitter_665 (
        .a(n_0880_),
        .b(new_Jinkela_wire_8717),
        .c(new_Jinkela_wire_8718)
    );

    bfr new_Jinkela_buffer_7019 (
        .din(new_Jinkela_wire_8671),
        .dout(new_Jinkela_wire_8672)
    );

    spl2 new_Jinkela_splitter_327 (
        .a(new_Jinkela_wire_5414),
        .b(new_Jinkela_wire_5415),
        .c(new_Jinkela_wire_5416)
    );

    bfr new_Jinkela_buffer_4540 (
        .din(new_Jinkela_wire_5407),
        .dout(new_Jinkela_wire_5408)
    );

    spl2 new_Jinkela_splitter_664 (
        .a(n_1072_),
        .b(new_Jinkela_wire_8715),
        .c(new_Jinkela_wire_8716)
    );

    bfr new_Jinkela_buffer_7047 (
        .din(new_Jinkela_wire_8701),
        .dout(new_Jinkela_wire_8702)
    );

    bfr new_Jinkela_buffer_7020 (
        .din(new_Jinkela_wire_8672),
        .dout(new_Jinkela_wire_8673)
    );

    bfr new_Jinkela_buffer_4541 (
        .din(new_Jinkela_wire_5408),
        .dout(new_Jinkela_wire_5409)
    );

    bfr new_Jinkela_buffer_7021 (
        .din(new_Jinkela_wire_8673),
        .dout(new_Jinkela_wire_8674)
    );

    bfr new_Jinkela_buffer_4581 (
        .din(new_Jinkela_wire_5459),
        .dout(new_Jinkela_wire_5460)
    );

    bfr new_Jinkela_buffer_4542 (
        .din(new_Jinkela_wire_5409),
        .dout(new_Jinkela_wire_5410)
    );

    spl4L new_Jinkela_splitter_667 (
        .a(n_1069_),
        .d(new_Jinkela_wire_8749),
        .b(new_Jinkela_wire_8750),
        .e(new_Jinkela_wire_8751),
        .c(new_Jinkela_wire_8752)
    );

    spl2 new_Jinkela_splitter_661 (
        .a(new_Jinkela_wire_8702),
        .b(new_Jinkela_wire_8703),
        .c(new_Jinkela_wire_8704)
    );

    bfr new_Jinkela_buffer_7022 (
        .din(new_Jinkela_wire_8674),
        .dout(new_Jinkela_wire_8675)
    );

    bfr new_Jinkela_buffer_4549 (
        .din(new_Jinkela_wire_5421),
        .dout(new_Jinkela_wire_5422)
    );

    bfr new_Jinkela_buffer_4543 (
        .din(new_Jinkela_wire_5410),
        .dout(new_Jinkela_wire_5411)
    );

    bfr new_Jinkela_buffer_7023 (
        .din(new_Jinkela_wire_8675),
        .dout(new_Jinkela_wire_8676)
    );

    spl2 new_Jinkela_splitter_329 (
        .a(new_Jinkela_wire_5449),
        .b(new_Jinkela_wire_5450),
        .c(new_Jinkela_wire_5451)
    );

    bfr new_Jinkela_buffer_4550 (
        .din(new_Jinkela_wire_5422),
        .dout(new_Jinkela_wire_5423)
    );

    bfr new_Jinkela_buffer_7024 (
        .din(new_Jinkela_wire_8676),
        .dout(new_Jinkela_wire_8677)
    );

    bfr new_Jinkela_buffer_4577 (
        .din(new_Jinkela_wire_5451),
        .dout(new_Jinkela_wire_5452)
    );

    bfr new_Jinkela_buffer_4621 (
        .din(n_0310_),
        .dout(new_Jinkela_wire_5500)
    );

    bfr new_Jinkela_buffer_7050 (
        .din(new_Jinkela_wire_8710),
        .dout(new_Jinkela_wire_8711)
    );

    bfr new_Jinkela_buffer_4551 (
        .din(new_Jinkela_wire_5423),
        .dout(new_Jinkela_wire_5424)
    );

    bfr new_Jinkela_buffer_7025 (
        .din(new_Jinkela_wire_8677),
        .dout(new_Jinkela_wire_8678)
    );

    bfr new_Jinkela_buffer_7051 (
        .din(new_Jinkela_wire_8711),
        .dout(new_Jinkela_wire_8712)
    );

    bfr new_Jinkela_buffer_4552 (
        .din(new_Jinkela_wire_5424),
        .dout(new_Jinkela_wire_5425)
    );

    bfr new_Jinkela_buffer_7026 (
        .din(new_Jinkela_wire_8678),
        .dout(new_Jinkela_wire_8679)
    );

    bfr new_Jinkela_buffer_4623 (
        .din(n_0867_),
        .dout(new_Jinkela_wire_5502)
    );

    bfr new_Jinkela_buffer_7054 (
        .din(new_net_2523),
        .dout(new_Jinkela_wire_8719)
    );

    bfr new_Jinkela_buffer_4553 (
        .din(new_Jinkela_wire_5425),
        .dout(new_Jinkela_wire_5426)
    );

    spl2 new_Jinkela_splitter_666 (
        .a(n_0618_),
        .b(new_Jinkela_wire_8747),
        .c(new_Jinkela_wire_8748)
    );

    bfr new_Jinkela_buffer_2613 (
        .din(new_Jinkela_wire_3018),
        .dout(new_Jinkela_wire_3019)
    );

    bfr new_Jinkela_buffer_2614 (
        .din(new_Jinkela_wire_3019),
        .dout(new_Jinkela_wire_3020)
    );

    bfr new_Jinkela_buffer_2615 (
        .din(new_Jinkela_wire_3020),
        .dout(new_Jinkela_wire_3021)
    );

    bfr new_Jinkela_buffer_2660 (
        .din(new_Jinkela_wire_3069),
        .dout(new_Jinkela_wire_3070)
    );

    bfr new_Jinkela_buffer_1262 (
        .din(new_Jinkela_wire_1582),
        .dout(new_Jinkela_wire_1583)
    );

    bfr new_Jinkela_buffer_724 (
        .din(new_Jinkela_wire_780),
        .dout(new_Jinkela_wire_781)
    );

    bfr new_Jinkela_buffer_6219 (
        .din(new_Jinkela_wire_7592),
        .dout(new_Jinkela_wire_7593)
    );

    bfr new_Jinkela_buffer_6169 (
        .din(new_Jinkela_wire_7534),
        .dout(new_Jinkela_wire_7535)
    );

    bfr new_Jinkela_buffer_1372 (
        .din(new_Jinkela_wire_1697),
        .dout(new_Jinkela_wire_1698)
    );

    bfr new_Jinkela_buffer_616 (
        .din(new_Jinkela_wire_664),
        .dout(new_Jinkela_wire_665)
    );

    bfr new_Jinkela_buffer_6187 (
        .din(new_Jinkela_wire_7560),
        .dout(new_Jinkela_wire_7561)
    );

    bfr new_Jinkela_buffer_1263 (
        .din(new_Jinkela_wire_1583),
        .dout(new_Jinkela_wire_1584)
    );

    bfr new_Jinkela_buffer_660 (
        .din(new_Jinkela_wire_712),
        .dout(new_Jinkela_wire_713)
    );

    bfr new_Jinkela_buffer_6170 (
        .din(new_Jinkela_wire_7535),
        .dout(new_Jinkela_wire_7536)
    );

    bfr new_Jinkela_buffer_1309 (
        .din(new_Jinkela_wire_1634),
        .dout(new_Jinkela_wire_1635)
    );

    bfr new_Jinkela_buffer_617 (
        .din(new_Jinkela_wire_665),
        .dout(new_Jinkela_wire_666)
    );

    bfr new_Jinkela_buffer_1264 (
        .din(new_Jinkela_wire_1584),
        .dout(new_Jinkela_wire_1585)
    );

    bfr new_Jinkela_buffer_722 (
        .din(new_Jinkela_wire_778),
        .dout(new_Jinkela_wire_779)
    );

    bfr new_Jinkela_buffer_6171 (
        .din(new_Jinkela_wire_7536),
        .dout(new_Jinkela_wire_7537)
    );

    bfr new_Jinkela_buffer_1375 (
        .din(new_Jinkela_wire_1702),
        .dout(new_Jinkela_wire_1703)
    );

    bfr new_Jinkela_buffer_618 (
        .din(new_Jinkela_wire_666),
        .dout(new_Jinkela_wire_667)
    );

    bfr new_Jinkela_buffer_1378 (
        .din(N254),
        .dout(new_Jinkela_wire_1706)
    );

    bfr new_Jinkela_buffer_6188 (
        .din(new_Jinkela_wire_7561),
        .dout(new_Jinkela_wire_7562)
    );

    bfr new_Jinkela_buffer_1265 (
        .din(new_Jinkela_wire_1585),
        .dout(new_Jinkela_wire_1586)
    );

    bfr new_Jinkela_buffer_661 (
        .din(new_Jinkela_wire_713),
        .dout(new_Jinkela_wire_714)
    );

    bfr new_Jinkela_buffer_6172 (
        .din(new_Jinkela_wire_7537),
        .dout(new_Jinkela_wire_7538)
    );

    bfr new_Jinkela_buffer_1310 (
        .din(new_Jinkela_wire_1635),
        .dout(new_Jinkela_wire_1636)
    );

    bfr new_Jinkela_buffer_619 (
        .din(new_Jinkela_wire_667),
        .dout(new_Jinkela_wire_668)
    );

    bfr new_Jinkela_buffer_6306 (
        .din(new_Jinkela_wire_7687),
        .dout(new_Jinkela_wire_7688)
    );

    bfr new_Jinkela_buffer_1266 (
        .din(new_Jinkela_wire_1586),
        .dout(new_Jinkela_wire_1587)
    );

    bfr new_Jinkela_buffer_731 (
        .din(N208),
        .dout(new_Jinkela_wire_788)
    );

    bfr new_Jinkela_buffer_6220 (
        .din(new_Jinkela_wire_7593),
        .dout(new_Jinkela_wire_7594)
    );

    spl2 new_Jinkela_splitter_537 (
        .a(new_Jinkela_wire_7538),
        .b(new_Jinkela_wire_7539),
        .c(new_Jinkela_wire_7540)
    );

    bfr new_Jinkela_buffer_620 (
        .din(new_Jinkela_wire_668),
        .dout(new_Jinkela_wire_669)
    );

    bfr new_Jinkela_buffer_1267 (
        .din(new_Jinkela_wire_1587),
        .dout(new_Jinkela_wire_1588)
    );

    bfr new_Jinkela_buffer_662 (
        .din(new_Jinkela_wire_714),
        .dout(new_Jinkela_wire_715)
    );

    bfr new_Jinkela_buffer_6278 (
        .din(new_Jinkela_wire_7655),
        .dout(new_Jinkela_wire_7656)
    );

    bfr new_Jinkela_buffer_6189 (
        .din(new_Jinkela_wire_7562),
        .dout(new_Jinkela_wire_7563)
    );

    bfr new_Jinkela_buffer_1311 (
        .din(new_Jinkela_wire_1636),
        .dout(new_Jinkela_wire_1637)
    );

    bfr new_Jinkela_buffer_621 (
        .din(new_Jinkela_wire_669),
        .dout(new_Jinkela_wire_670)
    );

    bfr new_Jinkela_buffer_6190 (
        .din(new_Jinkela_wire_7563),
        .dout(new_Jinkela_wire_7564)
    );

    bfr new_Jinkela_buffer_1268 (
        .din(new_Jinkela_wire_1588),
        .dout(new_Jinkela_wire_1589)
    );

    bfr new_Jinkela_buffer_725 (
        .din(new_Jinkela_wire_781),
        .dout(new_Jinkela_wire_782)
    );

    bfr new_Jinkela_buffer_622 (
        .din(new_Jinkela_wire_670),
        .dout(new_Jinkela_wire_671)
    );

    bfr new_Jinkela_buffer_6221 (
        .din(new_Jinkela_wire_7594),
        .dout(new_Jinkela_wire_7595)
    );

    bfr new_Jinkela_buffer_6191 (
        .din(new_Jinkela_wire_7564),
        .dout(new_Jinkela_wire_7565)
    );

    bfr new_Jinkela_buffer_1269 (
        .din(new_Jinkela_wire_1589),
        .dout(new_Jinkela_wire_1590)
    );

    bfr new_Jinkela_buffer_663 (
        .din(new_Jinkela_wire_715),
        .dout(new_Jinkela_wire_716)
    );

    bfr new_Jinkela_buffer_1312 (
        .din(new_Jinkela_wire_1637),
        .dout(new_Jinkela_wire_1638)
    );

    bfr new_Jinkela_buffer_623 (
        .din(new_Jinkela_wire_671),
        .dout(new_Jinkela_wire_672)
    );

    spl2 new_Jinkela_splitter_545 (
        .a(n_1332_),
        .b(new_Jinkela_wire_7730),
        .c(new_Jinkela_wire_7731)
    );

    bfr new_Jinkela_buffer_6192 (
        .din(new_Jinkela_wire_7565),
        .dout(new_Jinkela_wire_7566)
    );

    bfr new_Jinkela_buffer_1270 (
        .din(new_Jinkela_wire_1590),
        .dout(new_Jinkela_wire_1591)
    );

    bfr new_Jinkela_buffer_728 (
        .din(new_Jinkela_wire_784),
        .dout(new_Jinkela_wire_785)
    );

    bfr new_Jinkela_buffer_2618 (
        .din(new_Jinkela_wire_3023),
        .dout(new_Jinkela_wire_3024)
    );

    bfr new_Jinkela_buffer_1376 (
        .din(new_Jinkela_wire_1703),
        .dout(new_Jinkela_wire_1704)
    );

    bfr new_Jinkela_buffer_624 (
        .din(new_Jinkela_wire_672),
        .dout(new_Jinkela_wire_673)
    );

    bfr new_Jinkela_buffer_6222 (
        .din(new_Jinkela_wire_7595),
        .dout(new_Jinkela_wire_7596)
    );

    bfr new_Jinkela_buffer_6193 (
        .din(new_Jinkela_wire_7566),
        .dout(new_Jinkela_wire_7567)
    );

    bfr new_Jinkela_buffer_1271 (
        .din(new_Jinkela_wire_1591),
        .dout(new_Jinkela_wire_1592)
    );

    bfr new_Jinkela_buffer_664 (
        .din(new_Jinkela_wire_716),
        .dout(new_Jinkela_wire_717)
    );

    bfr new_Jinkela_buffer_1313 (
        .din(new_Jinkela_wire_1638),
        .dout(new_Jinkela_wire_1639)
    );

    bfr new_Jinkela_buffer_625 (
        .din(new_Jinkela_wire_673),
        .dout(new_Jinkela_wire_674)
    );

    bfr new_Jinkela_buffer_6279 (
        .din(new_Jinkela_wire_7656),
        .dout(new_Jinkela_wire_7657)
    );

    bfr new_Jinkela_buffer_6194 (
        .din(new_Jinkela_wire_7567),
        .dout(new_Jinkela_wire_7568)
    );

    bfr new_Jinkela_buffer_1272 (
        .din(new_Jinkela_wire_1592),
        .dout(new_Jinkela_wire_1593)
    );

    bfr new_Jinkela_buffer_726 (
        .din(new_Jinkela_wire_782),
        .dout(new_Jinkela_wire_783)
    );

    bfr new_Jinkela_buffer_1379 (
        .din(new_Jinkela_wire_1706),
        .dout(new_Jinkela_wire_1707)
    );

    bfr new_Jinkela_buffer_626 (
        .din(new_Jinkela_wire_674),
        .dout(new_Jinkela_wire_675)
    );

    bfr new_Jinkela_buffer_6223 (
        .din(new_Jinkela_wire_7596),
        .dout(new_Jinkela_wire_7597)
    );

    bfr new_Jinkela_buffer_6195 (
        .din(new_Jinkela_wire_7568),
        .dout(new_Jinkela_wire_7569)
    );

    bfr new_Jinkela_buffer_1273 (
        .din(new_Jinkela_wire_1593),
        .dout(new_Jinkela_wire_1594)
    );

    bfr new_Jinkela_buffer_665 (
        .din(new_Jinkela_wire_717),
        .dout(new_Jinkela_wire_718)
    );

    bfr new_Jinkela_buffer_1314 (
        .din(new_Jinkela_wire_1639),
        .dout(new_Jinkela_wire_1640)
    );

    bfr new_Jinkela_buffer_627 (
        .din(new_Jinkela_wire_675),
        .dout(new_Jinkela_wire_676)
    );

    bfr new_Jinkela_buffer_6350 (
        .din(n_0514_),
        .dout(new_Jinkela_wire_7736)
    );

    bfr new_Jinkela_buffer_6196 (
        .din(new_Jinkela_wire_7569),
        .dout(new_Jinkela_wire_7570)
    );

    bfr new_Jinkela_buffer_1274 (
        .din(new_Jinkela_wire_1594),
        .dout(new_Jinkela_wire_1595)
    );

    bfr new_Jinkela_buffer_735 (
        .din(N155),
        .dout(new_Jinkela_wire_792)
    );

    bfr new_Jinkela_buffer_6345 (
        .din(new_Jinkela_wire_7728),
        .dout(new_Jinkela_wire_7729)
    );

    bfr new_Jinkela_buffer_1377 (
        .din(new_Jinkela_wire_1704),
        .dout(new_Jinkela_wire_1705)
    );

    bfr new_Jinkela_buffer_628 (
        .din(new_Jinkela_wire_676),
        .dout(new_Jinkela_wire_677)
    );

    bfr new_Jinkela_buffer_6224 (
        .din(new_Jinkela_wire_7597),
        .dout(new_Jinkela_wire_7598)
    );

    bfr new_Jinkela_buffer_6197 (
        .din(new_Jinkela_wire_7570),
        .dout(new_Jinkela_wire_7571)
    );

    bfr new_Jinkela_buffer_1275 (
        .din(new_Jinkela_wire_1595),
        .dout(new_Jinkela_wire_1596)
    );

    bfr new_Jinkela_buffer_666 (
        .din(new_Jinkela_wire_718),
        .dout(new_Jinkela_wire_719)
    );

    bfr new_Jinkela_buffer_2619 (
        .din(new_Jinkela_wire_3024),
        .dout(new_Jinkela_wire_3025)
    );

    bfr new_Jinkela_buffer_1315 (
        .din(new_Jinkela_wire_1640),
        .dout(new_Jinkela_wire_1641)
    );

    bfr new_Jinkela_buffer_629 (
        .din(new_Jinkela_wire_677),
        .dout(new_Jinkela_wire_678)
    );

    bfr new_Jinkela_buffer_6280 (
        .din(new_Jinkela_wire_7657),
        .dout(new_Jinkela_wire_7658)
    );

    bfr new_Jinkela_buffer_6198 (
        .din(new_Jinkela_wire_7571),
        .dout(new_Jinkela_wire_7572)
    );

    bfr new_Jinkela_buffer_1276 (
        .din(new_Jinkela_wire_1596),
        .dout(new_Jinkela_wire_1597)
    );

    bfr new_Jinkela_buffer_729 (
        .din(new_Jinkela_wire_785),
        .dout(new_Jinkela_wire_786)
    );

    bfr new_Jinkela_buffer_667 (
        .din(new_Jinkela_wire_719),
        .dout(new_Jinkela_wire_720)
    );

    bfr new_Jinkela_buffer_1446 (
        .din(N53),
        .dout(new_Jinkela_wire_1779)
    );

    bfr new_Jinkela_buffer_6225 (
        .din(new_Jinkela_wire_7598),
        .dout(new_Jinkela_wire_7599)
    );

    bfr new_Jinkela_buffer_6199 (
        .din(new_Jinkela_wire_7572),
        .dout(new_Jinkela_wire_7573)
    );

    bfr new_Jinkela_buffer_1277 (
        .din(new_Jinkela_wire_1597),
        .dout(new_Jinkela_wire_1598)
    );

    bfr new_Jinkela_buffer_732 (
        .din(new_Jinkela_wire_788),
        .dout(new_Jinkela_wire_789)
    );

    bfr new_Jinkela_buffer_1316 (
        .din(new_Jinkela_wire_1641),
        .dout(new_Jinkela_wire_1642)
    );

    bfr new_Jinkela_buffer_668 (
        .din(new_Jinkela_wire_720),
        .dout(new_Jinkela_wire_721)
    );

    bfr new_Jinkela_buffer_6307 (
        .din(new_Jinkela_wire_7688),
        .dout(new_Jinkela_wire_7689)
    );

    bfr new_Jinkela_buffer_6200 (
        .din(new_Jinkela_wire_7573),
        .dout(new_Jinkela_wire_7574)
    );

    bfr new_Jinkela_buffer_1278 (
        .din(new_Jinkela_wire_1598),
        .dout(new_Jinkela_wire_1599)
    );

    bfr new_Jinkela_buffer_730 (
        .din(new_Jinkela_wire_786),
        .dout(new_Jinkela_wire_787)
    );

    bfr new_Jinkela_buffer_1380 (
        .din(new_Jinkela_wire_1707),
        .dout(new_Jinkela_wire_1708)
    );

    bfr new_Jinkela_buffer_669 (
        .din(new_Jinkela_wire_721),
        .dout(new_Jinkela_wire_722)
    );

    bfr new_Jinkela_buffer_6226 (
        .din(new_Jinkela_wire_7599),
        .dout(new_Jinkela_wire_7600)
    );

    bfr new_Jinkela_buffer_6201 (
        .din(new_Jinkela_wire_7574),
        .dout(new_Jinkela_wire_7575)
    );

    bfr new_Jinkela_buffer_1279 (
        .din(new_Jinkela_wire_1599),
        .dout(new_Jinkela_wire_1600)
    );

    bfr new_Jinkela_buffer_739 (
        .din(N94),
        .dout(new_Jinkela_wire_796)
    );

    bfr new_Jinkela_buffer_1317 (
        .din(new_Jinkela_wire_1642),
        .dout(new_Jinkela_wire_1643)
    );

    bfr new_Jinkela_buffer_670 (
        .din(new_Jinkela_wire_722),
        .dout(new_Jinkela_wire_723)
    );

    bfr new_Jinkela_buffer_6281 (
        .din(new_Jinkela_wire_7658),
        .dout(new_Jinkela_wire_7659)
    );

    bfr new_Jinkela_buffer_6202 (
        .din(new_Jinkela_wire_7575),
        .dout(new_Jinkela_wire_7576)
    );

    bfr new_Jinkela_buffer_1280 (
        .din(new_Jinkela_wire_1600),
        .dout(new_Jinkela_wire_1601)
    );

    bfr new_Jinkela_buffer_733 (
        .din(new_Jinkela_wire_789),
        .dout(new_Jinkela_wire_790)
    );

    bfr new_Jinkela_buffer_2620 (
        .din(new_Jinkela_wire_3025),
        .dout(new_Jinkela_wire_3026)
    );

    bfr new_Jinkela_buffer_1443 (
        .din(new_Jinkela_wire_1775),
        .dout(new_Jinkela_wire_1776)
    );

    bfr new_Jinkela_buffer_671 (
        .din(new_Jinkela_wire_723),
        .dout(new_Jinkela_wire_724)
    );

    bfr new_Jinkela_buffer_1442 (
        .din(N193),
        .dout(new_Jinkela_wire_1775)
    );

    bfr new_Jinkela_buffer_6227 (
        .din(new_Jinkela_wire_7600),
        .dout(new_Jinkela_wire_7601)
    );

    bfr new_Jinkela_buffer_6203 (
        .din(new_Jinkela_wire_7576),
        .dout(new_Jinkela_wire_7577)
    );

    bfr new_Jinkela_buffer_1281 (
        .din(new_Jinkela_wire_1601),
        .dout(new_Jinkela_wire_1602)
    );

    bfr new_Jinkela_buffer_736 (
        .din(new_Jinkela_wire_792),
        .dout(new_Jinkela_wire_793)
    );

    bfr new_Jinkela_buffer_1318 (
        .din(new_Jinkela_wire_1643),
        .dout(new_Jinkela_wire_1644)
    );

    bfr new_Jinkela_buffer_672 (
        .din(new_Jinkela_wire_724),
        .dout(new_Jinkela_wire_725)
    );

    bfr new_Jinkela_buffer_6204 (
        .din(new_Jinkela_wire_7577),
        .dout(new_Jinkela_wire_7578)
    );

    bfr new_Jinkela_buffer_1282 (
        .din(new_Jinkela_wire_1602),
        .dout(new_Jinkela_wire_1603)
    );

    bfr new_Jinkela_buffer_734 (
        .din(new_Jinkela_wire_790),
        .dout(new_Jinkela_wire_791)
    );

    bfr new_Jinkela_buffer_6228 (
        .din(new_Jinkela_wire_7601),
        .dout(new_Jinkela_wire_7602)
    );

endmodule
