module c3540(G25,G47,G30,G50,G27,G3,G31,G19,G9,G13,G39,G34,G8,G46,G14,G18,G32,G42,G11,G48,G22,G4,G17,G35,G23,G21,G36,G41,G5,G38,G26,G7,G1,G28,G6,G24,G20,G43,G44,G12,G40,G10,G29,G16,G33,G37,G45,G49,G15,G2);
    wire new_Jinkela_wire_1621;
    wire new_Jinkela_wire_2646;
    wire new_Jinkela_wire_621;
    wire new_Jinkela_wire_338;
    wire new_Jinkela_wire_1956;
    wire new_Jinkela_wire_839;
    wire new_Jinkela_wire_1714;
    wire new_Jinkela_wire_1061;
    wire new_Jinkela_wire_2333;
    wire _0257_;
    wire new_Jinkela_wire_234;
    wire new_Jinkela_wire_37;
    wire new_Jinkela_wire_1211;
    wire new_Jinkela_wire_541;
    wire new_Jinkela_wire_2608;
    wire new_Jinkela_wire_2947;
    wire new_Jinkela_wire_3086;
    wire _0109_;
    wire _0205_;
    wire new_Jinkela_wire_1183;
    wire new_Jinkela_wire_436;
    wire new_Jinkela_wire_77;
    wire new_Jinkela_wire_3286;
    wire new_Jinkela_wire_2184;
    wire _0178_;
    wire new_Jinkela_wire_1008;
    wire new_Jinkela_wire_2629;
    wire new_Jinkela_wire_1187;
    wire new_Jinkela_wire_116;
    wire new_Jinkela_wire_3295;
    wire new_Jinkela_wire_2494;
    wire new_Jinkela_wire_3158;
    wire new_Jinkela_wire_905;
    wire new_Jinkela_wire_760;
    wire new_Jinkela_wire_2221;
    wire _0405_;
    wire new_Jinkela_wire_1695;
    wire new_Jinkela_wire_2672;
    wire new_Jinkela_wire_1507;
    wire new_Jinkela_wire_2702;
    wire new_Jinkela_wire_2680;
    wire new_Jinkela_wire_4;
    wire new_Jinkela_wire_470;
    wire _0605_;
    wire new_Jinkela_wire_1220;
    wire new_Jinkela_wire_530;
    wire new_Jinkela_wire_419;
    wire _0253_;
    wire new_Jinkela_wire_1645;
    wire new_Jinkela_wire_2300;
    wire _0242_;
    wire new_Jinkela_wire_1655;
    wire new_Jinkela_wire_2175;
    wire new_Jinkela_wire_2801;
    wire new_Jinkela_wire_3077;
    wire new_Jinkela_wire_955;
    wire new_Jinkela_wire_14;
    wire new_Jinkela_wire_654;
    wire new_Jinkela_wire_2634;
    wire new_Jinkela_wire_3114;
    wire new_Jinkela_wire_850;
    wire new_Jinkela_wire_1567;
    wire _0333_;
    wire new_Jinkela_wire_45;
    wire new_Jinkela_wire_1736;
    wire new_Jinkela_wire_2633;
    wire _0527_;
    wire new_Jinkela_wire_1962;
    wire _0095_;
    wire _0571_;
    wire new_Jinkela_wire_1088;
    wire new_Jinkela_wire_709;
    wire new_Jinkela_wire_762;
    wire new_Jinkela_wire_2186;
    wire _0536_;
    wire new_Jinkela_wire_2438;
    wire new_Jinkela_wire_1678;
    wire new_Jinkela_wire_1555;
    wire _0681_;
    wire _0583_;
    wire new_Jinkela_wire_2986;
    wire new_Jinkela_wire_1089;
    wire new_Jinkela_wire_2290;
    wire new_Jinkela_wire_2682;
    wire _0685_;
    wire _0121_;
    wire new_Jinkela_wire_2032;
    wire new_Jinkela_wire_1791;
    wire new_Jinkela_wire_524;
    wire _0290_;
    wire new_Jinkela_wire_3180;
    wire _0044_;
    wire new_Jinkela_wire_2984;
    wire new_Jinkela_wire_632;
    wire new_Jinkela_wire_2211;
    wire _0190_;
    wire new_Jinkela_wire_2442;
    wire new_Jinkela_wire_1981;
    wire new_Jinkela_wire_2408;
    wire _0162_;
    wire new_Jinkela_wire_2164;
    wire new_Jinkela_wire_781;
    wire new_Jinkela_wire_151;
    wire new_Jinkela_wire_1828;
    wire new_Jinkela_wire_1097;
    wire new_Jinkela_wire_611;
    wire new_Jinkela_wire_3188;
    wire new_Jinkela_wire_1819;
    wire new_Jinkela_wire_3045;
    wire _0614_;
    wire _0293_;
    wire new_Jinkela_wire_539;
    wire new_Jinkela_wire_986;
    wire new_Jinkela_wire_3261;
    wire new_Jinkela_wire_738;
    wire new_Jinkela_wire_423;
    wire new_Jinkela_wire_1232;
    wire _0755_;
    wire new_Jinkela_wire_793;
    wire _0072_;
    wire _0395_;
    wire _0676_;
    wire new_Jinkela_wire_2039;
    wire new_Jinkela_wire_1532;
    wire new_Jinkela_wire_1110;
    wire new_Jinkela_wire_2339;
    wire new_Jinkela_wire_31;
    wire new_Jinkela_wire_3297;
    wire new_Jinkela_wire_1948;
    wire _0092_;
    wire _0345_;
    wire new_Jinkela_wire_1995;
    wire new_Jinkela_wire_2141;
    wire new_Jinkela_wire_2722;
    wire new_Jinkela_wire_2497;
    wire new_Jinkela_wire_1672;
    wire new_Jinkela_wire_2054;
    wire new_Jinkela_wire_2108;
    wire new_net_1481;
    wire _0415_;
    wire new_Jinkela_wire_18;
    wire new_Jinkela_wire_677;
    wire new_Jinkela_wire_461;
    wire new_Jinkela_wire_1776;
    wire new_Jinkela_wire_853;
    wire new_Jinkela_wire_1950;
    wire new_Jinkela_wire_1733;
    wire new_Jinkela_wire_2085;
    wire _0754_;
    wire new_Jinkela_wire_1909;
    wire new_Jinkela_wire_2907;
    wire new_Jinkela_wire_1949;
    wire _0557_;
    wire new_Jinkela_wire_468;
    wire new_Jinkela_wire_2152;
    wire new_Jinkela_wire_157;
    wire new_Jinkela_wire_3139;
    wire new_Jinkela_wire_1018;
    wire new_Jinkela_wire_432;
    wire _0339_;
    wire _0456_;
    wire _0600_;
    wire new_Jinkela_wire_2921;
    wire new_Jinkela_wire_1556;
    wire new_Jinkela_wire_2909;
    wire new_Jinkela_wire_3309;
    wire new_Jinkela_wire_2307;
    wire new_Jinkela_wire_1345;
    wire new_Jinkela_wire_2312;
    wire new_Jinkela_wire_2717;
    wire new_Jinkela_wire_1186;
    wire new_Jinkela_wire_686;
    wire new_Jinkela_wire_1894;
    wire new_Jinkela_wire_1297;
    wire new_Jinkela_wire_1474;
    wire new_Jinkela_wire_1533;
    wire new_Jinkela_wire_3135;
    wire new_Jinkela_wire_3307;
    wire new_Jinkela_wire_2761;
    wire _0734_;
    wire _0678_;
    wire new_Jinkela_wire_610;
    wire new_Jinkela_wire_1338;
    wire new_Jinkela_wire_545;
    wire new_Jinkela_wire_2506;
    wire new_Jinkela_wire_661;
    wire new_Jinkela_wire_966;
    wire _0228_;
    wire new_Jinkela_wire_1479;
    wire new_Jinkela_wire_2075;
    wire new_Jinkela_wire_3207;
    wire _0312_;
    wire new_Jinkela_wire_3257;
    wire new_Jinkela_wire_1332;
    wire new_Jinkela_wire_958;
    wire new_Jinkela_wire_154;
    wire _0107_;
    wire new_Jinkela_wire_442;
    wire new_Jinkela_wire_629;
    wire new_Jinkela_wire_495;
    wire new_Jinkela_wire_2034;
    wire new_Jinkela_wire_1007;
    wire _0512_;
    wire new_Jinkela_wire_502;
    wire new_Jinkela_wire_2264;
    wire new_Jinkela_wire_1830;
    wire new_Jinkela_wire_134;
    wire _0428_;
    wire new_Jinkela_wire_148;
    wire new_Jinkela_wire_1149;
    wire new_Jinkela_wire_114;
    wire _0038_;
    wire new_Jinkela_wire_2177;
    wire new_Jinkela_wire_2235;
    wire new_Jinkela_wire_2547;
    wire new_Jinkela_wire_2055;
    wire new_Jinkela_wire_2397;
    wire new_Jinkela_wire_135;
    wire new_Jinkela_wire_1397;
    wire _0464_;
    wire new_Jinkela_wire_124;
    wire _0660_;
    wire new_Jinkela_wire_101;
    wire new_Jinkela_wire_1625;
    wire _0201_;
    wire new_Jinkela_wire_2410;
    wire new_Jinkela_wire_1697;
    wire _0629_;
    wire new_Jinkela_wire_585;
    wire new_Jinkela_wire_2481;
    wire new_Jinkela_wire_1738;
    wire new_Jinkela_wire_277;
    wire _0299_;
    wire new_Jinkela_wire_2550;
    wire new_Jinkela_wire_2860;
    wire _0354_;
    wire new_Jinkela_wire_1368;
    wire new_Jinkela_wire_3196;
    wire new_Jinkela_wire_1364;
    wire new_Jinkela_wire_491;
    wire new_Jinkela_wire_2588;
    wire new_Jinkela_wire_2248;
    wire new_Jinkela_wire_1017;
    wire new_Jinkela_wire_649;
    wire new_Jinkela_wire_1650;
    wire new_Jinkela_wire_2600;
    wire new_Jinkela_wire_670;
    wire new_Jinkela_wire_161;
    wire new_Jinkela_wire_1190;
    wire new_Jinkela_wire_34;
    wire _0429_;
    wire new_Jinkela_wire_1319;
    wire new_Jinkela_wire_2779;
    wire new_Jinkela_wire_1925;
    wire new_Jinkela_wire_2580;
    wire _0383_;
    wire new_Jinkela_wire_982;
    wire new_Jinkela_wire_1189;
    wire new_Jinkela_wire_1315;
    wire new_Jinkela_wire_247;
    wire new_Jinkela_wire_3271;
    wire new_Jinkela_wire_2526;
    wire new_Jinkela_wire_2068;
    wire _0402_;
    wire new_Jinkela_wire_582;
    wire new_Jinkela_wire_39;
    wire new_Jinkela_wire_1928;
    wire new_Jinkela_wire_657;
    wire _0142_;
    wire new_Jinkela_wire_3106;
    wire new_Jinkela_wire_1227;
    wire new_Jinkela_wire_2127;
    wire new_Jinkela_wire_69;
    wire new_Jinkela_wire_1699;
    wire new_Jinkela_wire_110;
    wire new_Jinkela_wire_1122;
    wire new_Jinkela_wire_2544;
    wire new_Jinkela_wire_3098;
    wire new_Jinkela_wire_2697;
    wire _0249_;
    wire new_Jinkela_wire_2698;
    wire new_Jinkela_wire_2231;
    wire new_Jinkela_wire_1762;
    wire new_Jinkela_wire_925;
    wire new_Jinkela_wire_98;
    wire new_Jinkela_wire_2082;
    wire new_Jinkela_wire_1970;
    wire new_Jinkela_wire_609;
    wire new_Jinkela_wire_2813;
    wire new_Jinkela_wire_2884;
    wire new_Jinkela_wire_2374;
    wire new_Jinkela_wire_984;
    wire new_Jinkela_wire_2181;
    wire new_Jinkela_wire_1282;
    wire new_Jinkela_wire_918;
    wire new_Jinkela_wire_3224;
    wire new_Jinkela_wire_1549;
    wire new_Jinkela_wire_2450;
    wire new_Jinkela_wire_747;
    wire new_Jinkela_wire_3242;
    wire new_Jinkela_wire_1912;
    wire new_Jinkela_wire_1947;
    wire new_Jinkela_wire_1420;
    wire _0470_;
    wire new_Jinkela_wire_2893;
    wire new_Jinkela_wire_3277;
    wire new_Jinkela_wire_2100;
    wire new_Jinkela_wire_1328;
    wire new_Jinkela_wire_1863;
    wire new_Jinkela_wire_224;
    wire _0327_;
    wire new_Jinkela_wire_1945;
    wire new_Jinkela_wire_406;
    wire new_Jinkela_wire_763;
    wire new_Jinkela_wire_2216;
    wire new_Jinkela_wire_2019;
    wire new_Jinkela_wire_1073;
    wire new_Jinkela_wire_464;
    wire new_Jinkela_wire_2518;
    wire new_Jinkela_wire_477;
    wire _0133_;
    wire new_Jinkela_wire_3117;
    wire new_Jinkela_wire_3179;
    wire new_Jinkela_wire_1418;
    wire new_Jinkela_wire_2687;
    wire new_Jinkela_wire_2625;
    wire new_Jinkela_wire_932;
    wire new_Jinkela_wire_250;
    wire new_Jinkela_wire_2218;
    wire new_Jinkela_wire_2236;
    wire new_Jinkela_wire_1323;
    wire new_Jinkela_wire_1582;
    wire new_Jinkela_wire_1045;
    wire new_Jinkela_wire_1812;
    wire new_Jinkela_wire_716;
    wire new_Jinkela_wire_325;
    wire new_Jinkela_wire_936;
    wire new_Jinkela_wire_3234;
    wire new_Jinkela_wire_100;
    wire new_Jinkela_wire_264;
    wire new_Jinkela_wire_2477;
    wire new_Jinkela_wire_1066;
    wire _0344_;
    wire new_Jinkela_wire_1885;
    wire new_Jinkela_wire_536;
    wire new_Jinkela_wire_2999;
    wire new_Jinkela_wire_861;
    wire new_Jinkela_wire_2570;
    wire new_Jinkela_wire_3330;
    wire new_Jinkela_wire_2642;
    wire new_Jinkela_wire_2768;
    wire new_Jinkela_wire_210;
    wire new_Jinkela_wire_182;
    wire _0732_;
    wire new_Jinkela_wire_3047;
    wire new_Jinkela_wire_1669;
    wire new_Jinkela_wire_3033;
    wire new_Jinkela_wire_322;
    wire new_Jinkela_wire_1916;
    wire new_Jinkela_wire_707;
    wire _0188_;
    wire _0638_;
    wire _0321_;
    wire new_Jinkela_wire_726;
    wire new_Jinkela_wire_1935;
    wire _0328_;
    wire new_Jinkela_wire_447;
    wire new_Jinkela_wire_765;
    wire new_Jinkela_wire_99;
    wire _0018_;
    wire new_Jinkela_wire_1768;
    wire new_Jinkela_wire_1664;
    wire new_Jinkela_wire_174;
    wire new_Jinkela_wire_2166;
    wire _0064_;
    wire new_Jinkela_wire_231;
    wire new_Jinkela_wire_2542;
    wire new_Jinkela_wire_1419;
    wire _0274_;
    wire new_Jinkela_wire_2179;
    wire new_Jinkela_wire_140;
    wire new_Jinkela_wire_1797;
    wire new_Jinkela_wire_316;
    wire new_Jinkela_wire_2029;
    wire new_Jinkela_wire_1987;
    wire _0586_;
    wire _0125_;
    wire new_Jinkela_wire_2033;
    wire new_Jinkela_wire_3247;
    wire new_Jinkela_wire_2095;
    wire new_Jinkela_wire_1596;
    wire new_Jinkela_wire_2284;
    wire _0364_;
    wire new_Jinkela_wire_2173;
    wire new_Jinkela_wire_729;
    wire new_Jinkela_wire_1710;
    wire new_Jinkela_wire_2879;
    wire new_Jinkela_wire_1551;
    wire new_Jinkela_wire_2837;
    wire _0214_;
    wire new_Jinkela_wire_352;
    wire new_Jinkela_wire_1792;
    wire new_Jinkela_wire_3149;
    wire new_Jinkela_wire_884;
    wire new_Jinkela_wire_2237;
    wire _0255_;
    wire new_Jinkela_wire_3273;
    wire new_Jinkela_wire_2667;
    wire new_Jinkela_wire_1197;
    wire _0714_;
    wire new_Jinkela_wire_970;
    wire new_Jinkela_wire_3012;
    wire new_Jinkela_wire_2614;
    wire new_Jinkela_wire_476;
    wire new_Jinkela_wire_2661;
    wire new_Jinkela_wire_1417;
    wire new_Jinkela_wire_1734;
    wire new_Jinkela_wire_1735;
    wire new_Jinkela_wire_728;
    wire new_Jinkela_wire_2567;
    wire new_Jinkela_wire_2522;
    wire new_Jinkela_wire_1991;
    wire new_Jinkela_wire_2167;
    wire _0400_;
    wire new_Jinkela_wire_1673;
    wire new_Jinkela_wire_44;
    wire _0508_;
    wire new_Jinkela_wire_758;
    wire _0173_;
    wire new_Jinkela_wire_401;
    wire new_Jinkela_wire_1270;
    wire new_Jinkela_wire_787;
    wire new_Jinkela_wire_2692;
    wire new_Jinkela_wire_3008;
    wire _0342_;
    wire new_Jinkela_wire_1721;
    wire new_Jinkela_wire_1614;
    wire new_Jinkela_wire_3275;
    wire new_Jinkela_wire_838;
    wire new_Jinkela_wire_2769;
    wire new_Jinkela_wire_1468;
    wire new_Jinkela_wire_1386;
    wire new_Jinkela_wire_1000;
    wire _0305_;
    wire new_Jinkela_wire_1992;
    wire new_Jinkela_wire_2533;
    wire new_Jinkela_wire_425;
    wire new_Jinkela_wire_652;
    wire new_Jinkela_wire_521;
    wire new_Jinkela_wire_3042;
    wire new_Jinkela_wire_2249;
    wire new_Jinkela_wire_2372;
    wire new_Jinkela_wire_2142;
    wire new_Jinkela_wire_1253;
    wire new_Jinkela_wire_1002;
    wire new_Jinkela_wire_293;
    wire new_Jinkela_wire_1399;
    wire new_Jinkela_wire_903;
    wire new_Jinkela_wire_1439;
    wire _0482_;
    wire new_Jinkela_wire_2589;
    wire _0659_;
    wire new_Jinkela_wire_2794;
    wire new_Jinkela_wire_1042;
    wire new_Jinkela_wire_2665;
    wire new_Jinkela_wire_2693;
    wire new_Jinkela_wire_3026;
    wire _0675_;
    wire new_Jinkela_wire_285;
    wire new_Jinkela_wire_934;
    wire new_Jinkela_wire_2320;
    wire new_Jinkela_wire_2172;
    wire new_Jinkela_wire_1362;
    wire new_Jinkela_wire_1952;
    wire new_Jinkela_wire_3160;
    wire new_Jinkela_wire_928;
    wire _0046_;
    wire new_Jinkela_wire_898;
    wire new_Jinkela_wire_3143;
    wire new_Jinkela_wire_633;
    wire new_Jinkela_wire_1291;
    wire new_Jinkela_wire_2861;
    wire new_Jinkela_wire_1493;
    wire new_Jinkela_wire_1453;
    wire new_Jinkela_wire_939;
    wire new_Jinkela_wire_2992;
    wire new_Jinkela_wire_66;
    wire new_Jinkela_wire_1443;
    wire _0151_;
    wire new_Jinkela_wire_1287;
    wire new_Jinkela_wire_1668;
    wire new_Jinkela_wire_241;
    wire new_Jinkela_wire_120;
    wire _0112_;
    wire new_Jinkela_wire_2245;
    wire _0615_;
    wire new_Jinkela_wire_2301;
    wire new_Jinkela_wire_1837;
    wire new_Jinkela_wire_403;
    wire _0521_;
    wire new_Jinkela_wire_19;
    wire new_Jinkela_wire_630;
    wire new_Jinkela_wire_53;
    wire new_Jinkela_wire_1146;
    wire new_Jinkela_wire_2936;
    wire new_Jinkela_wire_1815;
    wire new_Jinkela_wire_1084;
    wire new_Jinkela_wire_2728;
    wire new_Jinkela_wire_2243;
    wire new_Jinkela_wire_47;
    wire new_Jinkela_wire_2118;
    wire new_Jinkela_wire_2197;
    wire _0706_;
    wire _0725_;
    wire _0238_;
    wire new_Jinkela_wire_192;
    wire new_Jinkela_wire_2040;
    wire new_Jinkela_wire_3291;
    wire new_Jinkela_wire_2638;
    wire new_Jinkela_wire_2713;
    wire new_Jinkela_wire_2951;
    wire new_Jinkela_wire_2144;
    wire new_Jinkela_wire_2864;
    wire new_Jinkela_wire_2555;
    wire new_Jinkela_wire_1590;
    wire new_Jinkela_wire_377;
    wire _0147_;
    wire new_Jinkela_wire_119;
    wire new_Jinkela_wire_103;
    wire new_Jinkela_wire_2736;
    wire _0758_;
    wire new_Jinkela_wire_2356;
    wire new_Jinkela_wire_2014;
    wire new_Jinkela_wire_2354;
    wire _0700_;
    wire _0439_;
    wire new_Jinkela_wire_1891;
    wire new_Jinkela_wire_1787;
    wire new_Jinkela_wire_2240;
    wire _0411_;
    wire new_Jinkela_wire_2027;
    wire _0730_;
    wire new_Jinkela_wire_1626;
    wire _0207_;
    wire new_Jinkela_wire_1780;
    wire _0353_;
    wire new_Jinkela_wire_975;
    wire new_Jinkela_wire_2745;
    wire new_Jinkela_wire_938;
    wire _0245_;
    wire new_Jinkela_wire_1208;
    wire new_Jinkela_wire_896;
    wire new_Jinkela_wire_2676;
    wire new_Jinkela_wire_2666;
    wire new_Jinkela_wire_1589;
    wire new_Jinkela_wire_1172;
    wire new_Jinkela_wire_309;
    wire new_Jinkela_wire_1447;
    wire new_Jinkela_wire_926;
    wire new_Jinkela_wire_2826;
    wire new_Jinkela_wire_2962;
    wire new_Jinkela_wire_1041;
    wire new_Jinkela_wire_3146;
    wire new_Jinkela_wire_1184;
    wire new_Jinkela_wire_2432;
    wire new_Jinkela_wire_1961;
    wire new_Jinkela_wire_2792;
    wire new_Jinkela_wire_753;
    wire _0070_;
    wire new_Jinkela_wire_3294;
    wire new_Jinkela_wire_967;
    wire new_Jinkela_wire_2703;
    wire _0298_;
    wire new_Jinkela_wire_1155;
    wire new_Jinkela_wire_1381;
    wire new_Jinkela_wire_1435;
    wire _0138_;
    wire new_Jinkela_wire_1666;
    wire _0581_;
    wire _0680_;
    wire new_Jinkela_wire_2610;
    wire new_Jinkela_wire_1107;
    wire new_Jinkela_wire_2881;
    wire new_Jinkela_wire_488;
    wire _0059_;
    wire new_Jinkela_wire_2220;
    wire new_Jinkela_wire_696;
    wire new_Jinkela_wire_2516;
    wire new_Jinkela_wire_863;
    wire new_Jinkela_wire_2596;
    wire new_Jinkela_wire_782;
    wire _0480_;
    wire new_Jinkela_wire_588;
    wire new_Jinkela_wire_1506;
    wire _0540_;
    wire new_Jinkela_wire_1451;
    wire new_Jinkela_wire_2194;
    wire new_Jinkela_wire_1577;
    wire _0266_;
    wire new_Jinkela_wire_2929;
    wire _0444_;
    wire new_Jinkela_wire_332;
    wire new_Jinkela_wire_586;
    wire new_Jinkela_wire_2077;
    wire new_Jinkela_wire_879;
    wire new_Jinkela_wire_1739;
    wire new_Jinkela_wire_2063;
    wire new_Jinkela_wire_3312;
    wire _0598_;
    wire new_Jinkela_wire_923;
    wire new_Jinkela_wire_1478;
    wire new_Jinkela_wire_3239;
    wire _0309_;
    wire new_Jinkela_wire_1037;
    wire _0442_;
    wire new_Jinkela_wire_2615;
    wire new_Jinkela_wire_2799;
    wire _0647_;
    wire new_Jinkela_wire_2149;
    wire new_Jinkela_wire_1175;
    wire new_Jinkela_wire_214;
    wire new_Jinkela_wire_2804;
    wire new_Jinkela_wire_978;
    wire new_Jinkela_wire_1715;
    wire _0301_;
    wire new_Jinkela_wire_2989;
    wire new_Jinkela_wire_2502;
    wire new_Jinkela_wire_17;
    wire new_Jinkela_wire_538;
    wire new_Jinkela_wire_1450;
    wire _0111_;
    wire _0106_;
    wire new_Jinkela_wire_2705;
    wire new_Jinkela_wire_931;
    wire new_Jinkela_wire_1724;
    wire _0661_;
    wire new_Jinkela_wire_1281;
    wire new_Jinkela_wire_764;
    wire new_Jinkela_wire_1101;
    wire new_Jinkela_wire_272;
    wire new_Jinkela_wire_1712;
    wire _0055_;
    wire new_Jinkela_wire_2291;
    wire new_Jinkela_wire_1360;
    wire new_Jinkela_wire_323;
    wire new_Jinkela_wire_855;
    wire new_Jinkela_wire_215;
    wire _0363_;
    wire new_Jinkela_wire_1862;
    wire new_Jinkela_wire_1701;
    wire new_Jinkela_wire_1615;
    wire new_Jinkela_wire_636;
    wire new_Jinkela_wire_456;
    wire new_Jinkela_wire_2785;
    wire new_Jinkela_wire_2969;
    wire new_Jinkela_wire_115;
    wire new_Jinkela_wire_1059;
    wire new_Jinkela_wire_1584;
    wire _0717_;
    wire new_Jinkela_wire_1460;
    wire new_Jinkela_wire_949;
    wire new_Jinkela_wire_2593;
    wire new_Jinkela_wire_902;
    wire new_Jinkela_wire_727;
    wire new_Jinkela_wire_1286;
    wire _0001_;
    wire _0350_;
    wire new_Jinkela_wire_3078;
    wire new_Jinkela_wire_281;
    wire _0300_;
    wire new_Jinkela_wire_440;
    wire new_Jinkela_wire_1432;
    wire _0718_;
    wire new_Jinkela_wire_3326;
    wire new_Jinkela_wire_284;
    wire new_Jinkela_wire_972;
    wire new_Jinkela_wire_2454;
    wire new_Jinkela_wire_1160;
    wire new_Jinkela_wire_593;
    wire new_Jinkela_wire_104;
    wire _0017_;
    wire new_Jinkela_wire_2551;
    wire new_Jinkela_wire_1772;
    wire new_Jinkela_wire_1398;
    wire new_Jinkela_wire_2341;
    wire _0679_;
    wire new_Jinkela_wire_1694;
    wire _0037_;
    wire new_Jinkela_wire_365;
    wire new_Jinkela_wire_510;
    wire new_Jinkela_wire_1789;
    wire new_Jinkela_wire_129;
    wire new_Jinkela_wire_2122;
    wire new_Jinkela_wire_1711;
    wire new_Jinkela_wire_658;
    wire new_Jinkela_wire_2433;
    wire _0136_;
    wire new_Jinkela_wire_1019;
    wire _0194_;
    wire new_Jinkela_wire_1082;
    wire new_Jinkela_wire_832;
    wire _0099_;
    wire _0466_;
    wire new_Jinkela_wire_1370;
    wire _0236_;
    wire new_Jinkela_wire_1602;
    wire new_Jinkela_wire_2660;
    wire _0537_;
    wire new_Jinkela_wire_92;
    wire new_Jinkela_wire_2489;
    wire _0496_;
    wire new_Jinkela_wire_179;
    wire new_Jinkela_wire_574;
    wire new_Jinkela_wire_2370;
    wire new_Jinkela_wire_613;
    wire new_Jinkela_wire_2254;
    wire new_Jinkela_wire_1884;
    wire new_Jinkela_wire_1025;
    wire new_Jinkela_wire_1576;
    wire new_Jinkela_wire_3066;
    wire _0159_;
    wire _0391_;
    wire new_Jinkela_wire_2386;
    wire new_Jinkela_wire_2565;
    wire new_Jinkela_wire_1996;
    wire _0183_;
    wire _0416_;
    wire _0021_;
    wire new_Jinkela_wire_3193;
    wire new_Jinkela_wire_2482;
    wire new_Jinkela_wire_2889;
    wire new_Jinkela_wire_3067;
    wire new_Jinkela_wire_2624;
    wire new_Jinkela_wire_1684;
    wire new_Jinkela_wire_1483;
    wire new_Jinkela_wire_1910;
    wire new_Jinkela_wire_81;
    wire new_Jinkela_wire_381;
    wire new_Jinkela_wire_2225;
    wire _0131_;
    wire new_Jinkela_wire_2899;
    wire new_Jinkela_wire_1680;
    wire new_Jinkela_wire_2901;
    wire new_Jinkela_wire_2612;
    wire new_Jinkela_wire_2362;
    wire new_Jinkela_wire_1774;
    wire new_Jinkela_wire_2247;
    wire new_Jinkela_wire_3039;
    wire new_Jinkela_wire_1157;
    wire _0062_;
    wire new_Jinkela_wire_1499;
    wire new_Jinkela_wire_1706;
    wire new_Jinkela_wire_2970;
    wire new_Jinkela_wire_1401;
    wire new_Jinkela_wire_2467;
    wire new_Jinkela_wire_1001;
    wire new_Jinkela_wire_2348;
    wire new_Jinkela_wire_1844;
    wire new_Jinkela_wire_23;
    wire _0003_;
    wire _0119_;
    wire new_Jinkela_wire_559;
    wire new_Jinkela_wire_251;
    wire new_Jinkela_wire_2475;
    wire _0607_;
    wire new_Jinkela_wire_2787;
    wire new_Jinkela_wire_2347;
    wire new_Jinkela_wire_2091;
    wire new_Jinkela_wire_2020;
    wire new_Jinkela_wire_1702;
    wire new_Jinkela_wire_1492;
    wire _0619_;
    wire _0398_;
    wire new_Jinkela_wire_1210;
    wire new_Jinkela_wire_650;
    wire new_Jinkela_wire_226;
    wire new_Jinkela_wire_2212;
    wire new_Jinkela_wire_676;
    wire new_Jinkela_wire_1820;
    wire new_Jinkela_wire_1109;
    wire new_Jinkela_wire_3232;
    wire new_Jinkela_wire_1375;
    wire new_Jinkela_wire_480;
    wire _0096_;
    wire _0296_;
    wire new_Jinkela_wire_348;
    wire _0529_;
    wire new_Jinkela_wire_2350;
    wire new_Jinkela_wire_589;
    wire _0608_;
    wire _0694_;
    wire new_Jinkela_wire_708;
    wire new_Jinkela_wire_315;
    wire new_Jinkela_wire_2458;
    wire new_Jinkela_wire_2064;
    wire _0612_;
    wire new_Jinkela_wire_1480;
    wire new_Jinkela_wire_1773;
    wire new_Jinkela_wire_996;
    wire new_Jinkela_wire_2823;
    wire _0635_;
    wire new_Jinkela_wire_240;
    wire new_Jinkela_wire_417;
    wire _0225_;
    wire new_Jinkela_wire_910;
    wire new_Jinkela_wire_577;
    wire new_Jinkela_wire_603;
    wire new_Jinkela_wire_3302;
    wire _0705_;
    wire new_Jinkela_wire_255;
    wire _0195_;
    wire _0709_;
    wire new_Jinkela_wire_1092;
    wire new_Jinkela_wire_3195;
    wire _0757_;
    wire new_Jinkela_wire_1367;
    wire new_Jinkela_wire_1637;
    wire _0084_;
    wire new_Jinkela_wire_2139;
    wire new_Jinkela_wire_125;
    wire new_Jinkela_wire_2479;
    wire new_Jinkela_wire_683;
    wire new_Jinkela_wire_3003;
    wire new_Jinkela_wire_959;
    wire new_Jinkela_wire_1379;
    wire new_Jinkela_wire_518;
    wire new_Jinkela_wire_2795;
    wire new_Jinkela_wire_2332;
    wire new_Jinkela_wire_474;
    wire new_Jinkela_wire_803;
    wire _0283_;
    wire new_Jinkela_wire_3167;
    wire new_Jinkela_wire_1730;
    wire new_Jinkela_wire_3220;
    wire new_Jinkela_wire_1330;
    wire new_Jinkela_wire_6;
    wire new_Jinkela_wire_2441;
    wire new_Jinkela_wire_178;
    wire _0156_;
    wire new_Jinkela_wire_1455;
    wire new_Jinkela_wire_355;
    wire new_Jinkela_wire_977;
    wire new_Jinkela_wire_2285;
    wire new_Jinkela_wire_2130;
    wire new_Jinkela_wire_1428;
    wire new_Jinkela_wire_2297;
    wire new_Jinkela_wire_1023;
    wire new_Jinkela_wire_3034;
    wire new_Jinkela_wire_2812;
    wire new_Jinkela_wire_200;
    wire new_Jinkela_wire_1800;
    wire new_Jinkela_wire_3156;
    wire new_Jinkela_wire_1031;
    wire new_Jinkela_wire_1228;
    wire new_Jinkela_wire_2739;
    wire _0762_;
    wire new_Jinkela_wire_1914;
    wire new_Jinkela_wire_235;
    wire _0547_;
    wire new_Jinkela_wire_1842;
    wire new_Jinkela_wire_643;
    wire new_Jinkela_wire_1794;
    wire new_Jinkela_wire_286;
    wire new_Jinkela_wire_2330;
    wire new_Jinkela_wire_2955;
    wire new_Jinkela_wire_520;
    wire _0534_;
    wire new_Jinkela_wire_2321;
    wire new_Jinkela_wire_3258;
    wire new_Jinkela_wire_2088;
    wire new_Jinkela_wire_84;
    wire _0166_;
    wire new_Jinkela_wire_1817;
    wire _0079_;
    wire new_Jinkela_wire_2119;
    wire new_Jinkela_wire_1638;
    wire new_Jinkela_wire_2960;
    wire new_Jinkela_wire_547;
    wire new_Jinkela_wire_1595;
    wire new_Jinkela_wire_933;
    wire new_Jinkela_wire_1718;
    wire new_Jinkela_wire_489;
    wire new_Jinkela_wire_3153;
    wire new_Jinkela_wire_1448;
    wire new_Jinkela_wire_2659;
    wire new_Jinkela_wire_363;
    wire new_Jinkela_wire_2193;
    wire new_Jinkela_wire_2067;
    wire _0240_;
    wire _0378_;
    wire new_Jinkela_wire_1234;
    wire _0409_;
    wire new_Jinkela_wire_1355;
    wire _0441_;
    wire _0126_;
    wire _0020_;
    wire _0448_;
    wire new_Jinkela_wire_3134;
    wire new_Jinkela_wire_2050;
    wire _0784_;
    wire new_Jinkela_wire_868;
    wire new_Jinkela_wire_830;
    wire new_Jinkela_wire_1276;
    wire new_Jinkela_wire_1074;
    wire new_Jinkela_wire_1159;
    wire _0215_;
    wire _0209_;
    wire new_Jinkela_wire_2974;
    wire _0668_;
    wire _0663_;
    wire new_Jinkela_wire_3030;
    wire new_Jinkela_wire_3071;
    wire new_Jinkela_wire_908;
    wire new_Jinkela_wire_310;
    wire _0199_;
    wire _0281_;
    wire new_Jinkela_wire_1223;
    wire _0704_;
    wire new_Jinkela_wire_1578;
    wire new_Jinkela_wire_1058;
    wire new_Jinkela_wire_3151;
    wire new_Jinkela_wire_2116;
    wire new_Jinkela_wire_2669;
    wire new_Jinkela_wire_2373;
    wire new_Jinkela_wire_2763;
    wire new_Jinkela_wire_243;
    wire new_Jinkela_wire_1252;
    wire new_Jinkela_wire_1829;
    wire _0057_;
    wire _0031_;
    wire new_Jinkela_wire_1652;
    wire new_Jinkela_wire_2109;
    wire new_Jinkela_wire_1777;
    wire new_Jinkela_wire_3305;
    wire new_Jinkela_wire_385;
    wire _0782_;
    wire new_Jinkela_wire_1003;
    wire new_Jinkela_wire_2273;
    wire new_Jinkela_wire_1464;
    wire new_Jinkela_wire_3308;
    wire new_Jinkela_wire_2038;
    wire new_Jinkela_wire_2564;
    wire _0069_;
    wire _0655_;
    wire new_Jinkela_wire_2602;
    wire new_Jinkela_wire_416;
    wire _0108_;
    wire new_Jinkela_wire_2013;
    wire new_Jinkela_wire_1317;
    wire new_Jinkela_wire_2818;
    wire new_Jinkela_wire_2862;
    wire new_Jinkela_wire_2582;
    wire new_Jinkela_wire_2606;
    wire _0100_;
    wire new_Jinkela_wire_61;
    wire new_Jinkela_wire_463;
    wire new_Jinkela_wire_815;
    wire new_Jinkela_wire_1087;
    wire new_Jinkela_wire_3063;
    wire new_Jinkela_wire_317;
    wire _0776_;
    wire new_Jinkela_wire_1624;
    wire new_Jinkela_wire_3272;
    wire new_Jinkela_wire_712;
    wire _0672_;
    wire new_Jinkela_wire_3031;
    wire _0186_;
    wire new_Jinkela_wire_2700;
    wire new_Jinkela_wire_1238;
    wire new_Jinkela_wire_1038;
    wire new_Jinkela_wire_2670;
    wire new_Jinkela_wire_2066;
    wire new_Jinkela_wire_1274;
    wire new_Jinkela_wire_871;
    wire _0451_;
    wire _0462_;
    wire _0538_;
    wire new_Jinkela_wire_1850;
    wire new_Jinkela_wire_2983;
    wire new_Jinkela_wire_3006;
    wire _0330_;
    wire new_Jinkela_wire_3109;
    wire new_Jinkela_wire_2539;
    wire _0073_;
    wire new_Jinkela_wire_2244;
    wire new_Jinkela_wire_172;
    wire new_Jinkela_wire_95;
    wire new_Jinkela_wire_2647;
    wire new_Jinkela_wire_170;
    wire new_Jinkela_wire_1926;
    wire new_Jinkela_wire_1898;
    wire new_Jinkela_wire_1039;
    wire _0023_;
    wire new_Jinkela_wire_2423;
    wire new_Jinkela_wire_2155;
    wire new_Jinkela_wire_2603;
    wire new_Jinkela_wire_2530;
    wire new_Jinkela_wire_2808;
    wire new_Jinkela_wire_2885;
    wire new_Jinkela_wire_32;
    wire new_Jinkela_wire_1892;
    wire new_Jinkela_wire_2529;
    wire new_Jinkela_wire_1827;
    wire new_Jinkela_wire_1340;
    wire new_Jinkela_wire_48;
    wire new_Jinkela_wire_397;
    wire new_Jinkela_wire_2500;
    wire new_Jinkela_wire_212;
    wire _0294_;
    wire new_Jinkela_wire_964;
    wire new_Jinkela_wire_848;
    wire new_Jinkela_wire_3027;
    wire new_Jinkela_wire_410;
    wire new_Jinkela_wire_1458;
    wire new_Jinkela_wire_1202;
    wire _0187_;
    wire new_Jinkela_wire_2451;
    wire new_Jinkela_wire_2287;
    wire new_Jinkela_wire_3083;
    wire new_Jinkela_wire_302;
    wire new_Jinkela_wire_1134;
    wire new_Jinkela_wire_404;
    wire new_Jinkela_wire_1646;
    wire new_Jinkela_wire_3148;
    wire new_Jinkela_wire_922;
    wire new_Jinkela_wire_2584;
    wire new_Jinkela_wire_943;
    wire new_Jinkela_wire_549;
    wire new_Jinkela_wire_1811;
    wire new_Jinkela_wire_514;
    wire new_Jinkela_wire_270;
    wire new_Jinkela_wire_1053;
    wire new_Jinkela_wire_2623;
    wire _0407_;
    wire new_Jinkela_wire_2752;
    wire _0731_;
    wire new_Jinkela_wire_1090;
    wire new_Jinkela_wire_822;
    wire new_Jinkela_wire_1765;
    wire _0662_;
    wire new_Jinkela_wire_2251;
    wire new_Jinkela_wire_1060;
    wire new_Jinkela_wire_1429;
    wire new_Jinkela_wire_0;
    wire new_Jinkela_wire_1985;
    wire new_Jinkela_wire_1540;
    wire new_Jinkela_wire_568;
    wire _0030_;
    wire new_Jinkela_wire_1631;
    wire new_Jinkela_wire_2607;
    wire new_Jinkela_wire_1525;
    wire new_Jinkela_wire_1861;
    wire new_Jinkela_wire_503;
    wire _0317_;
    wire new_Jinkela_wire_645;
    wire new_Jinkela_wire_2894;
    wire new_Jinkela_wire_2888;
    wire new_Jinkela_wire_94;
    wire new_Jinkela_wire_2464;
    wire new_Jinkela_wire_1079;
    wire new_Jinkela_wire_875;
    wire new_Jinkela_wire_944;
    wire new_Jinkela_wire_438;
    wire new_Jinkela_wire_1723;
    wire new_Jinkela_wire_1969;
    wire new_Jinkela_wire_860;
    wire _0503_;
    wire _0268_;
    wire new_Jinkela_wire_3321;
    wire new_Jinkela_wire_1719;
    wire new_Jinkela_wire_3001;
    wire new_Jinkela_wire_791;
    wire new_Jinkela_wire_2559;
    wire new_Jinkela_wire_862;
    wire new_Jinkela_wire_1758;
    wire new_Jinkela_wire_3079;
    wire new_Jinkela_wire_2453;
    wire new_Jinkela_wire_2773;
    wire new_Jinkela_wire_1050;
    wire new_Jinkela_wire_2089;
    wire new_Jinkela_wire_2566;
    wire new_Jinkela_wire_2210;
    wire _0574_;
    wire new_Jinkela_wire_2844;
    wire new_Jinkela_wire_2753;
    wire new_Jinkela_wire_2416;
    wire new_Jinkela_wire_386;
    wire new_Jinkela_wire_3289;
    wire new_Jinkela_wire_2517;
    wire new_Jinkela_wire_2825;
    wire new_Jinkela_wire_2513;
    wire new_Jinkela_wire_1121;
    wire new_Jinkela_wire_1111;
    wire _0347_;
    wire new_Jinkela_wire_357;
    wire new_Jinkela_wire_366;
    wire new_Jinkela_wire_601;
    wire new_Jinkela_wire_2803;
    wire _0174_;
    wire new_Jinkela_wire_216;
    wire new_Jinkela_wire_1982;
    wire new_Jinkela_wire_2258;
    wire new_Jinkela_wire_3126;
    wire new_Jinkela_wire_1147;
    wire new_Jinkela_wire_2628;
    wire new_Jinkela_wire_1430;
    wire new_Jinkela_wire_1481;
    wire new_Jinkela_wire_118;
    wire new_Jinkela_wire_1633;
    wire new_Jinkela_wire_2326;
    wire _0362_;
    wire new_Jinkela_wire_3229;
    wire new_Jinkela_wire_1726;
    wire _0569_;
    wire new_Jinkela_wire_2772;
    wire new_Jinkela_wire_3267;
    wire new_Jinkela_wire_819;
    wire new_Jinkela_wire_1237;
    wire new_Jinkela_wire_1998;
    wire new_Jinkela_wire_2510;
    wire new_Jinkela_wire_2552;
    wire _0316_;
    wire new_Jinkela_wire_2001;
    wire new_Jinkela_wire_2024;
    wire new_Jinkela_wire_409;
    wire new_Jinkela_wire_2256;
    wire new_Jinkela_wire_2732;
    wire new_Jinkela_wire_320;
    wire new_Jinkela_wire_3228;
    wire new_Jinkela_wire_1106;
    wire new_Jinkela_wire_1378;
    wire new_Jinkela_wire_2782;
    wire new_Jinkela_wire_2867;
    wire new_Jinkela_wire_2910;
    wire new_Jinkela_wire_1230;
    wire new_Jinkela_wire_1327;
    wire new_Jinkela_wire_3246;
    wire new_Jinkela_wire_882;
    wire new_Jinkela_wire_2043;
    wire new_Jinkela_wire_2023;
    wire new_Jinkela_wire_1727;
    wire _0220_;
    wire new_Jinkela_wire_2828;
    wire new_Jinkela_wire_2296;
    wire new_Jinkela_wire_3265;
    wire _0403_;
    wire new_Jinkela_wire_2731;
    wire new_Jinkela_wire_1641;
    wire new_Jinkela_wire_72;
    wire new_Jinkela_wire_1078;
    wire new_Jinkela_wire_3112;
    wire _0241_;
    wire new_Jinkela_wire_1938;
    wire new_Jinkela_wire_2367;
    wire new_Jinkela_wire_1503;
    wire new_Jinkela_wire_2270;
    wire new_Jinkela_wire_2865;
    wire new_Jinkela_wire_1068;
    wire new_Jinkela_wire_3070;
    wire new_Jinkela_wire_2140;
    wire _0518_;
    wire new_Jinkela_wire_2465;
    wire new_Jinkela_wire_246;
    wire new_Jinkela_wire_1342;
    wire new_Jinkela_wire_188;
    wire new_Jinkela_wire_3002;
    wire new_Jinkela_wire_304;
    wire _0114_;
    wire new_Jinkela_wire_2571;
    wire new_Jinkela_wire_1627;
    wire _0443_;
    wire _0437_;
    wire new_Jinkela_wire_2973;
    wire _0585_;
    wire _0773_;
    wire new_Jinkela_wire_2846;
    wire new_Jinkela_wire_1836;
    wire new_Jinkela_wire_396;
    wire new_Jinkela_wire_2057;
    wire new_Jinkela_wire_581;
    wire new_Jinkela_wire_1569;
    wire new_Jinkela_wire_2310;
    wire new_Jinkela_wire_2685;
    wire new_Jinkela_wire_1163;
    wire new_Jinkela_wire_2543;
    wire new_net_1483;
    wire new_Jinkela_wire_1568;
    wire new_Jinkela_wire_486;
    wire new_Jinkela_wire_68;
    wire new_Jinkela_wire_2776;
    wire new_Jinkela_wire_519;
    wire new_Jinkela_wire_3144;
    wire new_Jinkela_wire_2076;
    wire new_Jinkela_wire_407;
    wire new_Jinkela_wire_2151;
    wire _0077_;
    wire new_Jinkela_wire_606;
    wire new_Jinkela_wire_2203;
    wire new_Jinkela_wire_3319;
    wire _0743_;
    wire new_Jinkela_wire_462;
    wire _0273_;
    wire new_Jinkela_wire_1741;
    wire new_Jinkela_wire_1732;
    wire new_Jinkela_wire_576;
    wire new_Jinkela_wire_743;
    wire new_Jinkela_wire_1670;
    wire new_Jinkela_wire_1583;
    wire new_Jinkela_wire_2587;
    wire _0587_;
    wire new_Jinkela_wire_336;
    wire new_Jinkela_wire_2616;
    wire new_Jinkela_wire_833;
    wire new_Jinkela_wire_354;
    wire new_Jinkela_wire_1144;
    wire new_Jinkela_wire_1977;
    wire new_Jinkela_wire_1832;
    wire _0191_;
    wire _0155_;
    wire new_Jinkela_wire_2654;
    wire _0609_;
    wire new_Jinkela_wire_783;
    wire new_Jinkela_wire_373;
    wire new_Jinkela_wire_3217;
    wire new_Jinkela_wire_1839;
    wire new_Jinkela_wire_1746;
    wire new_Jinkela_wire_2729;
    wire new_Jinkela_wire_681;
    wire _0625_;
    wire _0460_;
    wire new_Jinkela_wire_469;
    wire new_Jinkela_wire_988;
    wire new_Jinkela_wire_1620;
    wire new_Jinkela_wire_1491;
    wire new_Jinkela_wire_2521;
    wire _0247_;
    wire new_Jinkela_wire_457;
    wire new_Jinkela_wire_2664;
    wire new_Jinkela_wire_3097;
    wire new_Jinkela_wire_920;
    wire new_Jinkela_wire_3306;
    wire new_Jinkela_wire_3192;
    wire new_Jinkela_wire_2159;
    wire _0710_;
    wire new_Jinkela_wire_872;
    wire _0664_;
    wire new_Jinkela_wire_1939;
    wire _0541_;
    wire new_Jinkela_wire_2295;
    wire new_Jinkela_wire_1225;
    wire new_Jinkela_wire_1798;
    wire new_Jinkela_wire_2015;
    wire new_Jinkela_wire_2322;
    wire new_net_6;
    wire _0495_;
    wire new_Jinkela_wire_930;
    wire new_Jinkela_wire_2271;
    wire new_Jinkela_wire_702;
    wire new_Jinkela_wire_3094;
    wire new_Jinkela_wire_2388;
    wire new_Jinkela_wire_3298;
    wire _0721_;
    wire new_Jinkela_wire_3136;
    wire new_Jinkela_wire_2230;
    wire _0406_;
    wire new_Jinkela_wire_1153;
    wire new_Jinkela_wire_2783;
    wire new_Jinkela_wire_724;
    wire new_Jinkela_wire_1470;
    wire new_Jinkela_wire_2987;
    wire new_Jinkela_wire_816;
    wire new_Jinkela_wire_720;
    wire _0048_;
    wire new_Jinkela_wire_3262;
    wire new_Jinkela_wire_604;
    wire _0510_;
    wire new_Jinkela_wire_2575;
    wire new_Jinkela_wire_2224;
    wire new_Jinkela_wire_319;
    wire new_Jinkela_wire_41;
    wire new_Jinkela_wire_1056;
    wire new_Jinkela_wire_1886;
    wire _0475_;
    wire new_Jinkela_wire_2932;
    wire new_Jinkela_wire_1165;
    wire new_Jinkela_wire_1955;
    wire _0506_;
    wire new_Jinkela_wire_218;
    wire _0622_;
    wire _0578_;
    wire new_Jinkela_wire_1307;
    wire new_Jinkela_wire_2111;
    wire new_Jinkela_wire_2576;
    wire new_Jinkela_wire_809;
    wire new_Jinkela_wire_130;
    wire new_Jinkela_wire_481;
    wire new_Jinkela_wire_3154;
    wire new_Jinkela_wire_483;
    wire new_Jinkela_wire_1511;
    wire new_Jinkela_wire_2747;
    wire new_Jinkela_wire_1662;
    wire new_Jinkela_wire_2677;
    wire new_Jinkela_wire_3202;
    wire _0572_;
    wire new_Jinkela_wire_2868;
    wire new_Jinkela_wire_2751;
    wire new_Jinkela_wire_437;
    wire new_Jinkela_wire_2887;
    wire new_Jinkela_wire_350;
    wire new_Jinkela_wire_2171;
    wire new_Jinkela_wire_2688;
    wire new_Jinkela_wire_1752;
    wire new_Jinkela_wire_2990;
    wire new_Jinkela_wire_2836;
    wire new_Jinkela_wire_1989;
    wire new_Jinkela_wire_3287;
    wire new_Jinkela_wire_1128;
    wire _0110_;
    wire _0756_;
    wire new_Jinkela_wire_158;
    wire new_Jinkela_wire_2435;
    wire new_Jinkela_wire_3323;
    wire _0390_;
    wire new_Jinkela_wire_372;
    wire _0323_;
    wire new_Jinkela_wire_427;
    wire _0708_;
    wire new_Jinkela_wire_741;
    wire new_Jinkela_wire_232;
    wire new_Jinkela_wire_1069;
    wire new_Jinkela_wire_844;
    wire new_Jinkela_wire_1630;
    wire _0657_;
    wire new_Jinkela_wire_1877;
    wire new_Jinkela_wire_1348;
    wire new_Jinkela_wire_3122;
    wire _0684_;
    wire new_Jinkela_wire_718;
    wire new_Jinkela_wire_749;
    wire new_Jinkela_wire_2073;
    wire new_Jinkela_wire_1353;
    wire new_Jinkela_wire_1509;
    wire new_Jinkela_wire_3108;
    wire new_Jinkela_wire_2314;
    wire new_Jinkela_wire_1825;
    wire new_Jinkela_wire_2345;
    wire new_Jinkela_wire_3004;
    wire _0224_;
    wire new_Jinkela_wire_699;
    wire new_Jinkela_wire_1512;
    wire new_Jinkela_wire_571;
    wire _0531_;
    wire _0747_;
    wire _0753_;
    wire _0653_;
    wire new_Jinkela_wire_974;
    wire new_Jinkela_wire_126;
    wire new_Jinkela_wire_1923;
    wire new_Jinkela_wire_1659;
    wire new_Jinkela_wire_2933;
    wire new_Jinkela_wire_268;
    wire _0701_;
    wire new_Jinkela_wire_1136;
    wire _0075_;
    wire new_Jinkela_wire_2120;
    wire new_Jinkela_wire_3020;
    wire new_Jinkela_wire_810;
    wire new_Jinkela_wire_824;
    wire new_Jinkela_wire_527;
    wire new_Jinkela_wire_2232;
    wire new_Jinkela_wire_1951;
    wire new_Jinkela_wire_2133;
    wire new_Jinkela_wire_2758;
    wire new_Jinkela_wire_3084;
    wire new_Jinkela_wire_2710;
    wire new_Jinkela_wire_1094;
    wire new_Jinkela_wire_1528;
    wire new_Jinkela_wire_3157;
    wire new_Jinkela_wire_368;
    wire new_Jinkela_wire_2537;
    wire new_Jinkela_wire_1813;
    wire new_Jinkela_wire_719;
    wire _0197_;
    wire new_Jinkela_wire_1818;
    wire new_Jinkela_wire_306;
    wire new_Jinkela_wire_660;
    wire new_Jinkela_wire_3147;
    wire new_Jinkela_wire_2294;
    wire new_Jinkela_wire_3128;
    wire _0346_;
    wire new_Jinkela_wire_2842;
    wire new_Jinkela_wire_2313;
    wire new_Jinkela_wire_846;
    wire new_Jinkela_wire_1024;
    wire new_Jinkela_wire_3040;
    wire new_Jinkela_wire_3318;
    wire new_Jinkela_wire_3162;
    wire new_Jinkela_wire_1958;
    wire new_Jinkela_wire_786;
    wire new_Jinkela_wire_2132;
    wire _0632_;
    wire new_Jinkela_wire_1390;
    wire new_Jinkela_wire_108;
    wire new_Jinkela_wire_1098;
    wire _0422_;
    wire new_Jinkela_wire_2377;
    wire new_Jinkela_wire_1280;
    wire new_Jinkela_wire_888;
    wire new_Jinkela_wire_2594;
    wire new_Jinkela_wire_956;
    wire new_Jinkela_wire_482;
    wire new_Jinkela_wire_1182;
    wire new_Jinkela_wire_2487;
    wire new_Jinkela_wire_3222;
    wire new_Jinkela_wire_2945;
    wire _0011_;
    wire new_Jinkela_wire_735;
    wire _0744_;
    wire new_Jinkela_wire_91;
    wire new_Jinkela_wire_2746;
    wire new_Jinkela_wire_1461;
    wire new_Jinkela_wire_2874;
    wire new_Jinkela_wire_2940;
    wire new_Jinkela_wire_2044;
    wire _0787_;
    wire new_Jinkela_wire_2447;
    wire new_Jinkela_wire_2621;
    wire new_Jinkela_wire_811;
    wire _0554_;
    wire new_Jinkela_wire_2017;
    wire _0727_;
    wire new_Jinkela_wire_96;
    wire _0686_;
    wire new_Jinkela_wire_2026;
    wire new_Jinkela_wire_1749;
    wire new_Jinkela_wire_2514;
    wire new_Jinkela_wire_3132;
    wire new_Jinkela_wire_3055;
    wire new_Jinkela_wire_866;
    wire new_Jinkela_wire_1466;
    wire _0556_;
    wire _0337_;
    wire new_Jinkela_wire_725;
    wire _0693_;
    wire new_Jinkela_wire_493;
    wire new_Jinkela_wire_1648;
    wire new_Jinkela_wire_2592;
    wire new_Jinkela_wire_2086;
    wire _0171_;
    wire new_Jinkela_wire_54;
    wire new_Jinkela_wire_867;
    wire new_Jinkela_wire_672;
    wire new_Jinkela_wire_1888;
    wire new_Jinkela_wire_2009;
    wire new_Jinkela_wire_2740;
    wire new_Jinkela_wire_2205;
    wire new_Jinkela_wire_460;
    wire new_Jinkela_wire_3310;
    wire _0239_;
    wire new_Jinkela_wire_1879;
    wire new_Jinkela_wire_2281;
    wire _0006_;
    wire new_Jinkela_wire_2995;
    wire new_Jinkela_wire_647;
    wire new_Jinkela_wire_818;
    wire _0370_;
    wire new_Jinkela_wire_1204;
    wire new_Jinkela_wire_2261;
    wire new_Jinkela_wire_3197;
    wire _0417_;
    wire new_net_1463;
    wire new_Jinkela_wire_2892;
    wire new_Jinkela_wire_2771;
    wire new_Jinkela_wire_1764;
    wire new_Jinkela_wire_1139;
    wire new_Jinkela_wire_1559;
    wire new_Jinkela_wire_3145;
    wire new_Jinkela_wire_2257;
    wire new_Jinkela_wire_2704;
    wire new_Jinkela_wire_431;
    wire new_Jinkela_wire_2318;
    wire new_Jinkela_wire_168;
    wire _0211_;
    wire _0551_;
    wire _0033_;
    wire _0606_;
    wire new_Jinkela_wire_3235;
    wire new_Jinkela_wire_1613;
    wire new_Jinkela_wire_1441;
    wire new_Jinkela_wire_1477;
    wire new_Jinkela_wire_2793;
    wire new_Jinkela_wire_2327;
    wire _0276_;
    wire new_Jinkela_wire_2668;
    wire new_Jinkela_wire_360;
    wire new_Jinkela_wire_1168;
    wire new_Jinkela_wire_693;
    wire new_Jinkela_wire_2941;
    wire new_Jinkela_wire_2674;
    wire _0140_;
    wire new_Jinkela_wire_2262;
    wire new_Jinkela_wire_2527;
    wire new_Jinkela_wire_20;
    wire new_Jinkela_wire_1299;
    wire new_Jinkela_wire_1821;
    wire new_Jinkela_wire_653;
    wire new_Jinkela_wire_194;
    wire new_Jinkela_wire_3036;
    wire new_Jinkela_wire_177;
    wire new_Jinkela_wire_2165;
    wire new_Jinkela_wire_3266;
    wire new_Jinkela_wire_1527;
    wire new_Jinkela_wire_121;
    wire _0568_;
    wire new_Jinkela_wire_2279;
    wire new_Jinkela_wire_504;
    wire new_Jinkela_wire_2346;
    wire _0122_;
    wire new_Jinkela_wire_496;
    wire new_Jinkela_wire_67;
    wire new_Jinkela_wire_253;
    wire new_Jinkela_wire_428;
    wire new_Jinkela_wire_213;
    wire new_Jinkela_wire_767;
    wire _0473_;
    wire new_Jinkela_wire_1192;
    wire new_Jinkela_wire_459;
    wire new_Jinkela_wire_3090;
    wire new_Jinkela_wire_2756;
    wire new_Jinkela_wire_3100;
    wire new_Jinkela_wire_1859;
    wire new_Jinkela_wire_3327;
    wire new_Jinkela_wire_1166;
    wire _0399_;
    wire new_Jinkela_wire_537;
    wire new_Jinkela_wire_2645;
    wire new_Jinkela_wire_2641;
    wire new_Jinkela_wire_1212;
    wire new_Jinkela_wire_622;
    wire new_Jinkela_wire_2389;
    wire new_Jinkela_wire_3104;
    wire new_Jinkela_wire_2695;
    wire new_Jinkela_wire_523;
    wire new_Jinkela_wire_1530;
    wire new_Jinkela_wire_2000;
    wire new_Jinkela_wire_2557;
    wire new_Jinkela_wire_895;
    wire _0277_;
    wire new_Jinkela_wire_1099;
    wire new_Jinkela_wire_1927;
    wire new_Jinkela_wire_433;
    wire new_Jinkela_wire_2579;
    wire new_Jinkela_wire_453;
    wire new_Jinkela_wire_314;
    wire new_Jinkela_wire_1125;
    wire _0656_;
    wire new_Jinkela_wire_1554;
    wire new_Jinkela_wire_1135;
    wire _0648_;
    wire _0711_;
    wire new_Jinkela_wire_3168;
    wire new_Jinkela_wire_641;
    wire _0118_;
    wire new_Jinkela_wire_1835;
    wire new_Jinkela_wire_3115;
    wire new_Jinkela_wire_573;
    wire new_Jinkela_wire_2719;
    wire _0689_;
    wire new_Jinkela_wire_1872;
    wire _0012_;
    wire new_Jinkela_wire_845;
    wire _0621_;
    wire new_Jinkela_wire_1242;
    wire new_Jinkela_wire_2985;
    wire new_Jinkela_wire_220;
    wire new_Jinkela_wire_141;
    wire new_Jinkela_wire_3174;
    wire new_Jinkela_wire_62;
    wire new_Jinkela_wire_1006;
    wire new_Jinkela_wire_2848;
    wire _0061_;
    wire new_Jinkela_wire_2563;
    wire new_Jinkela_wire_1339;
    wire new_Jinkela_wire_1309;
    wire new_Jinkela_wire_553;
    wire new_Jinkela_wire_205;
    wire new_Jinkela_wire_841;
    wire new_Jinkela_wire_3165;
    wire new_Jinkela_wire_941;
    wire new_Jinkela_wire_1775;
    wire new_Jinkela_wire_454;
    wire new_Jinkela_wire_698;
    wire new_Jinkela_wire_2922;
    wire _0599_;
    wire new_Jinkela_wire_2613;
    wire _0575_;
    wire new_Jinkela_wire_3065;
    wire new_Jinkela_wire_2872;
    wire _0472_;
    wire new_Jinkela_wire_739;
    wire _0007_;
    wire new_Jinkela_wire_2124;
    wire _0740_;
    wire new_Jinkela_wire_2311;
    wire _0129_;
    wire _0039_;
    wire new_Jinkela_wire_2831;
    wire new_Jinkela_wire_1387;
    wire new_Jinkela_wire_2393;
    wire new_Jinkela_wire_3212;
    wire new_Jinkela_wire_2188;
    wire new_Jinkela_wire_1486;
    wire new_Jinkela_wire_2798;
    wire new_Jinkela_wire_2959;
    wire new_Jinkela_wire_2401;
    wire new_Jinkela_wire_1047;
    wire new_Jinkela_wire_618;
    wire new_Jinkela_wire_597;
    wire new_Jinkela_wire_1597;
    wire new_Jinkela_wire_107;
    wire new_Jinkela_wire_2446;
    wire _0032_;
    wire new_Jinkela_wire_2060;
    wire new_Jinkela_wire_3073;
    wire new_Jinkela_wire_2720;
    wire _0105_;
    wire new_Jinkela_wire_2743;
    wire _0459_;
    wire _0604_;
    wire new_Jinkela_wire_2366;
    wire _0573_;
    wire new_Jinkela_wire_3015;
    wire new_Jinkela_wire_2470;
    wire new_Jinkela_wire_713;
    wire new_Jinkela_wire_2561;
    wire _0794_;
    wire new_Jinkela_wire_230;
    wire _0768_;
    wire new_Jinkela_wire_820;
    wire _0590_;
    wire new_Jinkela_wire_2715;
    wire new_Jinkela_wire_1043;
    wire new_Jinkela_wire_1433;
    wire new_Jinkela_wire_1954;
    wire _0392_;
    wire new_Jinkela_wire_1229;
    wire new_Jinkela_wire_773;
    wire _0216_;
    wire new_Jinkela_wire_1703;
    wire new_Jinkela_wire_237;
    wire new_Jinkela_wire_619;
    wire new_Jinkela_wire_635;
    wire new_Jinkela_wire_2222;
    wire _0666_;
    wire new_Jinkela_wire_961;
    wire new_Jinkela_wire_1984;
    wire new_Jinkela_wire_3186;
    wire new_Jinkela_wire_1538;
    wire _0413_;
    wire new_Jinkela_wire_1900;
    wire _0764_;
    wire new_Jinkela_wire_769;
    wire _0036_;
    wire _0759_;
    wire new_Jinkela_wire_2436;
    wire new_Jinkela_wire_2324;
    wire _0172_;
    wire _0302_;
    wire new_Jinkela_wire_2460;
    wire new_Jinkela_wire_1054;
    wire new_Jinkela_wire_1264;
    wire new_Jinkela_wire_1677;
    wire new_Jinkela_wire_2384;
    wire new_Jinkela_wire_992;
    wire _0288_;
    wire new_Jinkela_wire_186;
    wire new_Jinkela_wire_551;
    wire _0120_;
    wire new_Jinkela_wire_2617;
    wire new_Jinkela_wire_1519;
    wire new_Jinkela_wire_1676;
    wire new_Jinkela_wire_2895;
    wire new_Jinkela_wire_1272;
    wire new_Jinkela_wire_772;
    wire _0058_;
    wire new_Jinkela_wire_3284;
    wire new_Jinkela_wire_339;
    wire new_Jinkela_wire_307;
    wire new_Jinkela_wire_2426;
    wire new_Jinkela_wire_2636;
    wire new_Jinkela_wire_814;
    wire new_Jinkela_wire_671;
    wire new_Jinkela_wire_2534;
    wire _0654_;
    wire new_Jinkela_wire_7;
    wire new_Jinkela_wire_1565;
    wire new_Jinkela_wire_2548;
    wire new_Jinkela_wire_257;
    wire new_Jinkela_wire_3211;
    wire new_Jinkela_wire_2094;
    wire new_Jinkela_wire_2138;
    wire new_Jinkela_wire_2701;
    wire new_Jinkela_wire_2260;
    wire new_Jinkela_wire_2409;
    wire new_Jinkela_wire_2733;
    wire new_Jinkela_wire_3301;
    wire _0278_;
    wire new_Jinkela_wire_2556;
    wire new_Jinkela_wire_754;
    wire new_Jinkela_wire_2382;
    wire new_Jinkela_wire_2238;
    wire new_Jinkela_wire_2081;
    wire _0497_;
    wire _0564_;
    wire new_Jinkela_wire_1651;
    wire new_Jinkela_wire_2965;
    wire new_Jinkela_wire_1217;
    wire new_Jinkela_wire_2185;
    wire new_Jinkela_wire_1854;
    wire new_Jinkela_wire_3058;
    wire new_Jinkela_wire_3260;
    wire new_Jinkela_wire_3150;
    wire new_Jinkela_wire_24;
    wire new_Jinkela_wire_1195;
    wire new_Jinkela_wire_823;
    wire new_Jinkela_wire_3032;
    wire new_Jinkela_wire_1933;
    wire new_Jinkela_wire_1973;
    wire _0377_;
    wire _0161_;
    wire new_Jinkela_wire_2036;
    wire new_Jinkela_wire_1895;
    wire _0692_;
    wire new_Jinkela_wire_881;
    wire new_Jinkela_wire_275;
    wire _0271_;
    wire new_Jinkela_wire_894;
    wire new_Jinkela_wire_399;
    wire new_Jinkela_wire_1708;
    wire new_Jinkela_wire_2609;
    wire new_Jinkela_wire_1236;
    wire new_Jinkela_wire_1080;
    wire _0533_;
    wire new_Jinkela_wire_2652;
    wire new_Jinkela_wire_455;
    wire new_Jinkela_wire_2724;
    wire new_Jinkela_wire_1363;
    wire new_Jinkela_wire_1547;
    wire _0235_;
    wire new_Jinkela_wire_2948;
    wire new_Jinkela_wire_2683;
    wire new_Jinkela_wire_2112;
    wire new_Jinkela_wire_2568;
    wire _0427_;
    wire new_Jinkela_wire_1391;
    wire new_Jinkela_wire_1846;
    wire _0181_;
    wire new_Jinkela_wire_228;
    wire new_Jinkela_wire_2158;
    wire new_Jinkela_wire_2946;
    wire new_Jinkela_wire_340;
    wire new_Jinkela_wire_1261;
    wire new_Jinkela_wire_1268;
    wire new_Jinkela_wire_522;
    wire new_Jinkela_wire_3018;
    wire new_Jinkela_wire_3118;
    wire new_Jinkela_wire_1075;
    wire _0544_;
    wire new_Jinkela_wire_3069;
    wire _0063_;
    wire new_Jinkela_wire_1104;
    wire _0707_;
    wire new_Jinkela_wire_2546;
    wire new_Jinkela_wire_2545;
    wire new_Jinkela_wire_1035;
    wire new_Jinkela_wire_897;
    wire _0677_;
    wire new_Jinkela_wire_3101;
    wire _0262_;
    wire new_Jinkela_wire_2491;
    wire _0227_;
    wire new_Jinkela_wire_3024;
    wire new_Jinkela_wire_1847;
    wire new_Jinkela_wire_1974;
    wire new_Jinkela_wire_1393;
    wire new_Jinkela_wire_2845;
    wire new_Jinkela_wire_3283;
    wire new_Jinkela_wire_1352;
    wire new_Jinkela_wire_624;
    wire new_Jinkela_wire_3219;
    wire new_Jinkela_wire_1544;
    wire new_Jinkela_wire_1180;
    wire new_Jinkela_wire_2096;
    wire _0043_;
    wire new_Jinkela_wire_1618;
    wire new_net_7;
    wire new_Jinkela_wire_679;
    wire _0797_;
    wire new_Jinkela_wire_471;
    wire new_Jinkela_wire_3017;
    wire new_Jinkela_wire_2532;
    wire new_Jinkela_wire_3270;
    wire new_Jinkela_wire_56;
    wire new_Jinkela_wire_1196;
    wire _0016_;
    wire new_Jinkela_wire_2775;
    wire new_net_1467;
    wire new_Jinkela_wire_227;
    wire _0449_;
    wire new_Jinkela_wire_2156;
    wire _0601_;
    wire new_Jinkela_wire_2437;
    wire new_Jinkela_wire_3296;
    wire new_Jinkela_wire_49;
    wire new_Jinkela_wire_2689;
    wire new_Jinkela_wire_3199;
    wire new_Jinkela_wire_1924;
    wire _0483_;
    wire new_Jinkela_wire_1890;
    wire new_Jinkela_wire_1012;
    wire _0371_;
    wire _0770_;
    wire new_Jinkela_wire_1566;
    wire new_Jinkela_wire_2201;
    wire new_Jinkela_wire_999;
    wire new_Jinkela_wire_2383;
    wire new_Jinkela_wire_1452;
    wire new_Jinkela_wire_3181;
    wire new_Jinkela_wire_2135;
    wire new_Jinkela_wire_1403;
    wire new_Jinkela_wire_2495;
    wire _0014_;
    wire new_Jinkela_wire_2090;
    wire new_Jinkela_wire_249;
    wire new_Jinkela_wire_1628;
    wire new_Jinkela_wire_2840;
    wire _0083_;
    wire new_Jinkela_wire_628;
    wire new_Jinkela_wire_2214;
    wire new_Jinkela_wire_2637;
    wire new_Jinkela_wire_558;
    wire new_Jinkela_wire_1937;
    wire new_Jinkela_wire_362;
    wire new_Jinkela_wire_60;
    wire new_Jinkela_wire_441;
    wire _0372_;
    wire new_Jinkela_wire_3328;
    wire new_Jinkela_wire_1071;
    wire new_Jinkela_wire_478;
    wire _0468_;
    wire new_Jinkela_wire_2471;
    wire new_Jinkela_wire_701;
    wire new_Jinkela_wire_1869;
    wire new_Jinkela_wire_2114;
    wire _0504_;
    wire new_Jinkela_wire_1245;
    wire new_Jinkela_wire_3140;
    wire new_Jinkela_wire_2452;
    wire new_Jinkela_wire_784;
    wire new_Jinkela_wire_29;
    wire new_Jinkela_wire_3113;
    wire new_Jinkela_wire_379;
    wire new_Jinkela_wire_3274;
    wire new_Jinkela_wire_2601;
    wire new_Jinkela_wire_2851;
    wire new_Jinkela_wire_1851;
    wire new_Jinkela_wire_3129;
    wire new_Jinkela_wire_2644;
    wire new_Jinkela_wire_1988;
    wire new_Jinkela_wire_337;
    wire new_Jinkela_wire_885;
    wire new_Jinkela_wire_274;
    wire _0595_;
    wire new_Jinkela_wire_2630;
    wire _0260_;
    wire new_Jinkela_wire_223;
    wire new_Jinkela_wire_1262;
    wire new_Jinkela_wire_398;
    wire new_Jinkela_wire_222;
    wire _0292_;
    wire new_Jinkela_wire_3022;
    wire new_Jinkela_wire_1304;
    wire new_Jinkela_wire_1696;
    wire new_Jinkela_wire_1783;
    wire new_Jinkela_wire_2440;
    wire new_Jinkela_wire_3052;
    wire new_Jinkela_wire_344;
    wire new_Jinkela_wire_2351;
    wire new_Jinkela_wire_3259;
    wire new_Jinkela_wire_2807;
    wire new_Jinkela_wire_2422;
    wire _0520_;
    wire new_Jinkela_wire_1513;
    wire new_Jinkela_wire_1318;
    wire new_Jinkela_wire_58;
    wire _0616_;
    wire new_Jinkela_wire_2051;
    wire new_Jinkela_wire_2620;
    wire new_Jinkela_wire_290;
    wire new_Jinkela_wire_295;
    wire new_Jinkela_wire_717;
    wire new_Jinkela_wire_2093;
    wire new_Jinkela_wire_1517;
    wire _0359_;
    wire new_Jinkela_wire_1423;
    wire new_Jinkela_wire_2381;
    wire new_Jinkela_wire_1305;
    wire new_Jinkela_wire_1311;
    wire new_Jinkela_wire_1769;
    wire new_Jinkela_wire_1788;
    wire _0421_;
    wire _0326_;
    wire new_Jinkela_wire_1896;
    wire new_Jinkela_wire_807;
    wire new_Jinkela_wire_2207;
    wire new_Jinkela_wire_2176;
    wire new_Jinkela_wire_1809;
    wire new_Jinkela_wire_1707;
    wire new_Jinkela_wire_1705;
    wire _0384_;
    wire _0367_;
    wire _0745_;
    wire new_Jinkela_wire_1802;
    wire new_Jinkela_wire_994;
    wire new_Jinkela_wire_950;
    wire new_Jinkela_wire_9;
    wire new_Jinkela_wire_951;
    wire new_Jinkela_wire_2590;
    wire _0465_;
    wire new_Jinkela_wire_2368;
    wire new_Jinkela_wire_380;
    wire new_Jinkela_wire_298;
    wire new_Jinkela_wire_1557;
    wire new_Jinkela_wire_911;
    wire new_Jinkela_wire_1608;
    wire _0093_;
    wire new_Jinkela_wire_662;
    wire _0546_;
    wire _0042_;
    wire new_Jinkela_wire_876;
    wire new_Jinkela_wire_326;
    wire new_Jinkela_wire_700;
    wire new_Jinkela_wire_2821;
    wire new_Jinkela_wire_2217;
    wire new_Jinkela_wire_1611;
    wire new_Jinkela_wire_2206;
    wire new_Jinkela_wire_1490;
    wire _0351_;
    wire new_Jinkela_wire_1331;
    wire new_Jinkela_wire_395;
    wire _0049_;
    wire new_Jinkela_wire_2289;
    wire new_Jinkela_wire_184;
    wire new_Jinkela_wire_1179;
    wire new_Jinkela_wire_2790;
    wire _0771_;
    wire new_Jinkela_wire_2448;
    wire new_Jinkela_wire_695;
    wire new_Jinkela_wire_2190;
    wire new_Jinkela_wire_1524;
    wire new_Jinkela_wire_705;
    wire new_Jinkela_wire_2978;
    wire new_Jinkela_wire_145;
    wire _0670_;
    wire new_Jinkela_wire_1431;
    wire new_Jinkela_wire_312;
    wire _0474_;
    wire new_Jinkela_wire_1841;
    wire new_Jinkela_wire_2469;
    wire new_Jinkela_wire_1372;
    wire new_Jinkela_wire_260;
    wire new_Jinkela_wire_1849;
    wire new_Jinkela_wire_565;
    wire new_Jinkela_wire_2897;
    wire new_Jinkela_wire_843;
    wire new_Jinkela_wire_1965;
    wire new_Jinkela_wire_826;
    wire new_Jinkela_wire_2163;
    wire new_Jinkela_wire_1240;
    wire new_Jinkela_wire_1333;
    wire _0331_;
    wire new_Jinkela_wire_2427;
    wire new_Jinkela_wire_3051;
    wire _0165_;
    wire new_Jinkela_wire_204;
    wire new_Jinkela_wire_2765;
    wire _0580_;
    wire new_Jinkela_wire_563;
    wire new_Jinkela_wire_341;
    wire new_Jinkela_wire_2160;
    wire new_Jinkela_wire_2468;
    wire new_Jinkela_wire_2924;
    wire _0158_;
    wire _0184_;
    wire new_Jinkela_wire_1754;
    wire new_net_1485;
    wire new_Jinkela_wire_998;
    wire _0149_;
    wire new_Jinkela_wire_2991;
    wire _0559_;
    wire new_Jinkela_wire_16;
    wire new_Jinkela_wire_1132;
    wire _0232_;
    wire new_Jinkela_wire_2972;
    wire new_Jinkela_wire_1604;
    wire _0357_;
    wire _0026_;
    wire _0786_;
    wire _0500_;
    wire new_Jinkela_wire_1414;
    wire new_Jinkela_wire_1744;
    wire new_Jinkela_wire_2810;
    wire new_Jinkela_wire_1975;
    wire new_Jinkela_wire_614;
    wire new_Jinkela_wire_1336;
    wire new_Jinkela_wire_3281;
    wire new_Jinkela_wire_64;
    wire new_Jinkela_wire_2671;
    wire new_Jinkela_wire_887;
    wire new_Jinkela_wire_674;
    wire new_Jinkela_wire_2358;
    wire new_Jinkela_wire_1356;
    wire new_Jinkela_wire_466;
    wire new_Jinkela_wire_1674;
    wire new_Jinkela_wire_591;
    wire new_Jinkela_wire_2209;
    wire new_Jinkela_wire_570;
    wire new_Jinkela_wire_1867;
    wire new_Jinkela_wire_2662;
    wire _0735_;
    wire new_Jinkela_wire_2137;
    wire new_Jinkela_wire_2357;
    wire new_Jinkela_wire_697;
    wire new_Jinkela_wire_1667;
    wire new_Jinkela_wire_901;
    wire new_Jinkela_wire_211;
    wire new_Jinkela_wire_3060;
    wire new_Jinkela_wire_2507;
    wire new_Jinkela_wire_1860;
    wire new_Jinkela_wire_1522;
    wire new_Jinkela_wire_3325;
    wire _0244_;
    wire new_Jinkela_wire_2789;
    wire new_Jinkela_wire_3177;
    wire new_Jinkela_wire_2053;
    wire new_Jinkela_wire_2338;
    wire new_Jinkela_wire_1599;
    wire new_Jinkela_wire_46;
    wire new_Jinkela_wire_1941;
    wire new_Jinkela_wire_288;
    wire new_Jinkela_wire_90;
    wire new_Jinkela_wire_1959;
    wire new_Jinkela_wire_414;
    wire new_Jinkela_wire_1586;
    wire new_Jinkela_wire_2276;
    wire _0558_;
    wire new_Jinkela_wire_1889;
    wire _0234_;
    wire _0691_;
    wire new_Jinkela_wire_3169;
    wire _0263_;
    wire new_Jinkela_wire_1653;
    wire new_Jinkela_wire_1446;
    wire new_Jinkela_wire_2850;
    wire new_Jinkela_wire_1198;
    wire new_Jinkela_wire_1953;
    wire _0349_;
    wire _0004_;
    wire _0360_;
    wire new_Jinkela_wire_2802;
    wire new_Jinkela_wire_358;
    wire new_Jinkela_wire_2905;
    wire new_Jinkela_wire_351;
    wire _0088_;
    wire new_Jinkela_wire_3184;
    wire new_Jinkela_wire_408;
    wire new_Jinkela_wire_1770;
    wire new_Jinkela_wire_2012;
    wire new_Jinkela_wire_1142;
    wire _0772_;
    wire new_Jinkela_wire_375;
    wire new_Jinkela_wire_276;
    wire _0715_;
    wire new_Jinkela_wire_2686;
    wire _0646_;
    wire _0749_;
    wire new_Jinkela_wire_1366;
    wire new_Jinkela_wire_1357;
    wire new_Jinkela_wire_3059;
    wire _0644_;
    wire new_Jinkela_wire_656;
    wire new_Jinkela_wire_1377;
    wire _0763_;
    wire new_Jinkela_wire_1606;
    wire new_Jinkela_wire_1873;
    wire new_Jinkela_wire_2560;
    wire _0177_;
    wire new_Jinkela_wire_1550;
    wire new_Jinkela_wire_1337;
    wire _0620_;
    wire new_Jinkela_wire_3011;
    wire new_Jinkela_wire_2852;
    wire new_Jinkela_wire_2508;
    wire new_Jinkela_wire_2650;
    wire new_Jinkela_wire_542;
    wire new_Jinkela_wire_1116;
    wire new_Jinkela_wire_2778;
    wire new_Jinkela_wire_138;
    wire new_Jinkela_wire_418;
    wire new_Jinkela_wire_346;
    wire new_Jinkela_wire_917;
    wire new_Jinkela_wire_1644;
    wire new_Jinkela_wire_742;
    wire new_Jinkela_wire_435;
    wire new_Jinkela_wire_2226;
    wire new_Jinkela_wire_1562;
    wire _0549_;
    wire new_Jinkela_wire_30;
    wire new_Jinkela_wire_3000;
    wire new_Jinkela_wire_1572;
    wire _0127_;
    wire new_Jinkela_wire_1224;
    wire new_Jinkela_wire_1254;
    wire new_Jinkela_wire_1831;
    wire new_Jinkela_wire_2466;
    wire new_Jinkela_wire_1848;
    wire new_Jinkela_wire_2191;
    wire new_Jinkela_wire_2113;
    wire new_Jinkela_wire_711;
    wire new_Jinkela_wire_1188;
    wire new_Jinkela_wire_208;
    wire _0552_;
    wire new_Jinkela_wire_3046;
    wire new_Jinkela_wire_236;
    wire new_Jinkela_wire_2569;
    wire new_Jinkela_wire_1814;
    wire new_Jinkela_wire_1897;
    wire _0611_;
    wire new_Jinkela_wire_133;
    wire new_Jinkela_wire_2242;
    wire _0716_;
    wire new_Jinkela_wire_266;
    wire new_Jinkela_wire_451;
    wire new_Jinkela_wire_2935;
    wire new_Jinkela_wire_378;
    wire new_Jinkela_wire_2640;
    wire new_Jinkela_wire_1722;
    wire new_Jinkela_wire_1473;
    wire new_Jinkela_wire_2369;
    wire new_Jinkela_wire_2877;
    wire _0168_;
    wire new_Jinkela_wire_1185;
    wire new_Jinkela_wire_2414;
    wire new_Jinkela_wire_1502;
    wire new_Jinkela_wire_2949;
    wire new_Jinkela_wire_1946;
    wire new_Jinkela_wire_2512;
    wire new_Jinkela_wire_2673;
    wire new_Jinkela_wire_1292;
    wire new_Jinkela_wire_1308;
    wire new_Jinkela_wire_730;
    wire new_Jinkela_wire_1488;
    wire new_Jinkela_wire_59;
    wire new_Jinkela_wire_1575;
    wire new_Jinkela_wire_575;
    wire new_Jinkela_wire_2227;
    wire _0332_;
    wire new_Jinkela_wire_3091;
    wire new_Jinkela_wire_97;
    wire _0130_;
    wire new_Jinkela_wire_744;
    wire _0789_;
    wire _0507_;
    wire new_Jinkela_wire_2914;
    wire new_Jinkela_wire_1535;
    wire new_Jinkela_wire_80;
    wire new_Jinkela_wire_2480;
    wire new_Jinkela_wire_256;
    wire new_Jinkela_wire_544;
    wire new_Jinkela_wire_2859;
    wire new_Jinkela_wire_2402;
    wire new_Jinkela_wire_3172;
    wire _0065_;
    wire new_Jinkela_wire_620;
    wire new_Jinkela_wire_706;
    wire _0695_;
    wire new_Jinkela_wire_1857;
    wire new_Jinkela_wire_2443;
    wire _0040_;
    wire new_Jinkela_wire_2306;
    wire new_Jinkela_wire_2917;
    wire new_Jinkela_wire_827;
    wire _0785_;
    wire new_Jinkela_wire_983;
    wire new_Jinkela_wire_1219;
    wire _0356_;
    wire _0733_;
    wire new_Jinkela_wire_3014;
    wire new_Jinkela_wire_1063;
    wire _0152_;
    wire new_Jinkela_wire_55;
    wire new_Jinkela_wire_169;
    wire new_Jinkela_wire_1145;
    wire new_Jinkela_wire_2976;
    wire new_Jinkela_wire_128;
    wire new_Jinkela_wire_3019;
    wire _0650_;
    wire new_Jinkela_wire_1919;
    wire new_Jinkela_wire_1020;
    wire new_Jinkela_wire_2292;
    wire new_Jinkela_wire_318;
    wire new_Jinkela_wire_878;
    wire new_Jinkela_wire_1161;
    wire new_Jinkela_wire_86;
    wire new_Jinkela_wire_2760;
    wire _0401_;
    wire new_Jinkela_wire_2011;
    wire new_Jinkela_wire_668;
    wire new_Jinkela_wire_1856;
    wire new_Jinkela_wire_2492;
    wire new_Jinkela_wire_2101;
    wire new_Jinkela_wire_2280;
    wire new_Jinkela_wire_1349;
    wire new_Jinkela_wire_1275;
    wire new_Jinkela_wire_3041;
    wire new_Jinkela_wire_937;
    wire new_Jinkela_wire_2428;
    wire _0452_;
    wire new_net_1477;
    wire new_Jinkela_wire_388;
    wire new_Jinkela_wire_2956;
    wire new_Jinkela_wire_594;
    wire new_Jinkela_wire_1233;
    wire new_Jinkela_wire_1113;
    wire _0071_;
    wire new_Jinkela_wire_2223;
    wire _0412_;
    wire new_Jinkela_wire_1482;
    wire new_Jinkela_wire_2052;
    wire new_Jinkela_wire_906;
    wire _0052_;
    wire new_Jinkela_wire_245;
    wire new_Jinkela_wire_2577;
    wire new_Jinkela_wire_1440;
    wire new_Jinkela_wire_415;
    wire _0212_;
    wire _0430_;
    wire new_Jinkela_wire_1504;
    wire new_Jinkela_wire_3141;
    wire new_Jinkela_wire_2835;
    wire new_Jinkela_wire_2981;
    wire new_Jinkela_wire_865;
    wire new_Jinkela_wire_229;
    wire new_Jinkela_wire_1994;
    wire new_Jinkela_wire_2586;
    wire new_Jinkela_wire_387;
    wire new_Jinkela_wire_70;
    wire new_Jinkela_wire_73;
    wire new_Jinkela_wire_2531;
    wire new_Jinkela_wire_1248;
    wire _0213_;
    wire new_Jinkela_wire_2980;
    wire new_Jinkela_wire_2462;
    wire new_Jinkela_wire_1322;
    wire new_Jinkela_wire_1658;
    wire new_Jinkela_wire_1216;
    wire new_Jinkela_wire_1922;
    wire new_Jinkela_wire_2788;
    wire new_Jinkela_wire_2396;
    wire new_Jinkela_wire_785;
    wire new_Jinkela_wire_1394;
    wire new_Jinkela_wire_513;
    wire new_Jinkela_wire_2353;
    wire new_Jinkela_wire_2658;
    wire _0237_;
    wire new_Jinkela_wire_1277;
    wire new_Jinkela_wire_1215;
    wire new_Jinkela_wire_1014;
    wire new_Jinkela_wire_422;
    wire new_Jinkela_wire_3163;
    wire _0778_;
    wire new_Jinkela_wire_2102;
    wire new_Jinkela_wire_1601;
    wire new_net_1473;
    wire new_Jinkela_wire_3161;
    wire new_Jinkela_wire_1605;
    wire new_Jinkela_wire_2048;
    wire new_Jinkela_wire_76;
    wire new_Jinkela_wire_87;
    wire new_Jinkela_wire_1957;
    wire _0539_;
    wire new_Jinkela_wire_2762;
    wire _0198_;
    wire new_Jinkela_wire_2942;
    wire new_Jinkela_wire_2275;
    wire new_Jinkela_wire_1329;
    wire new_Jinkela_wire_1728;
    wire new_Jinkela_wire_3299;
    wire new_Jinkela_wire_1878;
    wire new_Jinkela_wire_185;
    wire new_Jinkela_wire_279;
    wire _0286_;
    wire new_Jinkela_wire_535;
    wire new_Jinkela_wire_2360;
    wire new_Jinkela_wire_2125;
    wire new_Jinkela_wire_640;
    wire new_Jinkela_wire_1341;
    wire new_Jinkela_wire_723;
    wire new_Jinkela_wire_508;
    wire new_Jinkela_wire_732;
    wire new_Jinkela_wire_2456;
    wire _0193_;
    wire new_Jinkela_wire_1531;
    wire _0431_;
    wire new_Jinkela_wire_173;
    wire new_Jinkela_wire_2246;
    wire new_Jinkela_wire_2605;
    wire new_Jinkela_wire_1203;
    wire new_Jinkela_wire_1622;
    wire new_Jinkela_wire_1193;
    wire new_Jinkela_wire_2365;
    wire new_Jinkela_wire_335;
    wire _0267_;
    wire new_Jinkela_wire_79;
    wire new_Jinkela_wire_3152;
    wire new_Jinkela_wire_2903;
    wire new_Jinkela_wire_987;
    wire new_Jinkela_wire_680;
    wire new_Jinkela_wire_1051;
    wire _0623_;
    wire _0210_;
    wire new_Jinkela_wire_2977;
    wire new_Jinkela_wire_36;
    wire new_Jinkela_wire_2145;
    wire new_Jinkela_wire_1901;
    wire new_Jinkela_wire_2611;
    wire new_Jinkela_wire_561;
    wire new_Jinkela_wire_2449;
    wire new_Jinkela_wire_2169;
    wire new_Jinkela_wire_2331;
    wire new_Jinkela_wire_2344;
    wire new_Jinkela_wire_2882;
    wire new_Jinkela_wire_3329;
    wire new_Jinkela_wire_3313;
    wire _0479_;
    wire new_Jinkela_wire_790;
    wire new_Jinkela_wire_1515;
    wire new_Jinkela_wire_1713;
    wire new_Jinkela_wire_2299;
    wire new_Jinkela_wire_3021;
    wire _0226_;
    wire _0617_;
    wire new_Jinkela_wire_642;
    wire new_Jinkela_wire_2691;
    wire new_Jinkela_wire_2183;
    wire new_Jinkela_wire_1740;
    wire _0501_;
    wire _0592_;
    wire new_Jinkela_wire_1778;
    wire new_Jinkela_wire_733;
    wire new_Jinkela_wire_1661;
    wire new_Jinkela_wire_347;
    wire new_Jinkela_wire_3123;
    wire new_Jinkela_wire_877;
    wire new_Jinkela_wire_1191;
    wire new_Jinkela_wire_1354;
    wire new_Jinkela_wire_3095;
    wire new_Jinkela_wire_2916;
    wire new_Jinkela_wire_2079;
    wire new_Jinkela_wire_1871;
    wire _0524_;
    wire new_Jinkela_wire_675;
    wire new_Jinkela_wire_1731;
    wire new_Jinkela_wire_689;
    wire new_Jinkela_wire_669;
    wire _0285_;
    wire new_Jinkela_wire_1561;
    wire new_Jinkela_wire_2334;
    wire new_Jinkela_wire_1266;
    wire _0222_;
    wire new_Jinkela_wire_2540;
    wire new_Jinkela_wire_371;
    wire _0570_;
    wire new_Jinkela_wire_2651;
    wire new_Jinkela_wire_2106;
    wire new_Jinkela_wire_1127;
    wire new_Jinkela_wire_2153;
    wire new_Jinkela_wire_2869;
    wire new_Jinkela_wire_2915;
    wire _0517_;
    wire new_Jinkela_wire_3238;
    wire new_Jinkela_wire_2062;
    wire new_Jinkela_wire_3282;
    wire new_Jinkela_wire_1687;
    wire _0146_;
    wire new_Jinkela_wire_2148;
    wire new_Jinkela_wire_2259;
    wire new_Jinkela_wire_1943;
    wire new_Jinkela_wire_1785;
    wire _0741_;
    wire _0603_;
    wire new_Jinkela_wire_2343;
    wire new_Jinkela_wire_1120;
    wire new_Jinkela_wire_1526;
    wire _0269_;
    wire new_Jinkela_wire_2364;
    wire new_Jinkela_wire_3009;
    wire _0561_;
    wire new_Jinkela_wire_278;
    wire _0642_;
    wire new_Jinkela_wire_2716;
    wire new_Jinkela_wire_2742;
    wire new_Jinkela_wire_2538;
    wire new_Jinkela_wire_1880;
    wire _0565_;
    wire new_Jinkela_wire_2415;
    wire new_Jinkela_wire_2390;
    wire new_Jinkela_wire_1209;
    wire new_Jinkela_wire_1009;
    wire new_Jinkela_wire_3215;
    wire new_Jinkela_wire_1972;
    wire _0113_;
    wire new_Jinkela_wire_1485;
    wire new_Jinkela_wire_1257;
    wire new_Jinkela_wire_180;
    wire new_Jinkela_wire_623;
    wire new_Jinkela_wire_93;
    wire new_Jinkela_wire_851;
    wire new_Jinkela_wire_2934;
    wire new_Jinkela_wire_2405;
    wire new_Jinkela_wire_137;
    wire _0208_;
    wire new_Jinkela_wire_269;
    wire new_Jinkela_wire_2714;
    wire new_Jinkela_wire_2117;
    wire new_Jinkela_wire_2675;
    wire new_Jinkela_wire_3290;
    wire new_Jinkela_wire_2908;
    wire new_Jinkela_wire_2827;
    wire new_Jinkela_wire_2626;
    wire new_Jinkela_wire_2195;
    wire _0634_;
    wire new_Jinkela_wire_1654;
    wire new_Jinkela_wire_1600;
    wire new_Jinkela_wire_2927;
    wire new_Jinkela_wire_1634;
    wire _0010_;
    wire new_net_0;
    wire _0477_;
    wire new_Jinkela_wire_448;
    wire new_Jinkela_wire_3200;
    wire new_Jinkela_wire_3205;
    wire new_Jinkela_wire_1763;
    wire _0009_;
    wire _0050_;
    wire _0200_;
    wire new_Jinkela_wire_3016;
    wire new_Jinkela_wire_529;
    wire new_Jinkela_wire_515;
    wire _0795_;
    wire new_Jinkela_wire_308;
    wire new_Jinkela_wire_1400;
    wire new_Jinkela_wire_631;
    wire new_Jinkela_wire_261;
    wire new_Jinkela_wire_2585;
    wire _0630_;
    wire new_Jinkela_wire_1796;
    wire new_Jinkela_wire_2619;
    wire new_Jinkela_wire_289;
    wire new_Jinkela_wire_2833;
    wire new_Jinkela_wire_1571;
    wire new_Jinkela_wire_1206;
    wire new_Jinkela_wire_1534;
    wire new_Jinkela_wire_1199;
    wire new_Jinkela_wire_1807;
    wire new_Jinkela_wire_2404;
    wire new_Jinkela_wire_3025;
    wire new_Jinkela_wire_2632;
    wire new_Jinkela_wire_1475;
    wire _0396_;
    wire _0767_;
    wire new_Jinkela_wire_389;
    wire new_Jinkela_wire_3190;
    wire _0388_;
    wire _0167_;
    wire _0777_;
    wire new_Jinkela_wire_799;
    wire new_Jinkela_wire_2004;
    wire _0436_;
    wire new_Jinkela_wire_804;
    wire new_Jinkela_wire_965;
    wire _0304_;
    wire new_Jinkela_wire_3320;
    wire new_Jinkela_wire_89;
    wire new_Jinkela_wire_25;
    wire new_Jinkela_wire_1444;
    wire _0176_;
    wire _0219_;
    wire new_Jinkela_wire_2078;
    wire new_Jinkela_wire_1344;
    wire new_Jinkela_wire_1285;
    wire new_Jinkela_wire_2853;
    wire _0137_;
    wire new_Jinkela_wire_2878;
    wire _0314_;
    wire new_Jinkela_wire_1755;
    wire _0380_;
    wire new_Jinkela_wire_2316;
    wire new_Jinkela_wire_2115;
    wire new_Jinkela_wire_1607;
    wire new_Jinkela_wire_912;
    wire new_Jinkela_wire_2930;
    wire _0041_;
    wire new_Jinkela_wire_1057;
    wire new_Jinkela_wire_644;
    wire _0361_;
    wire _0613_;
    wire new_Jinkela_wire_3170;
    wire new_Jinkela_wire_458;
    wire _0154_;
    wire new_Jinkela_wire_2376;
    wire new_Jinkela_wire_1374;
    wire new_Jinkela_wire_2841;
    wire _0275_;
    wire new_Jinkela_wire_2476;
    wire new_Jinkela_wire_3010;
    wire new_Jinkela_wire_1536;
    wire new_Jinkela_wire_2398;
    wire new_Jinkela_wire_900;
    wire new_Jinkela_wire_1086;
    wire new_Jinkela_wire_1004;
    wire new_Jinkela_wire_248;
    wire _0284_;
    wire new_Jinkela_wire_886;
    wire new_Jinkela_wire_655;
    wire new_Jinkela_wire_550;
    wire new_Jinkela_wire_1518;
    wire new_Jinkela_wire_1320;
    wire new_Jinkela_wire_193;
    wire new_Jinkela_wire_1361;
    wire new_Jinkela_wire_239;
    wire new_Jinkela_wire_3250;
    wire new_Jinkela_wire_608;
    wire new_Jinkela_wire_1964;
    wire new_Jinkela_wire_2400;
    wire new_Jinkela_wire_555;
    wire _0368_;
    wire new_Jinkela_wire_775;
    wire new_Jinkela_wire_1932;
    wire new_Jinkela_wire_2963;
    wire new_Jinkela_wire_2741;
    wire new_Jinkela_wire_3131;
    wire _0087_;
    wire new_Jinkela_wire_750;
    wire new_Jinkela_wire_2228;
    wire new_Jinkela_wire_334;
    wire new_Jinkela_wire_2684;
    wire new_Jinkela_wire_3178;
    wire new_Jinkela_wire_1424;
    wire new_Jinkela_wire_3331;
    wire new_Jinkela_wire_1640;
    wire new_Jinkela_wire_3105;
    wire new_Jinkela_wire_1799;
    wire new_Jinkela_wire_891;
    wire new_Jinkela_wire_1105;
    wire new_Jinkela_wire_301;
    wire new_Jinkela_wire_2635;
    wire new_Jinkela_wire_1426;
    wire new_Jinkela_wire_1759;
    wire _0526_;
    wire new_Jinkela_wire_2870;
    wire new_Jinkela_wire_796;
    wire new_Jinkela_wire_2278;
    wire _0481_;
    wire new_Jinkela_wire_2355;
    wire _0089_;
    wire _0408_;
    wire _0341_;
    wire new_Jinkela_wire_3237;
    wire new_Jinkela_wire_3125;
    wire new_Jinkela_wire_1647;
    wire _0752_;
    wire new_Jinkela_wire_2150;
    wire new_Jinkela_wire_2084;
    wire new_Jinkela_wire_1416;
    wire new_Jinkela_wire_2107;
    wire new_Jinkela_wire_1273;
    wire new_Jinkela_wire_835;
    wire _0682_;
    wire new_Jinkela_wire_1887;
    wire new_Jinkela_wire_1143;
    wire new_Jinkela_wire_203;
    wire _0189_;
    wire new_Jinkela_wire_3127;
    wire _0381_;
    wire new_Jinkela_wire_1693;
    wire _0280_;
    wire _0229_;
    wire new_Jinkela_wire_533;
    wire new_Jinkela_wire_1747;
    wire _0696_;
    wire new_Jinkela_wire_1246;
    wire new_Jinkela_wire_1176;
    wire new_Jinkela_wire_2434;
    wire new_Jinkela_wire_2411;
    wire new_Jinkela_wire_2511;
    wire new_Jinkela_wire_2371;
    wire new_Jinkela_wire_2979;
    wire new_Jinkela_wire_2046;
    wire new_Jinkela_wire_2417;
    wire new_Jinkela_wire_602;
    wire new_Jinkela_wire_1454;
    wire new_Jinkela_wire_1259;
    wire new_Jinkela_wire_1619;
    wire new_Jinkela_wire_131;
    wire _0013_;
    wire new_Jinkela_wire_2123;
    wire new_Jinkela_wire_2304;
    wire new_Jinkela_wire_1359;
    wire _0029_;
    wire new_Jinkela_wire_1990;
    wire new_Jinkela_wire_792;
    wire _0461_;
    wire _0252_;
    wire _0525_;
    wire new_Jinkela_wire_21;
    wire new_Jinkela_wire_1052;
    wire _0206_;
    wire new_Jinkela_wire_2627;
    wire new_Jinkela_wire_1293;
    wire new_Jinkela_wire_1580;
    wire new_Jinkela_wire_1592;
    wire new_Jinkela_wire_1376;
    wire new_Jinkela_wire_117;
    wire new_Jinkela_wire_2031;
    wire new_Jinkela_wire_2087;
    wire new_Jinkela_wire_566;
    wire new_Jinkela_wire_2317;
    wire new_Jinkela_wire_2202;
    wire new_Jinkela_wire_35;
    wire new_Jinkela_wire_617;
    wire _0192_;
    wire new_Jinkela_wire_3171;
    wire new_Jinkela_wire_443;
    wire new_Jinkela_wire_258;
    wire new_Jinkela_wire_858;
    wire _0674_;
    wire new_Jinkela_wire_420;
    wire new_Jinkela_wire_2873;
    wire new_Jinkela_wire_2337;
    wire new_Jinkela_wire_1552;
    wire new_Jinkela_wire_1235;
    wire new_Jinkela_wire_2342;
    wire new_Jinkela_wire_1389;
    wire new_Jinkela_wire_847;
    wire _0543_;
    wire new_Jinkela_wire_1030;
    wire new_Jinkela_wire_2952;
    wire _0582_;
    wire new_Jinkela_wire_722;
    wire new_Jinkela_wire_370;
    wire _0217_;
    wire _0005_;
    wire new_Jinkela_wire_907;
    wire new_Jinkela_wire_1310;
    wire new_Jinkela_wire_997;
    wire new_Jinkela_wire_2902;
    wire new_Jinkela_wire_1692;
    wire new_Jinkela_wire_1623;
    wire new_Jinkela_wire_1520;
    wire new_Jinkela_wire_1563;
    wire new_Jinkela_wire_2519;
    wire new_Jinkela_wire_1553;
    wire _0289_;
    wire new_Jinkela_wire_331;
    wire new_Jinkela_wire_479;
    wire new_Jinkela_wire_605;
    wire new_Jinkela_wire_2829;
    wire new_Jinkela_wire_71;
    wire _0019_;
    wire new_Jinkela_wire_2229;
    wire new_Jinkela_wire_1325;
    wire new_Jinkela_wire_1072;
    wire new_Jinkela_wire_2178;
    wire new_Jinkela_wire_40;
    wire new_Jinkela_wire_300;
    wire new_Jinkela_wire_2136;
    wire new_Jinkela_wire_2708;
    wire new_Jinkela_wire_3303;
    wire _0256_;
    wire new_Jinkela_wire_3209;
    wire new_Jinkela_wire_5;
    wire new_Jinkela_wire_1456;
    wire _0584_;
    wire new_Jinkela_wire_1214;
    wire new_Jinkela_wire_263;
    wire _0469_;
    wire new_Jinkela_wire_2711;
    wire new_Jinkela_wire_156;
    wire new_Jinkela_wire_1983;
    wire new_Jinkela_wire_798;
    wire new_Jinkela_wire_1383;
    wire new_Jinkela_wire_2420;
    wire new_Jinkela_wire_1603;
    wire _0124_;
    wire new_Jinkela_wire_1913;
    wire new_Jinkela_wire_1942;
    wire new_Jinkela_wire_2445;
    wire _0671_;
    wire new_Jinkela_wire_2213;
    wire new_Jinkela_wire_2378;
    wire new_Jinkela_wire_806;
    wire new_Jinkela_wire_3176;
    wire new_Jinkela_wire_197;
    wire new_Jinkela_wire_1494;
    wire _0522_;
    wire _0374_;
    wire new_Jinkela_wire_3251;
    wire new_Jinkela_wire_1290;
    wire new_Jinkela_wire_2302;
    wire _0643_;
    wire new_Jinkela_wire_1384;
    wire new_Jinkela_wire_2994;
    wire new_Jinkela_wire_1062;
    wire new_Jinkela_wire_1067;
    wire new_Jinkela_wire_1346;
    wire _0264_;
    wire _0246_;
    wire new_Jinkela_wire_788;
    wire new_Jinkela_wire_181;
    wire _0627_;
    wire new_Jinkela_wire_1150;
    wire new_Jinkela_wire_776;
    wire new_Jinkela_wire_2964;
    wire new_Jinkela_wire_836;
    wire new_Jinkela_wire_1980;
    wire new_Jinkela_wire_3236;
    wire new_Jinkela_wire_2631;
    wire new_Jinkela_wire_1716;
    wire new_Jinkela_wire_509;
    wire new_Jinkela_wire_774;
    wire new_Jinkela_wire_692;
    wire _0509_;
    wire new_Jinkela_wire_1529;
    wire new_Jinkela_wire_3080;
    wire new_Jinkela_wire_968;
    wire new_Jinkela_wire_345;
    wire new_Jinkela_wire_1997;
    wire new_Jinkela_wire_202;
    wire new_Jinkela_wire_1316;
    wire new_Jinkela_wire_1743;
    wire new_Jinkela_wire_2755;
    wire _0687_;
    wire new_Jinkela_wire_517;
    wire new_Jinkela_wire_1609;
    wire new_Jinkela_wire_1170;
    wire new_Jinkela_wire_2146;
    wire new_Jinkela_wire_616;
    wire new_Jinkela_wire_2520;
    wire new_Jinkela_wire_405;
    wire new_Jinkela_wire_915;
    wire new_Jinkela_wire_664;
    wire new_Jinkela_wire_1314;
    wire new_Jinkela_wire_746;
    wire _0434_;
    wire new_Jinkela_wire_2913;
    wire new_Jinkela_wire_1635;
    wire new_Jinkela_wire_2622;
    wire new_Jinkela_wire_2252;
    wire new_Jinkela_wire_2349;
    wire new_Jinkela_wire_913;
    wire _0231_;
    wire new_Jinkela_wire_132;
    wire new_Jinkela_wire_2599;
    wire new_Jinkela_wire_465;
    wire new_Jinkela_wire_359;
    wire new_Jinkela_wire_768;
    wire new_Jinkela_wire_2696;
    wire new_Jinkela_wire_2182;
    wire _0618_;
    wire _0376_;
    wire new_Jinkela_wire_3249;
    wire new_Jinkela_wire_3241;
    wire _0736_;
    wire new_Jinkela_wire_3252;
    wire new_Jinkela_wire_880;
    wire new_Jinkela_wire_1201;
    wire new_Jinkela_wire_690;
    wire new_Jinkela_wire_2461;
    wire new_Jinkela_wire_2944;
    wire new_Jinkela_wire_2806;
    wire new_Jinkela_wire_1231;
    wire new_Jinkela_wire_353;
    wire new_Jinkela_wire_2493;
    wire new_Jinkela_wire_1351;
    wire new_Jinkela_wire_2811;
    wire new_Jinkela_wire_123;
    wire new_Jinkela_wire_1993;
    wire _0324_;
    wire new_Jinkela_wire_3208;
    wire new_Jinkela_wire_1729;
    wire new_Jinkela_wire_757;
    wire new_Jinkela_wire_2407;
    wire new_Jinkela_wire_1472;
    wire new_Jinkela_wire_1944;
    wire new_Jinkela_wire_954;
    wire _0203_;
    wire new_Jinkela_wire_1406;
    wire new_Jinkela_wire_540;
    wire new_Jinkela_wire_2830;
    wire new_Jinkela_wire_1303;
    wire new_Jinkela_wire_592;
    wire new_Jinkela_wire_506;
    wire new_Jinkela_wire_666;
    wire new_Jinkela_wire_1239;
    wire new_Jinkela_wire_1335;
    wire new_Jinkela_wire_155;
    wire new_Jinkela_wire_2267;
    wire new_Jinkela_wire_2598;
    wire new_Jinkela_wire_2918;
    wire new_Jinkela_wire_242;
    wire _0493_;
    wire new_Jinkela_wire_500;
    wire new_Jinkela_wire_2875;
    wire new_Jinkela_wire_3062;
    wire new_Jinkela_wire_3085;
    wire _0179_;
    wire new_Jinkela_wire_1241;
    wire new_Jinkela_wire_942;
    wire new_Jinkela_wire_2394;
    wire new_Jinkela_wire_3155;
    wire new_Jinkela_wire_2721;
    wire new_Jinkela_wire_2679;
    wire new_Jinkela_wire_3138;
    wire new_Jinkela_wire_1893;
    wire new_Jinkela_wire_287;
    wire new_Jinkela_wire_935;
    wire _0148_;
    wire new_Jinkela_wire_1112;
    wire _0373_;
    wire new_Jinkela_wire_842;
    wire _0150_;
    wire new_Jinkela_wire_2286;
    wire new_Jinkela_wire_1221;
    wire new_Jinkela_wire_1131;
    wire new_Jinkela_wire_759;
    wire new_Jinkela_wire_1546;
    wire new_Jinkela_wire_2239;
    wire new_Jinkela_wire_1617;
    wire _0340_;
    wire _0343_;
    wire new_Jinkela_wire_3013;
    wire _0458_;
    wire new_Jinkela_wire_721;
    wire new_Jinkela_wire_3023;
    wire new_Jinkela_wire_1781;
    wire _0081_;
    wire new_Jinkela_wire_2754;
    wire _0746_;
    wire new_Jinkela_wire_2618;
    wire new_Jinkela_wire_1801;
    wire new_Jinkela_wire_1226;
    wire new_Jinkela_wire_3116;
    wire new_Jinkela_wire_1806;
    wire new_Jinkela_wire_2562;
    wire _0169_;
    wire _0450_;
    wire new_Jinkela_wire_2809;
    wire _0550_;
    wire new_Jinkela_wire_1508;
    wire new_net_4;
    wire new_Jinkela_wire_3269;
    wire new_Jinkela_wire_445;
    wire new_Jinkela_wire_1133;
    wire new_Jinkela_wire_1587;
    wire new_Jinkela_wire_2727;
    wire new_Jinkela_wire_321;
    wire new_Jinkela_wire_615;
    wire new_Jinkela_wire_948;
    wire _0315_;
    wire new_Jinkela_wire_1091;
    wire new_Jinkela_wire_105;
    wire new_Jinkela_wire_1115;
    wire new_Jinkela_wire_973;
    wire _0002_;
    wire new_Jinkela_wire_2192;
    wire new_Jinkela_wire_673;
    wire new_Jinkela_wire_3213;
    wire new_Jinkela_wire_1321;
    wire new_Jinkela_wire_2061;
    wire _0471_;
    wire new_Jinkela_wire_1306;
    wire new_Jinkela_wire_981;
    wire new_Jinkela_wire_1866;
    wire new_Jinkela_wire_1010;
    wire new_Jinkela_wire_1639;
    wire new_Jinkela_wire_2498;
    wire new_Jinkela_wire_651;
    wire new_Jinkela_wire_2655;
    wire new_Jinkela_wire_38;
    wire new_Jinkela_wire_554;
    wire new_Jinkela_wire_2092;
    wire new_Jinkela_wire_2770;
    wire new_Jinkela_wire_2315;
    wire new_Jinkela_wire_2961;
    wire new_Jinkela_wire_596;
    wire new_Jinkela_wire_1154;
    wire new_Jinkela_wire_3110;
    wire new_Jinkela_wire_789;
    wire new_Jinkela_wire_2982;
    wire new_Jinkela_wire_927;
    wire new_Jinkela_wire_1100;
    wire new_Jinkela_wire_2926;
    wire _0792_;
    wire new_Jinkela_wire_3124;
    wire new_Jinkela_wire_65;
    wire new_Jinkela_wire_3230;
    wire new_Jinkela_wire_1114;
    wire _0334_;
    wire new_Jinkela_wire_1300;
    wire new_Jinkela_wire_2699;
    wire _0516_;
    wire new_Jinkela_wire_189;
    wire new_Jinkela_wire_2786;
    wire new_Jinkela_wire_499;
    wire new_Jinkela_wire_1591;
    wire _0066_;
    wire new_Jinkela_wire_572;
    wire new_Jinkela_wire_282;
    wire new_Jinkela_wire_874;
    wire new_Jinkela_wire_3254;
    wire new_Jinkela_wire_1181;
    wire new_Jinkela_wire_1065;
    wire new_Jinkela_wire_1421;
    wire new_Jinkela_wire_2839;
    wire _0394_;
    wire new_Jinkela_wire_2843;
    wire new_Jinkela_wire_969;
    wire new_Jinkela_wire_817;
    wire new_Jinkela_wire_1408;
    wire new_Jinkela_wire_821;
    wire _0563_;
    wire new_Jinkela_wire_136;
    wire new_Jinkela_wire_271;
    wire _0261_;
    wire new_Jinkela_wire_2478;
    wire new_Jinkela_wire_1979;
    wire new_Jinkela_wire_1521;
    wire new_Jinkela_wire_1126;
    wire new_Jinkela_wire_1934;
    wire _0379_;
    wire new_Jinkela_wire_2097;
    wire new_Jinkela_wire_687;
    wire new_Jinkela_wire_492;
    wire new_Jinkela_wire_1438;
    wire new_Jinkela_wire_1725;
    wire new_Jinkela_wire_112;
    wire new_Jinkela_wire_1415;
    wire new_Jinkela_wire_2900;
    wire new_Jinkela_wire_2583;
    wire new_Jinkela_wire_83;
    wire new_Jinkela_wire_3317;
    wire new_Jinkela_wire_2709;
    wire new_Jinkela_wire_1034;
    wire _0640_;
    wire new_Jinkela_wire_1148;
    wire new_Jinkela_wire_1720;
    wire _0419_;
    wire new_Jinkela_wire_176;
    wire new_Jinkela_wire_497;
    wire new_Jinkela_wire_3276;
    wire _0602_;
    wire new_Jinkela_wire_3248;
    wire new_Jinkela_wire_929;
    wire new_Jinkela_wire_780;
    wire new_Jinkela_wire_2856;
    wire _0515_;
    wire new_Jinkela_wire_1594;
    wire new_Jinkela_wire_980;
    wire new_Jinkela_wire_2515;
    wire new_Jinkela_wire_1779;
    wire new_Jinkela_wire_3226;
    wire _0530_;
    wire _0375_;
    wire new_Jinkela_wire_1141;
    wire new_Jinkela_wire_2105;
    wire new_Jinkela_wire_1471;
    wire new_Jinkela_wire_1244;
    wire new_Jinkela_wire_3120;
    wire _0594_;
    wire new_Jinkela_wire_122;
    wire _0688_;
    wire _0035_;
    wire new_Jinkela_wire_952;
    wire new_Jinkela_wire_1840;
    wire new_Jinkela_wire_160;
    wire new_Jinkela_wire_2553;
    wire new_Jinkela_wire_971;
    wire new_Jinkela_wire_1289;
    wire _0577_;
    wire new_Jinkela_wire_1704;
    wire new_Jinkela_wire_3185;
    wire new_Jinkela_wire_1296;
    wire new_Jinkela_wire_3;
    wire new_Jinkela_wire_452;
    wire new_Jinkela_wire_1816;
    wire _0223_;
    wire new_net_1475;
    wire new_Jinkela_wire_761;
    wire new_Jinkela_wire_2998;
    wire new_Jinkela_wire_3227;
    wire new_Jinkela_wire_2509;
    wire new_Jinkela_wire_870;
    wire new_Jinkela_wire_1574;
    wire new_Jinkela_wire_2234;
    wire new_Jinkela_wire_1076;
    wire new_Jinkela_wire_2215;
    wire _0389_;
    wire new_Jinkela_wire_1689;
    wire new_Jinkela_wire_2392;
    wire new_Jinkela_wire_2403;
    wire _0720_;
    wire new_Jinkela_wire_1347;
    wire new_Jinkela_wire_1093;
    wire new_Jinkela_wire_2528;
    wire new_Jinkela_wire_3053;
    wire new_Jinkela_wire_2938;
    wire new_Jinkela_wire_1717;
    wire new_Jinkela_wire_26;
    wire new_Jinkela_wire_3119;
    wire new_Jinkela_wire_3096;
    wire _0076_;
    wire _0366_;
    wire new_Jinkela_wire_2757;
    wire new_Jinkela_wire_1449;
    wire new_Jinkela_wire_2282;
    wire _0793_;
    wire new_Jinkela_wire_3285;
    wire new_Jinkela_wire_3133;
    wire new_Jinkela_wire_1683;
    wire _0336_;
    wire new_Jinkela_wire_505;
    wire new_Jinkela_wire_1843;
    wire new_Jinkela_wire_612;
    wire _0435_;
    wire new_Jinkela_wire_1459;
    wire new_Jinkela_wire_962;
    wire new_Jinkela_wire_2006;
    wire new_Jinkela_wire_3264;
    wire new_Jinkela_wire_595;
    wire new_Jinkela_wire_1501;
    wire new_Jinkela_wire_1786;
    wire new_net_5;
    wire _0250_;
    wire new_Jinkela_wire_2098;
    wire new_Jinkela_wire_2380;
    wire new_Jinkela_wire_2656;
    wire new_net_1471;
    wire new_Jinkela_wire_1409;
    wire new_Jinkela_wire_1660;
    wire new_Jinkela_wire_2406;
    wire new_Jinkela_wire_2993;
    wire _0499_;
    wire new_Jinkela_wire_3130;
    wire _0024_;
    wire new_Jinkela_wire_1251;
    wire _0454_;
    wire new_Jinkela_wire_1343;
    wire new_Jinkela_wire_1085;
    wire new_Jinkela_wire_3191;
    wire _0528_;
    wire new_Jinkela_wire_1543;
    wire new_Jinkela_wire_1593;
    wire new_Jinkela_wire_356;
    wire new_Jinkela_wire_2866;
    wire new_Jinkela_wire_2857;
    wire new_Jinkela_wire_472;
    wire new_Jinkela_wire_802;
    wire new_Jinkela_wire_3333;
    wire _0348_;
    wire _0455_;
    wire _0303_;
    wire _0649_;
    wire _0008_;
    wire new_Jinkela_wire_2336;
    wire _0091_;
    wire new_Jinkela_wire_2554;
    wire _0307_;
    wire new_Jinkela_wire_296;
    wire new_Jinkela_wire_2080;
    wire _0258_;
    wire new_Jinkela_wire_1907;
    wire new_Jinkela_wire_2016;
    wire _0588_;
    wire _0404_;
    wire new_Jinkela_wire_3223;
    wire new_Jinkela_wire_2157;
    wire new_Jinkela_wire_756;
    wire new_Jinkela_wire_1865;
    wire _0639_;
    wire _0463_;
    wire new_Jinkela_wire_2800;
    wire new_Jinkela_wire_1784;
    wire new_Jinkela_wire_909;
    wire _0418_;
    wire new_Jinkela_wire_3043;
    wire new_Jinkela_wire_2265;
    wire new_Jinkela_wire_2128;
    wire new_Jinkela_wire_2957;
    wire new_Jinkela_wire_1040;
    wire new_Jinkela_wire_2022;
    wire new_Jinkela_wire_1137;
    wire new_Jinkela_wire_127;
    wire new_Jinkela_wire_1404;
    wire _0170_;
    wire new_Jinkela_wire_2849;
    wire new_Jinkela_wire_3244;
    wire new_Jinkela_wire_1269;
    wire new_Jinkela_wire_113;
    wire new_Jinkela_wire_2263;
    wire _0056_;
    wire new_Jinkela_wire_694;
    wire new_Jinkela_wire_2854;
    wire new_Jinkela_wire_1579;
    wire _0440_;
    wire new_Jinkela_wire_856;
    wire new_Jinkela_wire_3005;
    wire _0082_;
    wire new_Jinkela_wire_78;
    wire new_Jinkela_wire_2266;
    wire new_Jinkela_wire_1904;
    wire new_Jinkela_wire_267;
    wire new_Jinkela_wire_801;
    wire new_Jinkela_wire_752;
    wire _0322_;
    wire new_Jinkela_wire_634;
    wire new_Jinkela_wire_2573;
    wire new_Jinkela_wire_82;
    wire _0182_;
    wire new_Jinkela_wire_2200;
    wire _0123_;
    wire new_Jinkela_wire_600;
    wire new_Jinkela_wire_2953;
    wire new_Jinkela_wire_349;
    wire new_Jinkela_wire_857;
    wire new_Jinkela_wire_1484;
    wire new_Jinkela_wire_1410;
    wire new_Jinkela_wire_2967;
    wire _0476_;
    wire new_Jinkela_wire_1834;
    wire new_Jinkela_wire_556;
    wire _0489_;
    wire new_Jinkela_wire_3198;
    wire new_Jinkela_wire_1629;
    wire new_Jinkela_wire_2694;
    wire new_Jinkela_wire_3092;
    wire new_Jinkela_wire_1411;
    wire new_Jinkela_wire_313;
    wire _0761_;
    wire _0143_;
    wire new_Jinkela_wire_1402;
    wire new_Jinkela_wire_1422;
    wire new_Jinkela_wire_2817;
    wire new_Jinkela_wire_8;
    wire new_net_1469;
    wire new_Jinkela_wire_1876;
    wire new_Jinkela_wire_2681;
    wire new_Jinkela_wire_2923;
    wire new_Jinkela_wire_1745;
    wire _0175_;
    wire _0054_;
    wire new_Jinkela_wire_797;
    wire new_Jinkela_wire_2269;
    wire new_Jinkela_wire_3279;
    wire _0723_;
    wire new_Jinkela_wire_665;
    wire new_Jinkela_wire_1905;
    wire new_Jinkela_wire_1036;
    wire new_Jinkela_wire_2305;
    wire _0553_;
    wire _0729_;
    wire new_Jinkela_wire_1685;
    wire new_Jinkela_wire_834;
    wire _0279_;
    wire new_Jinkela_wire_1118;
    wire new_Jinkela_wire_361;
    wire new_Jinkela_wire_1642;
    wire new_Jinkela_wire_795;
    wire _0116_;
    wire new_Jinkela_wire_710;
    wire new_Jinkela_wire_740;
    wire new_Jinkela_wire_1158;
    wire _0355_;
    wire new_Jinkela_wire_800;
    wire new_Jinkela_wire_2525;
    wire new_Jinkela_wire_1915;
    wire new_Jinkela_wire_3057;
    wire new_Jinkela_wire_3240;
    wire _0433_;
    wire new_Jinkela_wire_2707;
    wire new_Jinkela_wire_2255;
    wire _0690_;
    wire new_Jinkela_wire_1883;
    wire _0487_;
    wire new_Jinkela_wire_1081;
    wire new_Jinkela_wire_2572;
    wire new_Jinkela_wire_1795;
    wire new_Jinkela_wire_995;
    wire _0513_;
    wire new_Jinkela_wire_2858;
    wire new_Jinkela_wire_102;
    wire new_Jinkela_wire_63;
    wire new_Jinkela_wire_3175;
    wire _0027_;
    wire new_Jinkela_wire_1761;
    wire new_Jinkela_wire_1049;
    wire new_Jinkela_wire_1649;
    wire new_Jinkela_wire_329;
    wire new_Jinkela_wire_149;
    wire new_Jinkela_wire_3194;
    wire new_Jinkela_wire_2904;
    wire new_Jinkela_wire_3268;
    wire new_Jinkela_wire_3072;
    wire new_Jinkela_wire_333;
    wire new_Jinkela_wire_33;
    wire new_Jinkela_wire_2323;
    wire new_Jinkela_wire_467;
    wire new_Jinkela_wire_429;
    wire _0566_;
    wire new_Jinkela_wire_2352;
    wire new_Jinkela_wire_3049;
    wire new_Jinkela_wire_703;
    wire new_Jinkela_wire_1968;
    wire new_Jinkela_wire_1029;
    wire new_Jinkela_wire_2749;
    wire new_Jinkela_wire_1267;
    wire new_Jinkela_wire_1805;
    wire new_Jinkela_wire_3334;
    wire new_Jinkela_wire_1514;
    wire _0393_;
    wire new_Jinkela_wire_3166;
    wire new_Jinkela_wire_413;
    wire new_Jinkela_wire_1265;
    wire new_Jinkela_wire_1523;
    wire new_Jinkela_wire_3189;
    wire new_Jinkela_wire_1760;
    wire new_Jinkela_wire_940;
    wire new_Jinkela_wire_2505;
    wire new_Jinkela_wire_299;
    wire new_Jinkela_wire_1016;
    wire new_Jinkela_wire_663;
    wire new_Jinkela_wire_1808;
    wire new_Jinkela_wire_206;
    wire new_Jinkela_wire_2595;
    wire new_Jinkela_wire_993;
    wire new_Jinkela_wire_2134;
    wire new_Jinkela_wire_1044;
    wire new_Jinkela_wire_2387;
    wire new_Jinkela_wire_2430;
    wire new_Jinkela_wire_755;
    wire _0025_;
    wire _0259_;
    wire _0788_;
    wire new_Jinkela_wire_963;
    wire _0665_;
    wire new_Jinkela_wire_2457;
    wire new_Jinkela_wire_2838;
    wire new_Jinkela_wire_579;
    wire new_Jinkela_wire_2504;
    wire new_Jinkela_wire_2735;
    wire _0492_;
    wire new_Jinkela_wire_2439;
    wire new_Jinkela_wire_1334;
    wire new_Jinkela_wire_207;
    wire new_Jinkela_wire_1610;
    wire new_Jinkela_wire_1911;
    wire _0053_;
    wire new_Jinkela_wire_1218;
    wire new_Jinkela_wire_625;
    wire new_Jinkela_wire_2832;
    wire new_Jinkela_wire_528;
    wire new_Jinkela_wire_2018;
    wire new_Jinkela_wire_1064;
    wire new_Jinkela_wire_2037;
    wire new_Jinkela_wire_3263;
    wire new_Jinkela_wire_2424;
    wire new_Jinkela_wire_1748;
    wire new_Jinkela_wire_51;
    wire new_Jinkela_wire_852;
    wire new_Jinkela_wire_1405;
    wire _0221_;
    wire _0230_;
    wire new_Jinkela_wire_1005;
    wire new_net_8;
    wire new_Jinkela_wire_1427;
    wire new_Jinkela_wire_1858;
    wire new_Jinkela_wire_2988;
    wire new_Jinkela_wire_487;
    wire new_Jinkela_wire_1960;
    wire _0308_;
    wire new_Jinkela_wire_2890;
    wire new_Jinkela_wire_1899;
    wire new_Jinkela_wire_2250;
    wire new_Jinkela_wire_2359;
    wire _0445_;
    wire new_Jinkela_wire_221;
    wire _0593_;
    wire _0712_;
    wire new_Jinkela_wire_892;
    wire _0104_;
    wire new_Jinkela_wire_1380;
    wire new_Jinkela_wire_291;
    wire new_Jinkela_wire_590;
    wire new_Jinkela_wire_330;
    wire new_Jinkela_wire_2219;
    wire new_Jinkela_wire_2968;
    wire new_Jinkela_wire_829;
    wire new_Jinkela_wire_1882;
    wire _0750_;
    wire _0748_;
    wire new_Jinkela_wire_166;
    wire new_Jinkela_wire_2863;
    wire new_Jinkela_wire_3300;
    wire new_Jinkela_wire_3102;
    wire _0291_;
    wire new_Jinkela_wire_1585;
    wire new_Jinkela_wire_238;
    wire new_Jinkela_wire_252;
    wire new_Jinkela_wire_2824;
    wire new_Jinkela_wire_283;
    wire new_Jinkela_wire_1302;
    wire new_Jinkela_wire_2208;
    wire _0542_;
    wire _0775_;
    wire new_Jinkela_wire_2444;
    wire new_Jinkela_wire_947;
    wire _0243_;
    wire new_Jinkela_wire_382;
    wire _0297_;
    wire _0673_;
    wire _0484_;
    wire new_Jinkela_wire_2425;
    wire new_Jinkela_wire_1463;
    wire new_Jinkela_wire_1462;
    wire new_Jinkela_wire_2578;
    wire new_Jinkela_wire_1022;
    wire new_Jinkela_wire_1487;
    wire new_Jinkela_wire_1027;
    wire new_Jinkela_wire_3061;
    wire new_Jinkela_wire_3159;
    wire new_Jinkela_wire_3064;
    wire new_Jinkela_wire_1823;
    wire new_Jinkela_wire_516;
    wire _0424_;
    wire _0478_;
    wire new_Jinkela_wire_3088;
    wire new_Jinkela_wire_1;
    wire new_Jinkela_wire_2069;
    wire new_Jinkela_wire_812;
    wire new_Jinkela_wire_3233;
    wire new_Jinkela_wire_1560;
    wire new_Jinkela_wire_1096;
    wire new_Jinkela_wire_2288;
    wire new_Jinkela_wire_1656;
    wire _0780_;
    wire new_Jinkela_wire_2943;
    wire _0488_;
    wire new_Jinkela_wire_2196;
    wire _0145_;
    wire new_Jinkela_wire_2161;
    wire new_Jinkela_wire_15;
    wire new_Jinkela_wire_2766;
    wire _0080_;
    wire new_Jinkela_wire_2375;
    wire new_Jinkela_wire_2796;
    wire new_Jinkela_wire_1222;
    wire new_Jinkela_wire_2021;
    wire new_Jinkela_wire_2070;
    wire new_Jinkela_wire_1663;
    wire new_Jinkela_wire_1138;
    wire _0335_;
    wire new_Jinkela_wire_914;
    wire _0141_;
    wire new_Jinkela_wire_1278;
    wire new_Jinkela_wire_1288;
    wire new_Jinkela_wire_254;
    wire new_Jinkela_wire_2268;
    wire new_Jinkela_wire_1588;
    wire new_Jinkela_wire_3315;
    wire _0329_;
    wire new_Jinkela_wire_2604;
    wire new_Jinkela_wire_3332;
    wire new_Jinkela_wire_376;
    wire new_Jinkela_wire_2912;
    wire new_Jinkela_wire_1108;
    wire new_Jinkela_wire_153;
    wire new_Jinkela_wire_190;
    wire new_Jinkela_wire_869;
    wire new_Jinkela_wire_945;
    wire new_Jinkela_wire_2121;
    wire new_Jinkela_wire_2777;
    wire new_Jinkela_wire_2010;
    wire new_Jinkela_wire_3218;
    wire new_Jinkela_wire_2726;
    wire new_Jinkela_wire_2725;
    wire new_Jinkela_wire_2253;
    wire new_Jinkela_wire_391;
    wire new_Jinkela_wire_1026;
    wire _0397_;
    wire new_Jinkela_wire_1558;
    wire new_Jinkela_wire_1971;
    wire new_Jinkela_wire_893;
    wire new_Jinkela_wire_678;
    wire new_Jinkela_wire_805;
    wire new_Jinkela_wire_1750;
    wire _0728_;
    wire new_Jinkela_wire_3107;
    wire new_Jinkela_wire_342;
    wire _0115_;
    wire new_Jinkela_wire_1978;
    wire new_Jinkela_wire_2657;
    wire new_Jinkela_wire_1564;
    wire new_Jinkela_wire_1671;
    wire _0139_;
    wire new_Jinkela_wire_3007;
    wire new_Jinkela_wire_548;
    wire new_Jinkela_wire_1167;
    wire new_Jinkela_wire_2997;
    wire new_Jinkela_wire_1213;
    wire new_Jinkela_wire_1465;
    wire new_Jinkela_wire_1936;
    wire new_Jinkela_wire_1803;
    wire _0128_;
    wire new_Jinkela_wire_165;
    wire _0641_;
    wire new_Jinkela_wire_394;
    wire new_Jinkela_wire_1124;
    wire new_Jinkela_wire_1598;
    wire new_Jinkela_wire_2274;
    wire new_Jinkela_wire_1679;
    wire new_Jinkela_wire_2496;
    wire _0254_;
    wire new_Jinkela_wire_2283;
    wire new_Jinkela_wire_2028;
    wire new_Jinkela_wire_2591;
    wire new_Jinkela_wire_3076;
    wire _0726_;
    wire new_Jinkela_wire_1810;
    wire new_Jinkela_wire_1140;
    wire new_Jinkela_wire_209;
    wire new_Jinkela_wire_1700;
    wire new_Jinkela_wire_2143;
    wire new_Jinkela_wire_2126;
    wire new_Jinkela_wire_2199;
    wire new_Jinkela_wire_439;
    wire new_Jinkela_wire_2883;
    wire new_Jinkela_wire_384;
    wire new_Jinkela_wire_731;
    wire new_Jinkela_wire_626;
    wire _0135_;
    wire new_Jinkela_wire_507;
    wire _0702_;
    wire new_Jinkela_wire_715;
    wire _0338_;
    wire new_Jinkela_wire_511;
    wire new_Jinkela_wire_1200;
    wire new_Jinkela_wire_2541;
    wire new_Jinkela_wire_1986;
    wire new_Jinkela_wire_779;
    wire new_Jinkela_wire_1855;
    wire new_Jinkela_wire_3324;
    wire new_Jinkela_wire_1256;
    wire new_Jinkela_wire_1874;
    wire new_Jinkela_wire_2499;
    wire new_Jinkela_wire_1369;
    wire new_net_2;
    wire _0090_;
    wire new_Jinkela_wire_2065;
    wire new_Jinkela_wire_2129;
    wire new_Jinkela_wire_1247;
    wire new_Jinkela_wire_685;
    wire new_Jinkela_wire_2501;
    wire new_Jinkela_wire_1782;
    wire new_Jinkela_wire_3173;
    wire new_Jinkela_wire_808;
    wire new_Jinkela_wire_424;
    wire new_Jinkela_wire_217;
    wire new_Jinkela_wire_498;
    wire new_net_1479;
    wire new_Jinkela_wire_2059;
    wire new_Jinkela_wire_2663;
    wire new_Jinkela_wire_2361;
    wire _0532_;
    wire _0180_;
    wire _0597_;
    wire new_Jinkela_wire_985;
    wire _0365_;
    wire new_Jinkela_wire_748;
    wire new_Jinkela_wire_648;
    wire _0414_;
    wire _0658_;
    wire new_Jinkela_wire_225;
    wire new_Jinkela_wire_1413;
    wire new_Jinkela_wire_1967;
    wire _0251_;
    wire new_Jinkela_wire_3210;
    wire _0796_;
    wire new_Jinkela_wire_1130;
    wire new_Jinkela_wire_393;
    wire new_Jinkela_wire_2204;
    wire _0560_;
    wire new_Jinkela_wire_587;
    wire _0791_;
    wire new_Jinkela_wire_1681;
    wire new_Jinkela_wire_1771;
    wire _0386_;
    wire new_Jinkela_wire_873;
    wire new_Jinkela_wire_864;
    wire new_Jinkela_wire_2643;
    wire new_Jinkela_wire_1632;
    wire new_Jinkela_wire_2429;
    wire new_Jinkela_wire_2419;
    wire _0272_;
    wire new_Jinkela_wire_109;
    wire new_Jinkela_wire_1032;
    wire new_Jinkela_wire_2958;
    wire new_Jinkela_wire_682;
    wire new_Jinkela_wire_953;
    wire new_Jinkela_wire_1930;
    wire new_Jinkela_wire_2180;
    wire new_Jinkela_wire_152;
    wire _0576_;
    wire new_Jinkela_wire_1358;
    wire _0697_;
    wire new_Jinkela_wire_599;
    wire new_Jinkela_wire_1709;
    wire _0426_;
    wire _0287_;
    wire new_Jinkela_wire_1686;
    wire _0352_;
    wire new_Jinkela_wire_421;
    wire new_Jinkela_wire_3111;
    wire new_Jinkela_wire_2045;
    wire _0196_;
    wire new_Jinkela_wire_187;
    wire new_Jinkela_wire_444;
    wire _0698_;
    wire new_Jinkela_wire_1260;
    wire _0022_;
    wire _0591_;
    wire new_Jinkela_wire_1510;
    wire new_Jinkela_wire_2925;
    wire new_Jinkela_wire_175;
    wire _0667_;
    wire new_Jinkela_wire_2920;
    wire new_Jinkela_wire_831;
    wire new_Jinkela_wire_201;
    wire new_Jinkela_wire_2503;
    wire _0369_;
    wire new_Jinkela_wire_1476;
    wire new_Jinkela_wire_383;
    wire new_Jinkela_wire_1279;
    wire new_Jinkela_wire_526;
    wire _0766_;
    wire new_Jinkela_wire_2005;
    wire _0425_;
    wire new_Jinkela_wire_2030;
    wire new_Jinkela_wire_2303;
    wire new_Jinkela_wire_369;
    wire new_Jinkela_wire_921;
    wire new_Jinkela_wire_2035;
    wire new_Jinkela_wire_1258;
    wire new_Jinkela_wire_1918;
    wire new_Jinkela_wire_637;
    wire _0164_;
    wire new_Jinkela_wire_303;
    wire new_Jinkela_wire_1573;
    wire _0589_;
    wire new_Jinkela_wire_1123;
    wire new_Jinkela_wire_2103;
    wire new_Jinkela_wire_1103;
    wire _0579_;
    wire _0086_;
    wire new_Jinkela_wire_1173;
    wire new_Jinkela_wire_2110;
    wire new_Jinkela_wire_3292;
    wire new_Jinkela_wire_1917;
    wire new_Jinkela_wire_2774;
    wire new_Jinkela_wire_1908;
    wire new_Jinkela_wire_2847;
    wire _0783_;
    wire new_Jinkela_wire_557;
    wire new_Jinkela_wire_2293;
    wire _0453_;
    wire new_Jinkela_wire_1903;
    wire new_Jinkela_wire_1931;
    wire new_Jinkela_wire_52;
    wire new_Jinkela_wire_567;
    wire new_Jinkela_wire_3243;
    wire new_Jinkela_wire_1102;
    wire new_Jinkela_wire_1822;
    wire new_Jinkela_wire_111;
    wire _0739_;
    wire new_Jinkela_wire_1156;
    wire new_Jinkela_wire_2759;
    wire new_Jinkela_wire_2797;
    wire new_Jinkela_wire_2187;
    wire _0074_;
    wire new_Jinkela_wire_3137;
    wire _0097_;
    wire new_Jinkela_wire_3029;
    wire new_Jinkela_wire_1790;
    wire new_Jinkela_wire_1845;
    wire new_Jinkela_wire_1753;
    wire _0781_;
    wire _0447_;
    wire new_Jinkela_wire_3316;
    wire new_Jinkela_wire_475;
    wire new_Jinkela_wire_3182;
    wire new_Jinkela_wire_43;
    wire _0248_;
    wire new_Jinkela_wire_1756;
    wire new_Jinkela_wire_3322;
    wire new_Jinkela_wire_607;
    wire new_Jinkela_wire_2413;
    wire new_Jinkela_wire_1541;
    wire new_Jinkela_wire_1581;
    wire new_Jinkela_wire_3245;
    wire new_Jinkela_wire_883;
    wire new_Jinkela_wire_3256;
    wire new_Jinkela_wire_890;
    wire new_Jinkela_wire_2911;
    wire new_Jinkela_wire_3304;
    wire new_Jinkela_wire_311;
    wire new_Jinkela_wire_426;
    wire new_Jinkela_wire_1469;
    wire new_Jinkela_wire_598;
    wire new_Jinkela_wire_1516;
    wire _0555_;
    wire new_Jinkela_wire_2820;
    wire new_Jinkela_wire_2058;
    wire _0204_;
    wire new_Jinkela_wire_3038;
    wire new_Jinkela_wire_2737;
    wire new_Jinkela_wire_411;
    wire new_Jinkela_wire_42;
    wire new_Jinkela_wire_889;
    wire new_Jinkela_wire_328;
    wire new_Jinkela_wire_2718;
    wire new_Jinkela_wire_106;
    wire new_Jinkela_wire_3054;
    wire _0134_;
    wire new_Jinkela_wire_2047;
    wire new_Jinkela_wire_1457;
    wire new_Jinkela_wire_2876;
    wire _0548_;
    wire new_Jinkela_wire_1171;
    wire new_Jinkela_wire_638;
    wire _0101_;
    wire new_Jinkela_wire_2042;
    wire new_Jinkela_wire_2744;
    wire new_Jinkela_wire_10;
    wire new_Jinkela_wire_3164;
    wire _0713_;
    wire new_Jinkela_wire_22;
    wire new_Jinkela_wire_146;
    wire new_Jinkela_wire_1392;
    wire _0722_;
    wire new_Jinkela_wire_1388;
    wire new_Jinkela_wire_1940;
    wire new_Jinkela_wire_2822;
    wire new_Jinkela_wire_244;
    wire new_Jinkela_wire_1500;
    wire new_Jinkela_wire_1070;
    wire _0765_;
    wire new_Jinkela_wire_2174;
    wire _0494_;
    wire new_Jinkela_wire_2277;
    wire new_Jinkela_wire_2814;
    wire new_Jinkela_wire_532;
    wire new_Jinkela_wire_3089;
    wire new_Jinkela_wire_2706;
    wire new_Jinkela_wire_1434;
    wire _0505_;
    wire new_Jinkela_wire_75;
    wire new_Jinkela_wire_1283;
    wire new_Jinkela_wire_1028;
    wire new_Jinkela_wire_991;
    wire new_Jinkela_wire_1243;
    wire new_Jinkela_wire_297;
    wire new_Jinkela_wire_144;
    wire new_Jinkela_wire_3081;
    wire new_Jinkela_wire_1164;
    wire new_Jinkela_wire_198;
    wire new_Jinkela_wire_2996;
    wire _0387_;
    wire new_Jinkela_wire_1826;
    wire new_Jinkela_wire_3037;
    wire new_Jinkela_wire_262;
    wire new_Jinkela_wire_392;
    wire _0514_;
    wire new_Jinkela_wire_3311;
    wire new_Jinkela_wire_794;
    wire new_Jinkela_wire_28;
    wire _0683_;
    wire new_Jinkela_wire_2483;
    wire new_Jinkela_wire_1162;
    wire new_Jinkela_wire_3028;
    wire new_Jinkela_wire_1537;
    wire new_Jinkela_wire_1875;
    wire new_Jinkela_wire_1852;
    wire _0085_;
    wire new_Jinkela_wire_580;
    wire new_Jinkela_wire_2074;
    wire new_Jinkela_wire_219;
    wire new_Jinkela_wire_1824;
    wire new_Jinkela_wire_688;
    wire new_Jinkela_wire_3216;
    wire new_Jinkela_wire_2975;
    wire new_Jinkela_wire_1177;
    wire new_Jinkela_wire_1207;
    wire new_Jinkela_wire_1690;
    wire new_Jinkela_wire_1921;
    wire new_Jinkela_wire_2966;
    wire _0423_;
    wire new_Jinkela_wire_2738;
    wire new_Jinkela_wire_1497;
    wire _0313_;
    wire _0382_;
    wire new_Jinkela_wire_11;
    wire new_Jinkela_wire_825;
    wire new_Jinkela_wire_473;
    wire new_Jinkela_wire_305;
    wire new_Jinkela_wire_233;
    wire _0636_;
    wire new_Jinkela_wire_2678;
    wire _0790_;
    wire new_Jinkela_wire_3099;
    wire _0669_;
    wire _0202_;
    wire new_Jinkela_wire_1295;
    wire new_Jinkela_wire_919;
    wire new_Jinkela_wire_2455;
    wire new_Jinkela_wire_552;
    wire new_Jinkela_wire_2083;
    wire new_Jinkela_wire_1445;
    wire _0719_;
    wire new_Jinkela_wire_1095;
    wire new_Jinkela_wire_2431;
    wire new_Jinkela_wire_1793;
    wire new_Jinkela_wire_2459;
    wire new_Jinkela_wire_904;
    wire new_Jinkela_wire_3075;
    wire new_Jinkela_wire_2816;
    wire _0306_;
    wire new_Jinkela_wire_88;
    wire new_Jinkela_wire_1152;
    wire new_Jinkela_wire_265;
    wire new_Jinkela_wire_2363;
    wire new_Jinkela_wire_667;
    wire new_Jinkela_wire_1425;
    wire new_Jinkela_wire_1412;
    wire new_Jinkela_wire_2928;
    wire new_Jinkela_wire_494;
    wire new_Jinkela_wire_714;
    wire new_Jinkela_wire_813;
    wire new_Jinkela_wire_2008;
    wire new_Jinkela_wire_485;
    wire new_Jinkela_wire_578;
    wire new_Jinkela_wire_1902;
    wire new_Jinkela_wire_3278;
    wire new_Jinkela_wire_3288;
    wire new_Jinkela_wire_2954;
    wire new_Jinkela_wire_374;
    wire new_Jinkela_wire_2730;
    wire new_net_1465;
    wire _0218_;
    wire _0094_;
    wire new_Jinkela_wire_3293;
    wire new_Jinkela_wire_3221;
    wire new_Jinkela_wire_2147;
    wire new_Jinkela_wire_294;
    wire new_Jinkela_wire_1767;
    wire new_Jinkela_wire_1833;
    wire _0410_;
    wire new_Jinkela_wire_412;
    wire new_Jinkela_wire_704;
    wire new_Jinkela_wire_639;
    wire new_Jinkela_wire_1495;
    wire new_Jinkela_wire_143;
    wire new_Jinkela_wire_1371;
    wire _0486_;
    wire _0467_;
    wire new_Jinkela_wire_1737;
    wire new_Jinkela_wire_1636;
    wire new_Jinkela_wire_2421;
    wire new_Jinkela_wire_2463;
    wire new_Jinkela_wire_543;
    wire _0738_;
    wire new_Jinkela_wire_1976;
    wire new_Jinkela_wire_770;
    wire _0163_;
    wire new_Jinkela_wire_1382;
    wire new_Jinkela_wire_1250;
    wire new_Jinkela_wire_979;
    wire _0626_;
    wire new_Jinkela_wire_1011;
    wire new_Jinkela_wire_2690;
    wire new_Jinkela_wire_1864;
    wire new_Jinkela_wire_1385;
    wire _0270_;
    wire new_Jinkela_wire_1906;
    wire new_Jinkela_wire_1929;
    wire new_Jinkela_wire_2764;
    wire new_Jinkela_wire_164;
    wire new_Jinkela_wire_837;
    wire new_Jinkela_wire_1966;
    wire new_Jinkela_wire_2781;
    wire new_Jinkela_wire_840;
    wire new_Jinkela_wire_2104;
    wire new_Jinkela_wire_3253;
    wire _0144_;
    wire new_Jinkela_wire_1326;
    wire new_Jinkela_wire_1691;
    wire _0265_;
    wire new_Jinkela_wire_2418;
    wire new_Jinkela_wire_2485;
    wire _0774_;
    wire new_Jinkela_wire_2536;
    wire new_Jinkela_wire_367;
    wire new_Jinkela_wire_196;
    wire new_Jinkela_wire_2308;
    wire new_Jinkela_wire_2871;
    wire new_Jinkela_wire_1055;
    wire _0485_;
    wire new_Jinkela_wire_3204;
    wire new_Jinkela_wire_2049;
    wire new_Jinkela_wire_2319;
    wire new_Jinkela_wire_183;
    wire new_Jinkela_wire_2535;
    wire _0028_;
    wire new_Jinkela_wire_960;
    wire new_Jinkela_wire_292;
    wire new_Jinkela_wire_3048;
    wire new_Jinkela_wire_324;
    wire new_Jinkela_wire_2549;
    wire new_Jinkela_wire_3044;
    wire new_Jinkela_wire_195;
    wire new_Jinkela_wire_2597;
    wire new_Jinkela_wire_27;
    wire new_Jinkela_wire_3183;
    wire new_Jinkela_wire_430;
    wire _0498_;
    wire new_Jinkela_wire_849;
    wire _0015_;
    wire new_Jinkela_wire_3035;
    wire new_Jinkela_wire_2329;
    wire new_Jinkela_wire_2891;
    wire new_net_1;
    wire _0318_;
    wire new_Jinkela_wire_2558;
    wire new_Jinkela_wire_490;
    wire new_Jinkela_wire_2819;
    wire new_Jinkela_wire_3103;
    wire new_Jinkela_wire_2484;
    wire new_Jinkela_wire_1489;
    wire new_Jinkela_wire_2815;
    wire new_Jinkela_wire_327;
    wire new_Jinkela_wire_2950;
    wire new_Jinkela_wire_2649;
    wire new_Jinkela_wire_1048;
    wire new_Jinkela_wire_1539;
    wire new_Jinkela_wire_1312;
    wire new_Jinkela_wire_1249;
    wire _0157_;
    wire new_Jinkela_wire_1804;
    wire new_Jinkela_wire_1015;
    wire new_Jinkela_wire_450;
    wire new_Jinkela_wire_150;
    wire _0103_;
    wire new_Jinkela_wire_2170;
    wire new_Jinkela_wire_484;
    wire new_Jinkela_wire_434;
    wire new_Jinkela_wire_859;
    wire _0320_;
    wire _0519_;
    wire new_Jinkela_wire_159;
    wire new_Jinkela_wire_1542;
    wire new_Jinkela_wire_3121;
    wire new_Jinkela_wire_828;
    wire new_Jinkela_wire_2834;
    wire _0596_;
    wire new_Jinkela_wire_1999;
    wire new_Jinkela_wire_3074;
    wire _0432_;
    wire new_Jinkela_wire_990;
    wire new_Jinkela_wire_1675;
    wire _0117_;
    wire new_Jinkela_wire_531;
    wire new_Jinkela_wire_3093;
    wire new_Jinkela_wire_1013;
    wire new_Jinkela_wire_2412;
    wire new_Jinkela_wire_957;
    wire new_Jinkela_wire_1436;
    wire _0310_;
    wire new_Jinkela_wire_3314;
    wire _0545_;
    wire new_Jinkela_wire_2233;
    wire new_Jinkela_wire_2298;
    wire new_Jinkela_wire_13;
    wire _0567_;
    wire new_Jinkela_wire_1616;
    wire new_Jinkela_wire_1365;
    wire new_Jinkela_wire_1870;
    wire _0319_;
    wire new_Jinkela_wire_1046;
    wire _0078_;
    wire _0562_;
    wire new_Jinkela_wire_854;
    wire new_Jinkela_wire_2340;
    wire new_Jinkela_wire_449;
    wire new_Jinkela_wire_737;
    wire new_Jinkela_wire_1868;
    wire new_Jinkela_wire_400;
    wire new_Jinkela_wire_273;
    wire new_Jinkela_wire_446;
    wire new_Jinkela_wire_1766;
    wire new_Jinkela_wire_976;
    wire new_Jinkela_wire_899;
    wire new_Jinkela_wire_3203;
    wire new_Jinkela_wire_777;
    wire new_Jinkela_wire_2072;
    wire _0068_;
    wire new_Jinkela_wire_2898;
    wire new_Jinkela_wire_3050;
    wire _0311_;
    wire _0385_;
    wire _0628_;
    wire new_Jinkela_wire_1437;
    wire new_Jinkela_wire_3214;
    wire _0102_;
    wire new_Jinkela_wire_778;
    wire new_Jinkela_wire_2272;
    wire new_Jinkela_wire_1757;
    wire _0724_;
    wire _0633_;
    wire _0000_;
    wire new_Jinkela_wire_684;
    wire new_Jinkela_wire_1324;
    wire _0737_;
    wire new_Jinkela_wire_584;
    wire _0651_;
    wire new_Jinkela_wire_85;
    wire new_Jinkela_wire_1301;
    wire _0325_;
    wire new_Jinkela_wire_2919;
    wire new_Jinkela_wire_562;
    wire new_Jinkela_wire_2241;
    wire new_Jinkela_wire_147;
    wire _0511_;
    wire new_Jinkela_wire_2805;
    wire _0185_;
    wire new_Jinkela_wire_1920;
    wire new_Jinkela_wire_2784;
    wire new_Jinkela_wire_916;
    wire new_Jinkela_wire_2099;
    wire new_Jinkela_wire_1396;
    wire new_Jinkela_wire_3087;
    wire new_Jinkela_wire_2154;
    wire _0160_;
    wire new_Jinkela_wire_2639;
    wire new_Jinkela_wire_2309;
    wire new_Jinkela_wire_2335;
    wire _0742_;
    wire new_Jinkela_wire_1117;
    wire _0047_;
    wire new_Jinkela_wire_2003;
    wire new_Jinkela_wire_564;
    wire new_Jinkela_wire_1963;
    wire new_Jinkela_wire_2723;
    wire new_Jinkela_wire_1255;
    wire new_Jinkela_wire_1467;
    wire _0132_;
    wire _0295_;
    wire new_Jinkela_wire_3280;
    wire new_Jinkela_wire_1505;
    wire new_Jinkela_wire_167;
    wire _0358_;
    wire new_Jinkela_wire_259;
    wire _0233_;
    wire new_Jinkela_wire_2574;
    wire new_net_3;
    wire _0034_;
    wire new_Jinkela_wire_569;
    wire new_Jinkela_wire_1294;
    wire new_Jinkela_wire_1742;
    wire _0282_;
    wire _0760_;
    wire _0446_;
    wire new_Jinkela_wire_1077;
    wire new_Jinkela_wire_163;
    wire new_Jinkela_wire_2971;
    wire new_Jinkela_wire_2162;
    wire new_Jinkela_wire_390;
    wire new_Jinkela_wire_1545;
    wire new_Jinkela_wire_1021;
    wire new_Jinkela_wire_2168;
    wire new_Jinkela_wire_2056;
    wire _0631_;
    wire new_Jinkela_wire_2855;
    wire new_Jinkela_wire_2041;
    wire new_Jinkela_wire_139;
    wire new_Jinkela_wire_3187;
    wire new_Jinkela_wire_1129;
    wire new_Jinkela_wire_1033;
    wire new_Jinkela_wire_546;
    wire new_Jinkela_wire_2486;
    wire new_Jinkela_wire_2025;
    wire new_Jinkela_wire_3225;
    wire new_Jinkela_wire_1263;
    wire new_Jinkela_wire_501;
    wire new_Jinkela_wire_2791;
    wire new_Jinkela_wire_3068;
    wire new_Jinkela_wire_1682;
    wire new_Jinkela_wire_3082;
    wire new_Jinkela_wire_2198;
    wire new_Jinkela_wire_1373;
    wire new_Jinkela_wire_2379;
    wire new_Jinkela_wire_2391;
    wire new_Jinkela_wire_3255;
    wire new_Jinkela_wire_745;
    wire new_Jinkela_wire_751;
    wire new_Jinkela_wire_1698;
    wire _0779_;
    wire _0420_;
    wire new_Jinkela_wire_2937;
    wire new_Jinkela_wire_2906;
    wire new_Jinkela_wire_736;
    wire new_Jinkela_wire_142;
    wire new_Jinkela_wire_402;
    wire new_Jinkela_wire_2523;
    wire _0645_;
    wire new_Jinkela_wire_2886;
    wire new_Jinkela_wire_1350;
    wire new_Jinkela_wire_1151;
    wire new_Jinkela_wire_560;
    wire new_Jinkela_wire_1205;
    wire new_Jinkela_wire_1271;
    wire _0610_;
    wire new_Jinkela_wire_659;
    wire new_Jinkela_wire_525;
    wire new_Jinkela_wire_1407;
    wire _0523_;
    wire new_Jinkela_wire_57;
    wire new_Jinkela_wire_162;
    wire new_Jinkela_wire_1174;
    wire new_Jinkela_wire_1838;
    wire new_Jinkela_wire_1853;
    wire new_Jinkela_wire_2780;
    wire new_Jinkela_wire_1284;
    wire new_Jinkela_wire_2395;
    wire new_Jinkela_wire_2648;
    wire _0699_;
    wire new_Jinkela_wire_3201;
    wire new_Jinkela_wire_1194;
    wire new_Jinkela_wire_1442;
    wire new_Jinkela_wire_3056;
    wire new_Jinkela_wire_1570;
    wire new_Jinkela_wire_766;
    wire new_Jinkela_wire_50;
    wire new_Jinkela_wire_2189;
    wire new_Jinkela_wire_2939;
    wire _0751_;
    wire _0067_;
    wire new_Jinkela_wire_2712;
    wire new_Jinkela_wire_2385;
    wire new_Jinkela_wire_2007;
    wire new_Jinkela_wire_1498;
    wire new_Jinkela_wire_583;
    wire new_Jinkela_wire_3206;
    wire new_Jinkela_wire_2473;
    wire new_Jinkela_wire_1612;
    wire _0637_;
    wire new_Jinkela_wire_2002;
    wire new_Jinkela_wire_2490;
    wire new_Jinkela_wire_691;
    wire new_Jinkela_wire_1395;
    wire new_Jinkela_wire_1298;
    wire new_Jinkela_wire_2748;
    wire new_Jinkela_wire_2750;
    wire new_Jinkela_wire_2767;
    wire new_Jinkela_wire_2472;
    wire new_Jinkela_wire_2;
    wire new_Jinkela_wire_2488;
    wire _0045_;
    wire new_Jinkela_wire_2896;
    wire _0491_;
    wire _0153_;
    wire new_Jinkela_wire_1313;
    wire new_Jinkela_wire_512;
    wire _0769_;
    wire new_Jinkela_wire_1119;
    wire new_Jinkela_wire_343;
    wire new_Jinkela_wire_2931;
    wire _0490_;
    wire new_Jinkela_wire_1688;
    wire new_Jinkela_wire_534;
    wire new_Jinkela_wire_1657;
    wire _0502_;
    wire new_Jinkela_wire_364;
    wire new_Jinkela_wire_989;
    wire new_Jinkela_wire_1643;
    wire _0438_;
    wire new_Jinkela_wire_771;
    wire new_Jinkela_wire_74;
    wire _0051_;
    wire new_Jinkela_wire_2474;
    wire new_Jinkela_wire_946;
    wire new_Jinkela_wire_12;
    wire new_Jinkela_wire_171;
    wire _0652_;
    wire new_Jinkela_wire_2325;
    wire new_Jinkela_wire_2328;
    wire new_Jinkela_wire_1496;
    wire _0060_;
    wire new_Jinkela_wire_1665;
    wire new_Jinkela_wire_2734;
    wire new_Jinkela_wire_280;
    wire new_Jinkela_wire_1881;
    wire _0098_;
    wire new_Jinkela_wire_2880;
    wire new_Jinkela_wire_3142;
    wire new_Jinkela_wire_2524;
    wire new_Jinkela_wire_2581;
    wire new_Jinkela_wire_2653;
    wire new_Jinkela_wire_627;
    wire new_Jinkela_wire_1178;
    wire new_Jinkela_wire_1169;
    wire new_Jinkela_wire_2071;
    wire _0535_;
    wire _0703_;
    wire new_Jinkela_wire_1751;
    wire _0457_;
    wire new_Jinkela_wire_734;
    wire new_Jinkela_wire_2131;
    wire new_Jinkela_wire_199;
    wire new_Jinkela_wire_2399;
    wire new_Jinkela_wire_191;
    wire _0624_;
    wire new_Jinkela_wire_1083;
    wire new_Jinkela_wire_646;
    wire new_Jinkela_wire_1548;
    wire new_Jinkela_wire_924;
    wire new_Jinkela_wire_3231;
    input G25;
    input G47;
    input G30;
    input G50;
    input G27;
    input G3;
    input G31;
    input G19;
    input G9;
    input G13;
    input G39;
    input G34;
    input G8;
    input G46;
    input G14;
    input G18;
    input G32;
    input G42;
    input G11;
    input G48;
    input G22;
    input G4;
    input G17;
    input G35;
    input G23;
    input G21;
    input G36;
    input G41;
    input G5;
    input G38;
    input G26;
    input G7;
    input G1;
    input G28;
    input G6;
    input G24;
    input G20;
    input G43;
    input G44;
    input G12;
    input G40;
    input G10;
    input G29;
    input G16;
    input G33;
    input G37;
    input G45;
    input G49;
    input G15;
    input G2;
    output G3528;
    output G3521;
    output G3527;
    output G3535;
    output G3531;
    output G3540;
    output G3520;
    output G3537;
    output G3538;
    output G3530;
    output G3519;
    output G3525;
    output G3539;
    output G3524;
    output G3533;
    output G3523;
    output G3522;
    output G3532;
    output G3529;
    output G3534;
    output G3526;
    output G3536;

    bfr new_Jinkela_buffer_206 (
        .din(new_Jinkela_wire_351),
        .dout(new_Jinkela_wire_352)
    );

    bfr new_Jinkela_buffer_263 (
        .din(new_Jinkela_wire_463),
        .dout(new_Jinkela_wire_464)
    );

    bfr new_Jinkela_buffer_207 (
        .din(new_Jinkela_wire_352),
        .dout(new_Jinkela_wire_353)
    );

    bfr new_Jinkela_buffer_262 (
        .din(new_Jinkela_wire_462),
        .dout(new_Jinkela_wire_463)
    );

    bfr new_Jinkela_buffer_246 (
        .din(new_Jinkela_wire_396),
        .dout(new_Jinkela_wire_397)
    );

    bfr new_Jinkela_buffer_208 (
        .din(new_Jinkela_wire_353),
        .dout(new_Jinkela_wire_354)
    );

    spl2 new_Jinkela_splitter_78 (
        .a(G23),
        .b(new_Jinkela_wire_486),
        .c(new_Jinkela_wire_487)
    );

    bfr new_Jinkela_buffer_209 (
        .din(new_Jinkela_wire_354),
        .dout(new_Jinkela_wire_355)
    );

    bfr new_Jinkela_buffer_247 (
        .din(new_Jinkela_wire_397),
        .dout(new_Jinkela_wire_398)
    );

    bfr new_Jinkela_buffer_210 (
        .din(new_Jinkela_wire_355),
        .dout(new_Jinkela_wire_356)
    );

    bfr new_Jinkela_buffer_248 (
        .din(new_Jinkela_wire_398),
        .dout(new_Jinkela_wire_399)
    );

    bfr new_Jinkela_buffer_211 (
        .din(new_Jinkela_wire_356),
        .dout(new_Jinkela_wire_357)
    );

    bfr new_Jinkela_buffer_212 (
        .din(new_Jinkela_wire_357),
        .dout(new_Jinkela_wire_358)
    );

    spl2 new_Jinkela_splitter_56 (
        .a(new_Jinkela_wire_399),
        .b(new_Jinkela_wire_400),
        .c(new_Jinkela_wire_401)
    );

    bfr new_Jinkela_buffer_213 (
        .din(new_Jinkela_wire_358),
        .dout(new_Jinkela_wire_359)
    );

    bfr new_Jinkela_buffer_249 (
        .din(new_Jinkela_wire_401),
        .dout(new_Jinkela_wire_402)
    );

    bfr new_Jinkela_buffer_214 (
        .din(new_Jinkela_wire_359),
        .dout(new_Jinkela_wire_360)
    );

    bfr new_Jinkela_buffer_215 (
        .din(new_Jinkela_wire_360),
        .dout(new_Jinkela_wire_361)
    );

    spl4L new_Jinkela_splitter_75 (
        .a(new_Jinkela_wire_475),
        .d(new_Jinkela_wire_476),
        .e(new_Jinkela_wire_477),
        .b(new_Jinkela_wire_478),
        .c(new_Jinkela_wire_479)
    );

    spl2 new_Jinkela_splitter_74 (
        .a(G35),
        .b(new_Jinkela_wire_473),
        .c(new_Jinkela_wire_475)
    );

    bfr new_Jinkela_buffer_216 (
        .din(new_Jinkela_wire_361),
        .dout(new_Jinkela_wire_362)
    );

    spl2 new_Jinkela_splitter_57 (
        .a(new_Jinkela_wire_402),
        .b(new_Jinkela_wire_403),
        .c(new_Jinkela_wire_404)
    );

    bfr new_Jinkela_buffer_217 (
        .din(new_Jinkela_wire_362),
        .dout(new_Jinkela_wire_363)
    );

    spl2 new_Jinkela_splitter_58 (
        .a(new_Jinkela_wire_404),
        .b(new_Jinkela_wire_405),
        .c(new_Jinkela_wire_406)
    );

    bfr new_Jinkela_buffer_218 (
        .din(new_Jinkela_wire_363),
        .dout(new_Jinkela_wire_364)
    );

    spl4L new_Jinkela_splitter_62 (
        .a(new_Jinkela_wire_416),
        .d(new_Jinkela_wire_417),
        .e(new_Jinkela_wire_418),
        .b(new_Jinkela_wire_419),
        .c(new_Jinkela_wire_420)
    );

    bfr new_Jinkela_buffer_219 (
        .din(new_Jinkela_wire_364),
        .dout(new_Jinkela_wire_365)
    );

    bfr new_Jinkela_buffer_251 (
        .din(new_Jinkela_wire_408),
        .dout(new_Jinkela_wire_409)
    );

    bfr new_Jinkela_buffer_220 (
        .din(new_Jinkela_wire_365),
        .dout(new_Jinkela_wire_366)
    );

    spl4L new_Jinkela_splitter_61 (
        .a(new_Jinkela_wire_411),
        .d(new_Jinkela_wire_412),
        .e(new_Jinkela_wire_413),
        .b(new_Jinkela_wire_414),
        .c(new_Jinkela_wire_415)
    );

    bfr new_Jinkela_buffer_221 (
        .din(new_Jinkela_wire_366),
        .dout(new_Jinkela_wire_367)
    );

    spl4L new_Jinkela_splitter_66 (
        .a(new_Jinkela_wire_431),
        .d(new_Jinkela_wire_432),
        .e(new_Jinkela_wire_433),
        .b(new_Jinkela_wire_434),
        .c(new_Jinkela_wire_435)
    );

    bfr new_Jinkela_buffer_222 (
        .din(new_Jinkela_wire_367),
        .dout(new_Jinkela_wire_368)
    );

    bfr new_Jinkela_buffer_223 (
        .din(new_Jinkela_wire_368),
        .dout(new_Jinkela_wire_369)
    );

    spl4L new_Jinkela_splitter_64 (
        .a(new_Jinkela_wire_426),
        .d(new_Jinkela_wire_427),
        .e(new_Jinkela_wire_431),
        .b(new_Jinkela_wire_436),
        .c(new_Jinkela_wire_441)
    );

    spl4L new_Jinkela_splitter_63 (
        .a(new_Jinkela_wire_421),
        .d(new_Jinkela_wire_422),
        .e(new_Jinkela_wire_423),
        .b(new_Jinkela_wire_424),
        .c(new_Jinkela_wire_425)
    );

    bfr new_Jinkela_buffer_224 (
        .din(new_Jinkela_wire_369),
        .dout(new_Jinkela_wire_370)
    );

    bfr new_Jinkela_buffer_271 (
        .din(new_Jinkela_wire_487),
        .dout(new_Jinkela_wire_488)
    );

    bfr new_Jinkela_buffer_225 (
        .din(new_Jinkela_wire_370),
        .dout(new_Jinkela_wire_371)
    );

    spl3L new_Jinkela_splitter_65 (
        .a(new_Jinkela_wire_427),
        .d(new_Jinkela_wire_428),
        .b(new_Jinkela_wire_429),
        .c(new_Jinkela_wire_430)
    );

    bfr new_Jinkela_buffer_226 (
        .din(new_Jinkela_wire_371),
        .dout(new_Jinkela_wire_372)
    );

    spl4L new_Jinkela_splitter_67 (
        .a(new_Jinkela_wire_436),
        .d(new_Jinkela_wire_437),
        .e(new_Jinkela_wire_438),
        .b(new_Jinkela_wire_439),
        .c(new_Jinkela_wire_440)
    );

    bfr new_Jinkela_buffer_498 (
        .din(_0557_),
        .dout(new_Jinkela_wire_892)
    );

    bfr new_Jinkela_buffer_1183 (
        .din(new_Jinkela_wire_1955),
        .dout(new_Jinkela_wire_1956)
    );

    bfr new_Jinkela_buffer_451 (
        .din(new_Jinkela_wire_844),
        .dout(new_Jinkela_wire_845)
    );

    bfr new_Jinkela_buffer_1177 (
        .din(new_Jinkela_wire_1949),
        .dout(new_Jinkela_wire_1950)
    );

    bfr new_Jinkela_buffer_454 (
        .din(new_Jinkela_wire_847),
        .dout(new_Jinkela_wire_848)
    );

    spl2 new_Jinkela_splitter_301 (
        .a(_0559_),
        .b(new_Jinkela_wire_2003),
        .c(new_Jinkela_wire_2004)
    );

    bfr new_Jinkela_buffer_1227 (
        .din(_0232_),
        .dout(new_Jinkela_wire_2005)
    );

    spl2 new_Jinkela_splitter_152 (
        .a(_0339_),
        .b(new_Jinkela_wire_898),
        .c(new_Jinkela_wire_899)
    );

    bfr new_Jinkela_buffer_1184 (
        .din(new_Jinkela_wire_1956),
        .dout(new_Jinkela_wire_1957)
    );

    spl3L new_Jinkela_splitter_153 (
        .a(_0456_),
        .d(new_Jinkela_wire_900),
        .b(new_Jinkela_wire_901),
        .c(new_Jinkela_wire_902)
    );

    bfr new_Jinkela_buffer_455 (
        .din(new_Jinkela_wire_848),
        .dout(new_Jinkela_wire_849)
    );

    bfr new_Jinkela_buffer_1210 (
        .din(new_Jinkela_wire_1985),
        .dout(new_Jinkela_wire_1986)
    );

    bfr new_Jinkela_buffer_499 (
        .din(new_Jinkela_wire_892),
        .dout(new_Jinkela_wire_893)
    );

    bfr new_Jinkela_buffer_1185 (
        .din(new_Jinkela_wire_1957),
        .dout(new_Jinkela_wire_1958)
    );

    bfr new_Jinkela_buffer_456 (
        .din(new_Jinkela_wire_849),
        .dout(new_Jinkela_wire_850)
    );

    bfr new_Jinkela_buffer_1229 (
        .din(_0500_),
        .dout(new_Jinkela_wire_2007)
    );

    spl3L new_Jinkela_splitter_156 (
        .a(_0464_),
        .d(new_Jinkela_wire_909),
        .b(new_Jinkela_wire_910),
        .c(new_Jinkela_wire_911)
    );

    bfr new_Jinkela_buffer_1186 (
        .din(new_Jinkela_wire_1958),
        .dout(new_Jinkela_wire_1959)
    );

    bfr new_Jinkela_buffer_457 (
        .din(new_Jinkela_wire_850),
        .dout(new_Jinkela_wire_851)
    );

    bfr new_Jinkela_buffer_1211 (
        .din(new_Jinkela_wire_1986),
        .dout(new_Jinkela_wire_1987)
    );

    bfr new_Jinkela_buffer_500 (
        .din(new_Jinkela_wire_893),
        .dout(new_Jinkela_wire_894)
    );

    bfr new_Jinkela_buffer_1187 (
        .din(new_Jinkela_wire_1959),
        .dout(new_Jinkela_wire_1960)
    );

    bfr new_Jinkela_buffer_458 (
        .din(new_Jinkela_wire_851),
        .dout(new_Jinkela_wire_852)
    );

    bfr new_Jinkela_buffer_1188 (
        .din(new_Jinkela_wire_1960),
        .dout(new_Jinkela_wire_1961)
    );

    spl3L new_Jinkela_splitter_155 (
        .a(_0228_),
        .d(new_Jinkela_wire_906),
        .b(new_Jinkela_wire_907),
        .c(new_Jinkela_wire_908)
    );

    bfr new_Jinkela_buffer_459 (
        .din(new_Jinkela_wire_852),
        .dout(new_Jinkela_wire_853)
    );

    bfr new_Jinkela_buffer_1212 (
        .din(new_Jinkela_wire_1987),
        .dout(new_Jinkela_wire_1988)
    );

    bfr new_Jinkela_buffer_501 (
        .din(new_Jinkela_wire_894),
        .dout(new_Jinkela_wire_895)
    );

    bfr new_Jinkela_buffer_1189 (
        .din(new_Jinkela_wire_1961),
        .dout(new_Jinkela_wire_1962)
    );

    bfr new_Jinkela_buffer_460 (
        .din(new_Jinkela_wire_853),
        .dout(new_Jinkela_wire_854)
    );

    bfr new_Jinkela_buffer_1228 (
        .din(_0026_),
        .dout(new_Jinkela_wire_2006)
    );

    bfr new_Jinkela_buffer_1190 (
        .din(new_Jinkela_wire_1962),
        .dout(new_Jinkela_wire_1963)
    );

    bfr new_Jinkela_buffer_505 (
        .din(_0660_),
        .dout(new_Jinkela_wire_912)
    );

    bfr new_Jinkela_buffer_461 (
        .din(new_Jinkela_wire_854),
        .dout(new_Jinkela_wire_855)
    );

    bfr new_Jinkela_buffer_1213 (
        .din(new_Jinkela_wire_1988),
        .dout(new_Jinkela_wire_1989)
    );

    bfr new_Jinkela_buffer_502 (
        .din(new_Jinkela_wire_895),
        .dout(new_Jinkela_wire_896)
    );

    bfr new_Jinkela_buffer_1191 (
        .din(new_Jinkela_wire_1963),
        .dout(new_Jinkela_wire_1964)
    );

    bfr new_Jinkela_buffer_462 (
        .din(new_Jinkela_wire_855),
        .dout(new_Jinkela_wire_856)
    );

    spl2 new_Jinkela_splitter_302 (
        .a(_0735_),
        .b(new_Jinkela_wire_2008),
        .c(new_Jinkela_wire_2009)
    );

    spl2 new_Jinkela_splitter_303 (
        .a(_0244_),
        .b(new_Jinkela_wire_2010),
        .c(new_Jinkela_wire_2011)
    );

    bfr new_Jinkela_buffer_504 (
        .din(new_Jinkela_wire_902),
        .dout(new_Jinkela_wire_903)
    );

    bfr new_Jinkela_buffer_1192 (
        .din(new_Jinkela_wire_1964),
        .dout(new_Jinkela_wire_1965)
    );

    bfr new_Jinkela_buffer_507 (
        .din(_0201_),
        .dout(new_Jinkela_wire_914)
    );

    bfr new_Jinkela_buffer_463 (
        .din(new_Jinkela_wire_856),
        .dout(new_Jinkela_wire_857)
    );

    bfr new_Jinkela_buffer_1214 (
        .din(new_Jinkela_wire_1989),
        .dout(new_Jinkela_wire_1990)
    );

    bfr new_Jinkela_buffer_503 (
        .din(new_Jinkela_wire_896),
        .dout(new_Jinkela_wire_897)
    );

    bfr new_Jinkela_buffer_1193 (
        .din(new_Jinkela_wire_1965),
        .dout(new_Jinkela_wire_1966)
    );

    bfr new_Jinkela_buffer_464 (
        .din(new_Jinkela_wire_857),
        .dout(new_Jinkela_wire_858)
    );

    bfr new_Jinkela_buffer_1194 (
        .din(new_Jinkela_wire_1966),
        .dout(new_Jinkela_wire_1967)
    );

    bfr new_Jinkela_buffer_465 (
        .din(new_Jinkela_wire_858),
        .dout(new_Jinkela_wire_859)
    );

    bfr new_Jinkela_buffer_1215 (
        .din(new_Jinkela_wire_1990),
        .dout(new_Jinkela_wire_1991)
    );

    spl2 new_Jinkela_splitter_154 (
        .a(new_Jinkela_wire_903),
        .b(new_Jinkela_wire_904),
        .c(new_Jinkela_wire_905)
    );

    bfr new_Jinkela_buffer_1195 (
        .din(new_Jinkela_wire_1967),
        .dout(new_Jinkela_wire_1968)
    );

    bfr new_Jinkela_buffer_466 (
        .din(new_Jinkela_wire_859),
        .dout(new_Jinkela_wire_860)
    );

    bfr new_Jinkela_buffer_506 (
        .din(new_Jinkela_wire_912),
        .dout(new_Jinkela_wire_913)
    );

    bfr new_Jinkela_buffer_1196 (
        .din(new_Jinkela_wire_1968),
        .dout(new_Jinkela_wire_1969)
    );

    bfr new_Jinkela_buffer_467 (
        .din(new_Jinkela_wire_860),
        .dout(new_Jinkela_wire_861)
    );

    bfr new_Jinkela_buffer_1216 (
        .din(new_Jinkela_wire_1991),
        .dout(new_Jinkela_wire_1992)
    );

    bfr new_Jinkela_buffer_1197 (
        .din(new_Jinkela_wire_1969),
        .dout(new_Jinkela_wire_1970)
    );

    bfr new_Jinkela_buffer_468 (
        .din(new_Jinkela_wire_861),
        .dout(new_Jinkela_wire_862)
    );

    spl2 new_Jinkela_splitter_304 (
        .a(_0558_),
        .b(new_Jinkela_wire_2012),
        .c(new_Jinkela_wire_2013)
    );

    bfr new_Jinkela_buffer_1231 (
        .din(new_Jinkela_wire_2014),
        .dout(new_Jinkela_wire_2015)
    );

    bfr new_Jinkela_buffer_510 (
        .din(_0299_),
        .dout(new_Jinkela_wire_917)
    );

    bfr new_Jinkela_buffer_1198 (
        .din(new_Jinkela_wire_1970),
        .dout(new_Jinkela_wire_1971)
    );

    bfr new_Jinkela_buffer_469 (
        .din(new_Jinkela_wire_862),
        .dout(new_Jinkela_wire_863)
    );

    bfr new_Jinkela_buffer_1217 (
        .din(new_Jinkela_wire_1992),
        .dout(new_Jinkela_wire_1993)
    );

    bfr new_Jinkela_buffer_508 (
        .din(new_Jinkela_wire_914),
        .dout(new_Jinkela_wire_915)
    );

    bfr new_Jinkela_buffer_1199 (
        .din(new_Jinkela_wire_1971),
        .dout(new_Jinkela_wire_1972)
    );

    bfr new_Jinkela_buffer_470 (
        .din(new_Jinkela_wire_863),
        .dout(new_Jinkela_wire_864)
    );

    bfr new_Jinkela_buffer_1230 (
        .din(_0234_),
        .dout(new_Jinkela_wire_2014)
    );

    bfr new_Jinkela_buffer_1238 (
        .din(_0360_),
        .dout(new_Jinkela_wire_2026)
    );

    spl2 new_Jinkela_splitter_157 (
        .a(_0354_),
        .b(new_Jinkela_wire_918),
        .c(new_Jinkela_wire_919)
    );

    bfr new_Jinkela_buffer_1200 (
        .din(new_Jinkela_wire_1972),
        .dout(new_Jinkela_wire_1973)
    );

    bfr new_Jinkela_buffer_511 (
        .din(_0383_),
        .dout(new_Jinkela_wire_920)
    );

    bfr new_Jinkela_buffer_471 (
        .din(new_Jinkela_wire_864),
        .dout(new_Jinkela_wire_865)
    );

    bfr new_Jinkela_buffer_1218 (
        .din(new_Jinkela_wire_1993),
        .dout(new_Jinkela_wire_1994)
    );

    bfr new_Jinkela_buffer_509 (
        .din(new_Jinkela_wire_915),
        .dout(new_Jinkela_wire_916)
    );

    bfr new_Jinkela_buffer_1201 (
        .din(new_Jinkela_wire_1973),
        .dout(new_Jinkela_wire_1974)
    );

    bfr new_Jinkela_buffer_472 (
        .din(new_Jinkela_wire_865),
        .dout(new_Jinkela_wire_866)
    );

    bfr new_Jinkela_buffer_1234 (
        .din(_0349_),
        .dout(new_Jinkela_wire_2018)
    );

    spl2 new_Jinkela_splitter_160 (
        .a(_0142_),
        .b(new_Jinkela_wire_933),
        .c(new_Jinkela_wire_934)
    );

    bfr new_Jinkela_buffer_1202 (
        .din(new_Jinkela_wire_1974),
        .dout(new_Jinkela_wire_1975)
    );

    bfr new_Jinkela_buffer_519 (
        .din(_0249_),
        .dout(new_Jinkela_wire_935)
    );

    bfr new_Jinkela_buffer_473 (
        .din(new_Jinkela_wire_866),
        .dout(new_Jinkela_wire_867)
    );

    bfr new_Jinkela_buffer_1219 (
        .din(new_Jinkela_wire_1994),
        .dout(new_Jinkela_wire_1995)
    );

    bfr new_Jinkela_buffer_1203 (
        .din(new_Jinkela_wire_1975),
        .dout(new_Jinkela_wire_1976)
    );

    and_bi _0911_ (
        .a(new_Jinkela_wire_2565),
        .b(new_Jinkela_wire_937),
        .c(_0083_)
    );

    bfr new_Jinkela_buffer_423 (
        .din(G2),
        .dout(new_Jinkela_wire_792)
    );

    spl2 new_Jinkela_splitter_145 (
        .a(_0109_),
        .b(new_Jinkela_wire_804),
        .c(new_Jinkela_wire_805)
    );

    or_bb _0912_ (
        .a(_0083_),
        .b(new_Jinkela_wire_2089),
        .c(_0084_)
    );

    bfr new_Jinkela_buffer_416 (
        .din(new_Jinkela_wire_784),
        .dout(new_Jinkela_wire_785)
    );

    and_ii _0913_ (
        .a(new_Jinkela_wire_486),
        .b(new_Jinkela_wire_645),
        .c(_0085_)
    );

    bfr new_Jinkela_buffer_421 (
        .din(new_Jinkela_wire_789),
        .dout(new_Jinkela_wire_790)
    );

    or_bb _0914_ (
        .a(new_Jinkela_wire_3063),
        .b(new_Jinkela_wire_936),
        .c(_0086_)
    );

    and_bi _0915_ (
        .a(new_Jinkela_wire_2088),
        .b(_0086_),
        .c(_0087_)
    );

    spl4L new_Jinkela_splitter_142 (
        .a(new_Jinkela_wire_792),
        .d(new_Jinkela_wire_793),
        .e(new_Jinkela_wire_794),
        .b(new_Jinkela_wire_795),
        .c(new_Jinkela_wire_796)
    );

    and_bi _0916_ (
        .a(new_Jinkela_wire_1229),
        .b(new_Jinkela_wire_2370),
        .c(_0088_)
    );

    bfr new_Jinkela_buffer_429 (
        .din(_0605_),
        .dout(new_Jinkela_wire_810)
    );

    or_bb _0917_ (
        .a(new_Jinkela_wire_2169),
        .b(new_Jinkela_wire_1061),
        .c(_0089_)
    );

    spl2 new_Jinkela_splitter_146 (
        .a(_0205_),
        .b(new_Jinkela_wire_806),
        .c(new_Jinkela_wire_807)
    );

    and_bi _0918_ (
        .a(new_Jinkela_wire_1055),
        .b(new_Jinkela_wire_3305),
        .c(_0090_)
    );

    or_bi _0919_ (
        .a(new_Jinkela_wire_2914),
        .b(_0089_),
        .c(_0091_)
    );

    bfr new_Jinkela_buffer_424 (
        .din(new_Jinkela_wire_798),
        .dout(new_Jinkela_wire_799)
    );

    spl2 new_Jinkela_splitter_143 (
        .a(new_Jinkela_wire_796),
        .b(new_Jinkela_wire_797),
        .c(new_Jinkela_wire_798)
    );

    or_ii _0920_ (
        .a(new_Jinkela_wire_2781),
        .b(new_Jinkela_wire_166),
        .c(_0092_)
    );

    bfr new_Jinkela_buffer_427 (
        .din(new_Jinkela_wire_807),
        .dout(new_Jinkela_wire_808)
    );

    inv _0921_ (
        .din(new_Jinkela_wire_196),
        .dout(_0093_)
    );

    bfr new_Jinkela_buffer_440 (
        .din(_0095_),
        .dout(new_Jinkela_wire_821)
    );

    spl3L new_Jinkela_splitter_148 (
        .a(_0571_),
        .d(new_Jinkela_wire_830),
        .b(new_Jinkela_wire_831),
        .c(new_Jinkela_wire_832)
    );

    and_bi _0922_ (
        .a(new_Jinkela_wire_1939),
        .b(new_Jinkela_wire_3328),
        .c(_0094_)
    );

    bfr new_Jinkela_buffer_430 (
        .din(new_Jinkela_wire_810),
        .dout(new_Jinkela_wire_811)
    );

    spl2 new_Jinkela_splitter_144 (
        .a(new_Jinkela_wire_799),
        .b(new_Jinkela_wire_800),
        .c(new_Jinkela_wire_801)
    );

    and_bi _0923_ (
        .a(new_Jinkela_wire_393),
        .b(new_Jinkela_wire_152),
        .c(_0095_)
    );

    bfr new_Jinkela_buffer_425 (
        .din(new_Jinkela_wire_801),
        .dout(new_Jinkela_wire_802)
    );

    and_bi _0924_ (
        .a(new_Jinkela_wire_822),
        .b(new_Jinkela_wire_446),
        .c(_0096_)
    );

    bfr new_Jinkela_buffer_428 (
        .din(new_Jinkela_wire_808),
        .dout(new_Jinkela_wire_809)
    );

    or_bb _0925_ (
        .a(new_Jinkela_wire_1192),
        .b(_0094_),
        .c(_0097_)
    );

    and_bi _0926_ (
        .a(new_Jinkela_wire_846),
        .b(_0097_),
        .c(_0098_)
    );

    bfr new_Jinkela_buffer_447 (
        .din(_0685_),
        .dout(new_Jinkela_wire_833)
    );

    bfr new_Jinkela_buffer_426 (
        .din(new_Jinkela_wire_802),
        .dout(new_Jinkela_wire_803)
    );

    and_bi _0927_ (
        .a(new_Jinkela_wire_3320),
        .b(_0098_),
        .c(_0099_)
    );

    or_bi _0928_ (
        .a(_0099_),
        .b(_0091_),
        .c(_0100_)
    );

    bfr new_Jinkela_buffer_431 (
        .din(new_Jinkela_wire_811),
        .dout(new_Jinkela_wire_812)
    );

    or_bi _0929_ (
        .a(new_Jinkela_wire_3220),
        .b(new_Jinkela_wire_177),
        .c(_0101_)
    );

    spl2 new_Jinkela_splitter_147 (
        .a(new_Jinkela_wire_821),
        .b(new_Jinkela_wire_822),
        .c(new_Jinkela_wire_823)
    );

    and_bi _0930_ (
        .a(new_Jinkela_wire_754),
        .b(new_Jinkela_wire_3035),
        .c(_0102_)
    );

    bfr new_Jinkela_buffer_432 (
        .din(new_Jinkela_wire_812),
        .dout(new_Jinkela_wire_813)
    );

    or_bb _0931_ (
        .a(new_Jinkela_wire_409),
        .b(new_Jinkela_wire_332),
        .c(_0103_)
    );

    bfr new_Jinkela_buffer_441 (
        .din(new_Jinkela_wire_823),
        .dout(new_Jinkela_wire_824)
    );

    and_bi _0932_ (
        .a(new_Jinkela_wire_425),
        .b(new_Jinkela_wire_39),
        .c(_0104_)
    );

    bfr new_Jinkela_buffer_433 (
        .din(new_Jinkela_wire_813),
        .dout(new_Jinkela_wire_814)
    );

    and_bi _0933_ (
        .a(new_Jinkela_wire_3177),
        .b(new_Jinkela_wire_2824),
        .c(_0105_)
    );

    bfr new_Jinkela_buffer_448 (
        .din(_0121_),
        .dout(new_Jinkela_wire_834)
    );

    or_bb _0934_ (
        .a(new_Jinkela_wire_1675),
        .b(_0102_),
        .c(_0106_)
    );

    bfr new_Jinkela_buffer_434 (
        .din(new_Jinkela_wire_814),
        .dout(new_Jinkela_wire_815)
    );

    and_bi _0935_ (
        .a(new_Jinkela_wire_3044),
        .b(_0106_),
        .c(_0107_)
    );

    spl2 new_Jinkela_splitter_149 (
        .a(_0162_),
        .b(new_Jinkela_wire_835),
        .c(new_Jinkela_wire_836)
    );

    and_bi _0936_ (
        .a(new_Jinkela_wire_1047),
        .b(_0107_),
        .c(_0108_)
    );

    bfr new_Jinkela_buffer_435 (
        .din(new_Jinkela_wire_815),
        .dout(new_Jinkela_wire_816)
    );

    or_bb _0937_ (
        .a(new_Jinkela_wire_1289),
        .b(new_Jinkela_wire_841),
        .c(_0109_)
    );

    spl2 new_Jinkela_splitter_151 (
        .a(_0395_),
        .b(new_Jinkela_wire_842),
        .c(new_Jinkela_wire_843)
    );

    bfr new_Jinkela_buffer_442 (
        .din(new_Jinkela_wire_824),
        .dout(new_Jinkela_wire_825)
    );

    and_bi _0938_ (
        .a(new_Jinkela_wire_2570),
        .b(new_Jinkela_wire_805),
        .c(_0110_)
    );

    bfr new_Jinkela_buffer_436 (
        .din(new_Jinkela_wire_816),
        .dout(new_Jinkela_wire_817)
    );

    or_bb _0939_ (
        .a(_0110_),
        .b(new_Jinkela_wire_1293),
        .c(_0111_)
    );

    bfr new_Jinkela_buffer_449 (
        .din(_0293_),
        .dout(new_Jinkela_wire_837)
    );

    or_bb _0940_ (
        .a(new_Jinkela_wire_804),
        .b(new_Jinkela_wire_3060),
        .c(_0112_)
    );

    bfr new_Jinkela_buffer_437 (
        .din(new_Jinkela_wire_817),
        .dout(new_Jinkela_wire_818)
    );

    and_bi _0941_ (
        .a(new_Jinkela_wire_1292),
        .b(_0112_),
        .c(_0113_)
    );

    bfr new_Jinkela_buffer_443 (
        .din(new_Jinkela_wire_825),
        .dout(new_Jinkela_wire_826)
    );

    and_bi _0942_ (
        .a(new_Jinkela_wire_1099),
        .b(new_Jinkela_wire_2283),
        .c(_0114_)
    );

    bfr new_Jinkela_buffer_438 (
        .din(new_Jinkela_wire_818),
        .dout(new_Jinkela_wire_819)
    );

    and_bb _0943_ (
        .a(new_Jinkela_wire_1364),
        .b(new_Jinkela_wire_2032),
        .c(_0115_)
    );

    inv _0944_ (
        .din(new_Jinkela_wire_736),
        .dout(_0116_)
    );

    bfr new_Jinkela_buffer_439 (
        .din(new_Jinkela_wire_819),
        .dout(new_Jinkela_wire_820)
    );

    and_bi _0945_ (
        .a(new_Jinkela_wire_3312),
        .b(new_Jinkela_wire_2952),
        .c(_0117_)
    );

    bfr new_Jinkela_buffer_444 (
        .din(new_Jinkela_wire_826),
        .dout(new_Jinkela_wire_827)
    );

    and_ii _0946_ (
        .a(new_Jinkela_wire_3190),
        .b(new_Jinkela_wire_2168),
        .c(_0118_)
    );

    or_bb _0947_ (
        .a(_0118_),
        .b(new_Jinkela_wire_2764),
        .c(_0119_)
    );

    spl4L new_Jinkela_splitter_150 (
        .a(_0072_),
        .d(new_Jinkela_wire_838),
        .e(new_Jinkela_wire_839),
        .b(new_Jinkela_wire_840),
        .c(new_Jinkela_wire_841)
    );

    bfr new_Jinkela_buffer_445 (
        .din(new_Jinkela_wire_827),
        .dout(new_Jinkela_wire_828)
    );

    and_bi _0948_ (
        .a(new_Jinkela_wire_3302),
        .b(new_Jinkela_wire_746),
        .c(_0120_)
    );

    or_bb _0949_ (
        .a(new_Jinkela_wire_1281),
        .b(new_Jinkela_wire_273),
        .c(_0121_)
    );

    bfr new_Jinkela_buffer_453 (
        .din(new_net_1481),
        .dout(new_Jinkela_wire_847)
    );

    bfr new_Jinkela_buffer_446 (
        .din(new_Jinkela_wire_828),
        .dout(new_Jinkela_wire_829)
    );

    and_bi _0950_ (
        .a(new_Jinkela_wire_2053),
        .b(new_Jinkela_wire_3333),
        .c(_0122_)
    );

    and_bi _0951_ (
        .a(new_Jinkela_wire_834),
        .b(_0122_),
        .c(_0123_)
    );

    bfr new_Jinkela_buffer_452 (
        .din(_0092_),
        .dout(new_Jinkela_wire_846)
    );

    and_bi _0952_ (
        .a(new_Jinkela_wire_3316),
        .b(_0123_),
        .c(_0124_)
    );

    bfr new_Jinkela_buffer_450 (
        .din(new_Jinkela_wire_843),
        .dout(new_Jinkela_wire_844)
    );

    bfr new_Jinkela_buffer_227 (
        .din(new_Jinkela_wire_372),
        .dout(new_Jinkela_wire_373)
    );

    bfr new_Jinkela_buffer_356 (
        .din(new_Jinkela_wire_655),
        .dout(new_Jinkela_wire_656)
    );

    bfr new_Jinkela_buffer_2086 (
        .din(_0502_),
        .dout(new_Jinkela_wire_3310)
    );

    spl2 new_Jinkela_splitter_69 (
        .a(new_Jinkela_wire_445),
        .b(new_Jinkela_wire_446),
        .c(new_Jinkela_wire_447)
    );

    spl3L new_Jinkela_splitter_466 (
        .a(new_Jinkela_wire_3270),
        .d(new_Jinkela_wire_3271),
        .b(new_Jinkela_wire_3272),
        .c(new_Jinkela_wire_3273)
    );

    bfr new_Jinkela_buffer_228 (
        .din(new_Jinkela_wire_373),
        .dout(new_Jinkela_wire_374)
    );

    spl4L new_Jinkela_splitter_470 (
        .a(new_Jinkela_wire_3303),
        .d(new_Jinkela_wire_3304),
        .e(new_Jinkela_wire_3305),
        .b(new_Jinkela_wire_3306),
        .c(new_Jinkela_wire_3307)
    );

    bfr new_Jinkela_buffer_357 (
        .din(new_Jinkela_wire_656),
        .dout(new_Jinkela_wire_657)
    );

    bfr new_Jinkela_buffer_2080 (
        .din(new_Jinkela_wire_3293),
        .dout(new_Jinkela_wire_3294)
    );

    spl4L new_Jinkela_splitter_68 (
        .a(new_Jinkela_wire_441),
        .d(new_Jinkela_wire_442),
        .e(new_Jinkela_wire_443),
        .b(new_Jinkela_wire_444),
        .c(new_Jinkela_wire_445)
    );

    bfr new_Jinkela_buffer_2063 (
        .din(new_Jinkela_wire_3273),
        .dout(new_Jinkela_wire_3274)
    );

    bfr new_Jinkela_buffer_363 (
        .din(new_Jinkela_wire_664),
        .dout(new_Jinkela_wire_665)
    );

    bfr new_Jinkela_buffer_229 (
        .din(new_Jinkela_wire_374),
        .dout(new_Jinkela_wire_375)
    );

    spl4L new_Jinkela_splitter_122 (
        .a(new_Jinkela_wire_704),
        .d(new_Jinkela_wire_705),
        .e(new_Jinkela_wire_706),
        .b(new_Jinkela_wire_707),
        .c(new_Jinkela_wire_708)
    );

    spl2 new_Jinkela_splitter_113 (
        .a(new_Jinkela_wire_657),
        .b(new_Jinkela_wire_658),
        .c(new_Jinkela_wire_659)
    );

    spl4L new_Jinkela_splitter_469 (
        .a(new_Jinkela_wire_3298),
        .d(new_Jinkela_wire_3299),
        .e(new_Jinkela_wire_3300),
        .b(new_Jinkela_wire_3301),
        .c(new_Jinkela_wire_3302)
    );

    bfr new_Jinkela_buffer_272 (
        .din(G21),
        .dout(new_Jinkela_wire_489)
    );

    bfr new_Jinkela_buffer_2064 (
        .din(new_Jinkela_wire_3274),
        .dout(new_Jinkela_wire_3275)
    );

    bfr new_Jinkela_buffer_264 (
        .din(new_Jinkela_wire_464),
        .dout(new_Jinkela_wire_465)
    );

    bfr new_Jinkela_buffer_364 (
        .din(new_Jinkela_wire_665),
        .dout(new_Jinkela_wire_666)
    );

    bfr new_Jinkela_buffer_230 (
        .din(new_Jinkela_wire_375),
        .dout(new_Jinkela_wire_376)
    );

    bfr new_Jinkela_buffer_2081 (
        .din(new_Jinkela_wire_3294),
        .dout(new_Jinkela_wire_3295)
    );

    bfr new_Jinkela_buffer_2065 (
        .din(new_Jinkela_wire_3275),
        .dout(new_Jinkela_wire_3276)
    );

    bfr new_Jinkela_buffer_371 (
        .din(new_Jinkela_wire_680),
        .dout(new_Jinkela_wire_681)
    );

    bfr new_Jinkela_buffer_231 (
        .din(new_Jinkela_wire_376),
        .dout(new_Jinkela_wire_377)
    );

    bfr new_Jinkela_buffer_365 (
        .din(new_Jinkela_wire_666),
        .dout(new_Jinkela_wire_667)
    );

    bfr new_Jinkela_buffer_252 (
        .din(new_Jinkela_wire_447),
        .dout(new_Jinkela_wire_448)
    );

    bfr new_Jinkela_buffer_2066 (
        .din(new_Jinkela_wire_3276),
        .dout(new_Jinkela_wire_3277)
    );

    bfr new_Jinkela_buffer_232 (
        .din(new_Jinkela_wire_377),
        .dout(new_Jinkela_wire_378)
    );

    bfr new_Jinkela_buffer_393 (
        .din(new_Jinkela_wire_732),
        .dout(new_Jinkela_wire_733)
    );

    spl3L new_Jinkela_splitter_114 (
        .a(new_Jinkela_wire_667),
        .d(new_Jinkela_wire_668),
        .b(new_Jinkela_wire_669),
        .c(new_Jinkela_wire_670)
    );

    bfr new_Jinkela_buffer_2082 (
        .din(new_Jinkela_wire_3295),
        .dout(new_Jinkela_wire_3296)
    );

    bfr new_Jinkela_buffer_280 (
        .din(G36),
        .dout(new_Jinkela_wire_508)
    );

    bfr new_Jinkela_buffer_2067 (
        .din(new_Jinkela_wire_3277),
        .dout(new_Jinkela_wire_3278)
    );

    bfr new_Jinkela_buffer_265 (
        .din(new_Jinkela_wire_465),
        .dout(new_Jinkela_wire_466)
    );

    bfr new_Jinkela_buffer_372 (
        .din(new_Jinkela_wire_681),
        .dout(new_Jinkela_wire_682)
    );

    bfr new_Jinkela_buffer_233 (
        .din(new_Jinkela_wire_378),
        .dout(new_Jinkela_wire_379)
    );

    spl3L new_Jinkela_splitter_115 (
        .a(new_Jinkela_wire_670),
        .d(new_Jinkela_wire_671),
        .b(new_Jinkela_wire_672),
        .c(new_Jinkela_wire_673)
    );

    bfr new_Jinkela_buffer_2068 (
        .din(new_Jinkela_wire_3278),
        .dout(new_Jinkela_wire_3279)
    );

    spl2 new_Jinkela_splitter_76 (
        .a(new_Jinkela_wire_479),
        .b(new_Jinkela_wire_480),
        .c(new_Jinkela_wire_481)
    );

    bfr new_Jinkela_buffer_378 (
        .din(new_Jinkela_wire_691),
        .dout(new_Jinkela_wire_692)
    );

    bfr new_Jinkela_buffer_234 (
        .din(new_Jinkela_wire_379),
        .dout(new_Jinkela_wire_380)
    );

    bfr new_Jinkela_buffer_366 (
        .din(new_Jinkela_wire_673),
        .dout(new_Jinkela_wire_674)
    );

    bfr new_Jinkela_buffer_2083 (
        .din(new_Jinkela_wire_3296),
        .dout(new_Jinkela_wire_3297)
    );

    bfr new_Jinkela_buffer_253 (
        .din(new_Jinkela_wire_448),
        .dout(new_Jinkela_wire_449)
    );

    bfr new_Jinkela_buffer_2069 (
        .din(new_Jinkela_wire_3279),
        .dout(new_Jinkela_wire_3280)
    );

    bfr new_Jinkela_buffer_373 (
        .din(new_Jinkela_wire_682),
        .dout(new_Jinkela_wire_683)
    );

    bfr new_Jinkela_buffer_235 (
        .din(new_Jinkela_wire_380),
        .dout(new_Jinkela_wire_381)
    );

    bfr new_Jinkela_buffer_367 (
        .din(new_Jinkela_wire_674),
        .dout(new_Jinkela_wire_675)
    );

    bfr new_Jinkela_buffer_2070 (
        .din(new_Jinkela_wire_3280),
        .dout(new_Jinkela_wire_3281)
    );

    spl3L new_Jinkela_splitter_123 (
        .a(new_Jinkela_wire_708),
        .d(new_Jinkela_wire_709),
        .b(new_Jinkela_wire_710),
        .c(new_Jinkela_wire_711)
    );

    bfr new_Jinkela_buffer_236 (
        .din(new_Jinkela_wire_381),
        .dout(new_Jinkela_wire_382)
    );

    spl3L new_Jinkela_splitter_475 (
        .a(_0652_),
        .d(new_Jinkela_wire_3322),
        .b(new_Jinkela_wire_3323),
        .c(new_Jinkela_wire_3324)
    );

    bfr new_Jinkela_buffer_368 (
        .din(new_Jinkela_wire_675),
        .dout(new_Jinkela_wire_676)
    );

    bfr new_Jinkela_buffer_2085 (
        .din(new_Jinkela_wire_3308),
        .dout(new_Jinkela_wire_3309)
    );

    bfr new_Jinkela_buffer_254 (
        .din(new_Jinkela_wire_449),
        .dout(new_Jinkela_wire_450)
    );

    bfr new_Jinkela_buffer_2071 (
        .din(new_Jinkela_wire_3281),
        .dout(new_Jinkela_wire_3282)
    );

    bfr new_Jinkela_buffer_374 (
        .din(new_Jinkela_wire_683),
        .dout(new_Jinkela_wire_684)
    );

    bfr new_Jinkela_buffer_237 (
        .din(new_Jinkela_wire_382),
        .dout(new_Jinkela_wire_383)
    );

    bfr new_Jinkela_buffer_379 (
        .din(new_Jinkela_wire_692),
        .dout(new_Jinkela_wire_693)
    );

    spl3L new_Jinkela_splitter_471 (
        .a(_0051_),
        .d(new_Jinkela_wire_3311),
        .b(new_Jinkela_wire_3312),
        .c(new_Jinkela_wire_3313)
    );

    spl3L new_Jinkela_splitter_91 (
        .a(G5),
        .d(new_Jinkela_wire_534),
        .b(new_Jinkela_wire_535),
        .c(new_Jinkela_wire_536)
    );

    spl2 new_Jinkela_splitter_125 (
        .a(new_Jinkela_wire_714),
        .b(new_Jinkela_wire_715),
        .c(new_Jinkela_wire_716)
    );

    bfr new_Jinkela_buffer_2072 (
        .din(new_Jinkela_wire_3282),
        .dout(new_Jinkela_wire_3283)
    );

    bfr new_Jinkela_buffer_266 (
        .din(new_Jinkela_wire_466),
        .dout(new_Jinkela_wire_467)
    );

    bfr new_Jinkela_buffer_375 (
        .din(new_Jinkela_wire_684),
        .dout(new_Jinkela_wire_685)
    );

    bfr new_Jinkela_buffer_238 (
        .din(new_Jinkela_wire_383),
        .dout(new_Jinkela_wire_384)
    );

    bfr new_Jinkela_buffer_2087 (
        .din(new_Jinkela_wire_3324),
        .dout(new_Jinkela_wire_3325)
    );

    bfr new_Jinkela_buffer_255 (
        .din(new_Jinkela_wire_450),
        .dout(new_Jinkela_wire_451)
    );

    bfr new_Jinkela_buffer_2073 (
        .din(new_Jinkela_wire_3283),
        .dout(new_Jinkela_wire_3284)
    );

    spl2 new_Jinkela_splitter_117 (
        .a(new_Jinkela_wire_685),
        .b(new_Jinkela_wire_686),
        .c(new_Jinkela_wire_687)
    );

    bfr new_Jinkela_buffer_239 (
        .din(new_Jinkela_wire_384),
        .dout(new_Jinkela_wire_385)
    );

    spl3L new_Jinkela_splitter_473 (
        .a(new_Jinkela_wire_3315),
        .d(new_Jinkela_wire_3316),
        .b(new_Jinkela_wire_3317),
        .c(new_Jinkela_wire_3318)
    );

    bfr new_Jinkela_buffer_376 (
        .din(new_Jinkela_wire_687),
        .dout(new_Jinkela_wire_688)
    );

    bfr new_Jinkela_buffer_269 (
        .din(new_Jinkela_wire_481),
        .dout(new_Jinkela_wire_482)
    );

    bfr new_Jinkela_buffer_267 (
        .din(new_Jinkela_wire_467),
        .dout(new_Jinkela_wire_468)
    );

    bfr new_Jinkela_buffer_380 (
        .din(new_Jinkela_wire_693),
        .dout(new_Jinkela_wire_694)
    );

    spl2 new_Jinkela_splitter_476 (
        .a(_0060_),
        .b(new_Jinkela_wire_3327),
        .c(new_Jinkela_wire_3330)
    );

    bfr new_Jinkela_buffer_240 (
        .din(new_Jinkela_wire_385),
        .dout(new_Jinkela_wire_386)
    );

    spl2 new_Jinkela_splitter_121 (
        .a(new_Jinkela_wire_701),
        .b(new_Jinkela_wire_702),
        .c(new_Jinkela_wire_703)
    );

    spl2 new_Jinkela_splitter_70 (
        .a(new_Jinkela_wire_451),
        .b(new_Jinkela_wire_452),
        .c(new_Jinkela_wire_453)
    );

    spl2 new_Jinkela_splitter_124 (
        .a(G40),
        .b(new_Jinkela_wire_713),
        .c(new_Jinkela_wire_714)
    );

    spl3L new_Jinkela_splitter_474 (
        .a(new_Jinkela_wire_3318),
        .d(new_Jinkela_wire_3319),
        .b(new_Jinkela_wire_3320),
        .c(new_Jinkela_wire_3321)
    );

    bfr new_Jinkela_buffer_381 (
        .din(new_Jinkela_wire_694),
        .dout(new_Jinkela_wire_695)
    );

    spl2 new_Jinkela_splitter_472 (
        .a(new_Jinkela_wire_3313),
        .b(new_Jinkela_wire_3314),
        .c(new_Jinkela_wire_3315)
    );

    bfr new_Jinkela_buffer_241 (
        .din(new_Jinkela_wire_386),
        .dout(new_Jinkela_wire_387)
    );

    spl3L new_Jinkela_splitter_71 (
        .a(new_Jinkela_wire_453),
        .d(new_Jinkela_wire_454),
        .b(new_Jinkela_wire_455),
        .c(new_Jinkela_wire_456)
    );

    bfr new_Jinkela_buffer_382 (
        .din(new_Jinkela_wire_695),
        .dout(new_Jinkela_wire_696)
    );

    bfr new_Jinkela_buffer_242 (
        .din(new_Jinkela_wire_387),
        .dout(new_Jinkela_wire_388)
    );

    bfr new_Jinkela_buffer_2088 (
        .din(new_Jinkela_wire_3325),
        .dout(new_Jinkela_wire_3326)
    );

    bfr new_Jinkela_buffer_383 (
        .din(new_Jinkela_wire_696),
        .dout(new_Jinkela_wire_697)
    );

    spl4L new_Jinkela_splitter_478 (
        .a(new_Jinkela_wire_3330),
        .d(new_Jinkela_wire_3331),
        .e(new_Jinkela_wire_3332),
        .b(new_Jinkela_wire_3333),
        .c(new_Jinkela_wire_3334)
    );

    bfr new_Jinkela_buffer_243 (
        .din(new_Jinkela_wire_388),
        .dout(new_Jinkela_wire_389)
    );

    spl2 new_Jinkela_splitter_130 (
        .a(G10),
        .b(new_Jinkela_wire_732),
        .c(new_Jinkela_wire_734)
    );

    spl2 new_Jinkela_splitter_72 (
        .a(new_Jinkela_wire_468),
        .b(new_Jinkela_wire_469),
        .c(new_Jinkela_wire_470)
    );

    spl2 new_Jinkela_splitter_119 (
        .a(new_Jinkela_wire_697),
        .b(new_Jinkela_wire_698),
        .c(new_Jinkela_wire_699)
    );

    spl2 new_Jinkela_splitter_477 (
        .a(new_Jinkela_wire_3327),
        .b(new_Jinkela_wire_3328),
        .c(new_Jinkela_wire_3329)
    );

    bfr new_Jinkela_buffer_244 (
        .din(new_Jinkela_wire_389),
        .dout(new_Jinkela_wire_390)
    );

    bfr new_Jinkela_buffer_384 (
        .din(new_Jinkela_wire_699),
        .dout(new_Jinkela_wire_700)
    );

    bfr new_Jinkela_buffer_256 (
        .din(new_Jinkela_wire_456),
        .dout(new_Jinkela_wire_457)
    );

    bfr new_Jinkela_buffer_385 (
        .din(new_Jinkela_wire_711),
        .dout(new_Jinkela_wire_712)
    );

    spl2 new_Jinkela_splitter_73 (
        .a(new_Jinkela_wire_470),
        .b(new_Jinkela_wire_471),
        .c(new_Jinkela_wire_472)
    );

    bfr new_Jinkela_buffer_401 (
        .din(G16),
        .dout(new_Jinkela_wire_755)
    );

    bfr new_Jinkela_buffer_257 (
        .din(new_Jinkela_wire_457),
        .dout(new_Jinkela_wire_458)
    );

    bfr new_Jinkela_buffer_410 (
        .din(G33),
        .dout(new_Jinkela_wire_766)
    );

    spl2 new_Jinkela_splitter_126 (
        .a(new_Jinkela_wire_716),
        .b(new_Jinkela_wire_717),
        .c(new_Jinkela_wire_718)
    );

    bfr new_Jinkela_buffer_397 (
        .din(new_Jinkela_wire_748),
        .dout(new_Jinkela_wire_749)
    );

    spl4L new_Jinkela_splitter_84 (
        .a(new_Jinkela_wire_508),
        .d(new_Jinkela_wire_509),
        .e(new_Jinkela_wire_510),
        .b(new_Jinkela_wire_511),
        .c(new_Jinkela_wire_512)
    );

    spl4L new_Jinkela_splitter_131 (
        .a(new_Jinkela_wire_734),
        .d(new_Jinkela_wire_735),
        .e(new_Jinkela_wire_736),
        .b(new_Jinkela_wire_737),
        .c(new_Jinkela_wire_738)
    );

    bfr new_Jinkela_buffer_258 (
        .din(new_Jinkela_wire_458),
        .dout(new_Jinkela_wire_459)
    );

    bfr new_Jinkela_buffer_396 (
        .din(G29),
        .dout(new_Jinkela_wire_748)
    );

    bfr new_Jinkela_buffer_283 (
        .din(G41),
        .dout(new_Jinkela_wire_519)
    );

    bfr new_Jinkela_buffer_386 (
        .din(new_Jinkela_wire_718),
        .dout(new_Jinkela_wire_719)
    );

    bfr new_Jinkela_buffer_259 (
        .din(new_Jinkela_wire_459),
        .dout(new_Jinkela_wire_460)
    );

    spl3L new_Jinkela_splitter_308 (
        .a(_0088_),
        .d(new_Jinkela_wire_2032),
        .b(new_Jinkela_wire_2033),
        .c(new_Jinkela_wire_2034)
    );

    bfr new_Jinkela_buffer_1204 (
        .din(new_Jinkela_wire_1976),
        .dout(new_Jinkela_wire_1977)
    );

    bfr new_Jinkela_buffer_1220 (
        .din(new_Jinkela_wire_1995),
        .dout(new_Jinkela_wire_1996)
    );

    bfr new_Jinkela_buffer_1205 (
        .din(new_Jinkela_wire_1977),
        .dout(new_Jinkela_wire_1978)
    );

    bfr new_Jinkela_buffer_1232 (
        .din(new_Jinkela_wire_2015),
        .dout(new_Jinkela_wire_2016)
    );

    bfr new_Jinkela_buffer_1206 (
        .din(new_Jinkela_wire_1978),
        .dout(new_Jinkela_wire_1979)
    );

    bfr new_Jinkela_buffer_1221 (
        .din(new_Jinkela_wire_1996),
        .dout(new_Jinkela_wire_1997)
    );

    bfr new_Jinkela_buffer_1239 (
        .din(new_Jinkela_wire_2026),
        .dout(new_Jinkela_wire_2027)
    );

    bfr new_Jinkela_buffer_1222 (
        .din(new_Jinkela_wire_1997),
        .dout(new_Jinkela_wire_1998)
    );

    bfr new_Jinkela_buffer_1233 (
        .din(new_Jinkela_wire_2016),
        .dout(new_Jinkela_wire_2017)
    );

    bfr new_Jinkela_buffer_1223 (
        .din(new_Jinkela_wire_1998),
        .dout(new_Jinkela_wire_1999)
    );

    bfr new_Jinkela_buffer_1236 (
        .din(new_Jinkela_wire_2019),
        .dout(new_Jinkela_wire_2020)
    );

    bfr new_Jinkela_buffer_1224 (
        .din(new_Jinkela_wire_1999),
        .dout(new_Jinkela_wire_2000)
    );

    bfr new_Jinkela_buffer_1235 (
        .din(new_Jinkela_wire_2018),
        .dout(new_Jinkela_wire_2019)
    );

    bfr new_Jinkela_buffer_1225 (
        .din(new_Jinkela_wire_2000),
        .dout(new_Jinkela_wire_2001)
    );

    spl4L new_Jinkela_splitter_307 (
        .a(new_Jinkela_wire_2027),
        .d(new_Jinkela_wire_2028),
        .e(new_Jinkela_wire_2029),
        .b(new_Jinkela_wire_2030),
        .c(new_Jinkela_wire_2031)
    );

    spl2 new_Jinkela_splitter_305 (
        .a(new_Jinkela_wire_2020),
        .b(new_Jinkela_wire_2021),
        .c(new_Jinkela_wire_2022)
    );

    bfr new_Jinkela_buffer_1237 (
        .din(new_Jinkela_wire_2022),
        .dout(new_Jinkela_wire_2023)
    );

    bfr new_Jinkela_buffer_1241 (
        .din(_0646_),
        .dout(new_Jinkela_wire_2036)
    );

    bfr new_Jinkela_buffer_1240 (
        .din(_0715_),
        .dout(new_Jinkela_wire_2035)
    );

    bfr new_Jinkela_buffer_1248 (
        .din(_0177_),
        .dout(new_Jinkela_wire_2045)
    );

    spl2 new_Jinkela_splitter_306 (
        .a(new_Jinkela_wire_2023),
        .b(new_Jinkela_wire_2024),
        .c(new_Jinkela_wire_2025)
    );

    bfr new_Jinkela_buffer_1249 (
        .din(new_Jinkela_wire_2045),
        .dout(new_Jinkela_wire_2046)
    );

    bfr new_Jinkela_buffer_1242 (
        .din(_0644_),
        .dout(new_Jinkela_wire_2037)
    );

    bfr new_Jinkela_buffer_1250 (
        .din(_0620_),
        .dout(new_Jinkela_wire_2047)
    );

    bfr new_Jinkela_buffer_1243 (
        .din(new_Jinkela_wire_2037),
        .dout(new_Jinkela_wire_2038)
    );

    bfr new_Jinkela_buffer_1244 (
        .din(new_Jinkela_wire_2038),
        .dout(new_Jinkela_wire_2039)
    );

    bfr new_Jinkela_buffer_1245 (
        .din(new_Jinkela_wire_2039),
        .dout(new_Jinkela_wire_2040)
    );

    bfr new_Jinkela_buffer_1259 (
        .din(_0127_),
        .dout(new_Jinkela_wire_2065)
    );

    bfr new_Jinkela_buffer_1251 (
        .din(new_Jinkela_wire_2047),
        .dout(new_Jinkela_wire_2048)
    );

    bfr new_Jinkela_buffer_1246 (
        .din(new_Jinkela_wire_2040),
        .dout(new_Jinkela_wire_2041)
    );

    bfr new_Jinkela_buffer_1263 (
        .din(_0168_),
        .dout(new_Jinkela_wire_2071)
    );

    spl2 new_Jinkela_splitter_309 (
        .a(new_Jinkela_wire_2041),
        .b(new_Jinkela_wire_2042),
        .c(new_Jinkela_wire_2043)
    );

    bfr new_Jinkela_buffer_1247 (
        .din(new_Jinkela_wire_2043),
        .dout(new_Jinkela_wire_2044)
    );

    spl4L new_Jinkela_splitter_312 (
        .a(_0549_),
        .d(new_Jinkela_wire_2061),
        .e(new_Jinkela_wire_2062),
        .b(new_Jinkela_wire_2063),
        .c(new_Jinkela_wire_2064)
    );

    bfr new_Jinkela_buffer_1252 (
        .din(new_Jinkela_wire_2050),
        .dout(new_Jinkela_wire_2051)
    );

    spl2 new_Jinkela_splitter_310 (
        .a(new_Jinkela_wire_2048),
        .b(new_Jinkela_wire_2049),
        .c(new_Jinkela_wire_2050)
    );

    spl2 new_Jinkela_splitter_313 (
        .a(_0611_),
        .b(new_Jinkela_wire_2066),
        .c(new_Jinkela_wire_2067)
    );

    bfr new_Jinkela_buffer_1260 (
        .din(new_Jinkela_wire_2067),
        .dout(new_Jinkela_wire_2068)
    );

    spl3L new_Jinkela_splitter_311 (
        .a(new_Jinkela_wire_2051),
        .d(new_Jinkela_wire_2052),
        .b(new_Jinkela_wire_2053),
        .c(new_Jinkela_wire_2054)
    );

    spl2 new_Jinkela_splitter_315 (
        .a(_0332_),
        .b(new_Jinkela_wire_2077),
        .c(new_Jinkela_wire_2078)
    );

    and_bi _1289_ (
        .a(_0457_),
        .b(_0458_),
        .c(_0459_)
    );

    or_bi _1290_ (
        .a(new_Jinkela_wire_2736),
        .b(new_Jinkela_wire_1678),
        .c(_0460_)
    );

    and_bi _1291_ (
        .a(new_Jinkela_wire_2735),
        .b(new_Jinkela_wire_1677),
        .c(_0461_)
    );

    and_bi _1292_ (
        .a(_0460_),
        .b(_0461_),
        .c(_0462_)
    );

    and_bi _1293_ (
        .a(_0454_),
        .b(new_Jinkela_wire_1308),
        .c(_0463_)
    );

    or_bb _1294_ (
        .a(_0463_),
        .b(new_Jinkela_wire_1860),
        .c(new_net_0)
    );

    or_bb _1295_ (
        .a(new_Jinkela_wire_2289),
        .b(new_Jinkela_wire_3163),
        .c(_0464_)
    );

    or_bb _1296_ (
        .a(new_Jinkela_wire_2109),
        .b(new_Jinkela_wire_3068),
        .c(_0465_)
    );

    and_bi _1297_ (
        .a(new_Jinkela_wire_669),
        .b(new_Jinkela_wire_1876),
        .c(_0466_)
    );

    and_bi _1298_ (
        .a(new_Jinkela_wire_1057),
        .b(new_Jinkela_wire_1739),
        .c(_0467_)
    );

    and_bi _1299_ (
        .a(new_Jinkela_wire_190),
        .b(new_Jinkela_wire_2368),
        .c(_0468_)
    );

    or_bb _1300_ (
        .a(_0468_),
        .b(new_Jinkela_wire_3131),
        .c(_0469_)
    );

    or_bb _1301_ (
        .a(_0469_),
        .b(new_Jinkela_wire_1153),
        .c(_0470_)
    );

    and_bi _1302_ (
        .a(new_Jinkela_wire_1697),
        .b(new_Jinkela_wire_3011),
        .c(_0471_)
    );

    and_bi _1303_ (
        .a(new_Jinkela_wire_405),
        .b(new_Jinkela_wire_1132),
        .c(_0472_)
    );

    or_bb _1304_ (
        .a(_0472_),
        .b(new_Jinkela_wire_454),
        .c(_0473_)
    );

    and_bi _1305_ (
        .a(new_Jinkela_wire_301),
        .b(new_Jinkela_wire_1122),
        .c(_0474_)
    );

    or_bi _1306_ (
        .a(new_Jinkela_wire_490),
        .b(new_Jinkela_wire_192),
        .c(_0475_)
    );

    and_bi _1307_ (
        .a(new_Jinkela_wire_1472),
        .b(new_Jinkela_wire_2413),
        .c(_0476_)
    );

    or_bb _1308_ (
        .a(new_Jinkela_wire_2739),
        .b(_0474_),
        .c(_0477_)
    );

    or_bb _1309_ (
        .a(new_Jinkela_wire_2301),
        .b(new_Jinkela_wire_1644),
        .c(_0478_)
    );

    or_bb _1310_ (
        .a(_0478_),
        .b(_0471_),
        .c(_0479_)
    );

    or_bb _1311_ (
        .a(_0479_),
        .b(new_Jinkela_wire_939),
        .c(_0480_)
    );

    and_bi _1312_ (
        .a(new_Jinkela_wire_1714),
        .b(new_Jinkela_wire_1741),
        .c(_0481_)
    );

    or_bi _1313_ (
        .a(new_Jinkela_wire_1883),
        .b(new_Jinkela_wire_725),
        .c(_0482_)
    );

    and_bi _1314_ (
        .a(_0482_),
        .b(new_Jinkela_wire_2374),
        .c(_0483_)
    );

    and_bi _1315_ (
        .a(new_Jinkela_wire_533),
        .b(new_Jinkela_wire_2367),
        .c(_0484_)
    );

    and_ii _1316_ (
        .a(new_Jinkela_wire_1006),
        .b(new_Jinkela_wire_2429),
        .c(_0485_)
    );

    or_bb _1317_ (
        .a(new_Jinkela_wire_3133),
        .b(_0484_),
        .c(_0486_)
    );

    and_bi _1318_ (
        .a(new_Jinkela_wire_1861),
        .b(_0486_),
        .c(_0487_)
    );

    and_bi _1319_ (
        .a(new_Jinkela_wire_932),
        .b(new_Jinkela_wire_2999),
        .c(_0488_)
    );

    and_bi _1320_ (
        .a(new_Jinkela_wire_277),
        .b(new_Jinkela_wire_310),
        .c(_0489_)
    );

    and_ii _1321_ (
        .a(new_Jinkela_wire_2748),
        .b(new_Jinkela_wire_1133),
        .c(_0490_)
    );

    or_bb _1322_ (
        .a(_0490_),
        .b(new_Jinkela_wire_3092),
        .c(_0491_)
    );

    or_bb _1323_ (
        .a(new_Jinkela_wire_3309),
        .b(_0488_),
        .c(_0492_)
    );

    and_bi _1324_ (
        .a(new_Jinkela_wire_2771),
        .b(_0492_),
        .c(_0493_)
    );

    and_bi _1325_ (
        .a(_0480_),
        .b(_0493_),
        .c(_0494_)
    );

    and_bi _1326_ (
        .a(new_Jinkela_wire_1909),
        .b(_0494_),
        .c(_0495_)
    );

    or_bb _1327_ (
        .a(_0495_),
        .b(new_Jinkela_wire_1342),
        .c(_0496_)
    );

    and_bi _1328_ (
        .a(_0465_),
        .b(new_Jinkela_wire_1162),
        .c(_0497_)
    );

    inv _1329_ (
        .din(new_Jinkela_wire_3),
        .dout(_0498_)
    );

    and_bi _1330_ (
        .a(new_Jinkela_wire_2318),
        .b(new_Jinkela_wire_3162),
        .c(_0499_)
    );

    bfr new_Jinkela_buffer_1576 (
        .din(new_Jinkela_wire_2558),
        .dout(new_Jinkela_wire_2559)
    );

    bfr new_Jinkela_buffer_387 (
        .din(new_Jinkela_wire_719),
        .dout(new_Jinkela_wire_720)
    );

    bfr new_Jinkela_buffer_1557 (
        .din(new_Jinkela_wire_2527),
        .dout(new_Jinkela_wire_2528)
    );

    spl3L new_Jinkela_splitter_132 (
        .a(new_Jinkela_wire_738),
        .d(new_Jinkela_wire_739),
        .b(new_Jinkela_wire_740),
        .c(new_Jinkela_wire_741)
    );

    bfr new_Jinkela_buffer_1584 (
        .din(new_net_1475),
        .dout(new_Jinkela_wire_2588)
    );

    bfr new_Jinkela_buffer_388 (
        .din(new_Jinkela_wire_720),
        .dout(new_Jinkela_wire_721)
    );

    bfr new_Jinkela_buffer_1582 (
        .din(new_Jinkela_wire_2581),
        .dout(new_Jinkela_wire_2582)
    );

    bfr new_Jinkela_buffer_1558 (
        .din(new_Jinkela_wire_2528),
        .dout(new_Jinkela_wire_2529)
    );

    bfr new_Jinkela_buffer_398 (
        .din(new_Jinkela_wire_751),
        .dout(new_Jinkela_wire_752)
    );

    spl2 new_Jinkela_splitter_381 (
        .a(new_Jinkela_wire_2559),
        .b(new_Jinkela_wire_2560),
        .c(new_Jinkela_wire_2561)
    );

    spl2 new_Jinkela_splitter_135 (
        .a(new_Jinkela_wire_749),
        .b(new_Jinkela_wire_750),
        .c(new_Jinkela_wire_751)
    );

    spl2 new_Jinkela_splitter_127 (
        .a(new_Jinkela_wire_721),
        .b(new_Jinkela_wire_722),
        .c(new_Jinkela_wire_723)
    );

    bfr new_Jinkela_buffer_1559 (
        .din(new_Jinkela_wire_2529),
        .dout(new_Jinkela_wire_2530)
    );

    bfr new_Jinkela_buffer_389 (
        .din(new_Jinkela_wire_723),
        .dout(new_Jinkela_wire_724)
    );

    spl2 new_Jinkela_splitter_382 (
        .a(new_Jinkela_wire_2561),
        .b(new_Jinkela_wire_2562),
        .c(new_Jinkela_wire_2566)
    );

    bfr new_Jinkela_buffer_1560 (
        .din(new_Jinkela_wire_2530),
        .dout(new_Jinkela_wire_2531)
    );

    spl2 new_Jinkela_splitter_140 (
        .a(G37),
        .b(new_Jinkela_wire_777),
        .c(new_Jinkela_wire_778)
    );

    bfr new_Jinkela_buffer_394 (
        .din(new_Jinkela_wire_743),
        .dout(new_Jinkela_wire_744)
    );

    spl2 new_Jinkela_splitter_128 (
        .a(new_Jinkela_wire_724),
        .b(new_Jinkela_wire_725),
        .c(new_Jinkela_wire_726)
    );

    bfr new_Jinkela_buffer_1561 (
        .din(new_Jinkela_wire_2531),
        .dout(new_Jinkela_wire_2532)
    );

    spl2 new_Jinkela_splitter_129 (
        .a(new_Jinkela_wire_726),
        .b(new_Jinkela_wire_727),
        .c(new_Jinkela_wire_728)
    );

    spl4L new_Jinkela_splitter_384 (
        .a(new_Jinkela_wire_2566),
        .d(new_Jinkela_wire_2567),
        .e(new_Jinkela_wire_2568),
        .b(new_Jinkela_wire_2569),
        .c(new_Jinkela_wire_2570)
    );

    spl2 new_Jinkela_splitter_375 (
        .a(new_Jinkela_wire_2532),
        .b(new_Jinkela_wire_2533),
        .c(new_Jinkela_wire_2534)
    );

    bfr new_Jinkela_buffer_390 (
        .din(new_Jinkela_wire_728),
        .dout(new_Jinkela_wire_729)
    );

    bfr new_Jinkela_buffer_1562 (
        .din(new_Jinkela_wire_2534),
        .dout(new_Jinkela_wire_2535)
    );

    spl2 new_Jinkela_splitter_133 (
        .a(new_Jinkela_wire_741),
        .b(new_Jinkela_wire_742),
        .c(new_Jinkela_wire_743)
    );

    spl3L new_Jinkela_splitter_383 (
        .a(new_Jinkela_wire_2562),
        .d(new_Jinkela_wire_2563),
        .b(new_Jinkela_wire_2564),
        .c(new_Jinkela_wire_2565)
    );

    bfr new_Jinkela_buffer_402 (
        .din(new_Jinkela_wire_755),
        .dout(new_Jinkela_wire_756)
    );

    bfr new_Jinkela_buffer_395 (
        .din(new_Jinkela_wire_744),
        .dout(new_Jinkela_wire_745)
    );

    bfr new_Jinkela_buffer_391 (
        .din(new_Jinkela_wire_729),
        .dout(new_Jinkela_wire_730)
    );

    spl2 new_Jinkela_splitter_389 (
        .a(_0076_),
        .b(new_Jinkela_wire_2638),
        .c(new_Jinkela_wire_2639)
    );

    bfr new_Jinkela_buffer_1563 (
        .din(new_Jinkela_wire_2535),
        .dout(new_Jinkela_wire_2536)
    );

    bfr new_Jinkela_buffer_1633 (
        .din(_0389_),
        .dout(new_Jinkela_wire_2637)
    );

    bfr new_Jinkela_buffer_419 (
        .din(G49),
        .dout(new_Jinkela_wire_788)
    );

    bfr new_Jinkela_buffer_392 (
        .din(new_Jinkela_wire_730),
        .dout(new_Jinkela_wire_731)
    );

    spl2 new_Jinkela_splitter_376 (
        .a(new_Jinkela_wire_2536),
        .b(new_Jinkela_wire_2537),
        .c(new_Jinkela_wire_2538)
    );

    spl2 new_Jinkela_splitter_138 (
        .a(new_Jinkela_wire_770),
        .b(new_Jinkela_wire_771),
        .c(new_Jinkela_wire_772)
    );

    bfr new_Jinkela_buffer_1564 (
        .din(new_Jinkela_wire_2538),
        .dout(new_Jinkela_wire_2539)
    );

    spl2 new_Jinkela_splitter_134 (
        .a(new_Jinkela_wire_745),
        .b(new_Jinkela_wire_746),
        .c(new_Jinkela_wire_747)
    );

    bfr new_Jinkela_buffer_1585 (
        .din(new_Jinkela_wire_2588),
        .dout(new_Jinkela_wire_2589)
    );

    bfr new_Jinkela_buffer_403 (
        .din(new_Jinkela_wire_756),
        .dout(new_Jinkela_wire_757)
    );

    bfr new_Jinkela_buffer_1634 (
        .din(_0366_),
        .dout(new_Jinkela_wire_2640)
    );

    bfr new_Jinkela_buffer_399 (
        .din(new_Jinkela_wire_752),
        .dout(new_Jinkela_wire_753)
    );

    bfr new_Jinkela_buffer_1586 (
        .din(new_Jinkela_wire_2589),
        .dout(new_Jinkela_wire_2590)
    );

    bfr new_Jinkela_buffer_1565 (
        .din(new_Jinkela_wire_2539),
        .dout(new_Jinkela_wire_2540)
    );

    bfr new_Jinkela_buffer_400 (
        .din(new_Jinkela_wire_753),
        .dout(new_Jinkela_wire_754)
    );

    spl3L new_Jinkela_splitter_391 (
        .a(_0336_),
        .d(new_Jinkela_wire_2646),
        .b(new_Jinkela_wire_2647),
        .c(new_Jinkela_wire_2648)
    );

    bfr new_Jinkela_buffer_1566 (
        .din(new_Jinkela_wire_2540),
        .dout(new_Jinkela_wire_2541)
    );

    bfr new_Jinkela_buffer_404 (
        .din(new_Jinkela_wire_757),
        .dout(new_Jinkela_wire_758)
    );

    bfr new_Jinkela_buffer_1635 (
        .din(new_Jinkela_wire_2640),
        .dout(new_Jinkela_wire_2641)
    );

    bfr new_Jinkela_buffer_1587 (
        .din(new_Jinkela_wire_2590),
        .dout(new_Jinkela_wire_2591)
    );

    spl2 new_Jinkela_splitter_377 (
        .a(new_Jinkela_wire_2541),
        .b(new_Jinkela_wire_2542),
        .c(new_Jinkela_wire_2543)
    );

    bfr new_Jinkela_buffer_405 (
        .din(new_Jinkela_wire_758),
        .dout(new_Jinkela_wire_759)
    );

    bfr new_Jinkela_buffer_1567 (
        .din(new_Jinkela_wire_2543),
        .dout(new_Jinkela_wire_2544)
    );

    spl4L new_Jinkela_splitter_137 (
        .a(new_Jinkela_wire_766),
        .d(new_Jinkela_wire_767),
        .e(new_Jinkela_wire_768),
        .b(new_Jinkela_wire_769),
        .c(new_Jinkela_wire_770)
    );

    bfr new_Jinkela_buffer_406 (
        .din(new_Jinkela_wire_759),
        .dout(new_Jinkela_wire_760)
    );

    spl3L new_Jinkela_splitter_141 (
        .a(new_Jinkela_wire_778),
        .d(new_Jinkela_wire_779),
        .b(new_Jinkela_wire_780),
        .c(new_Jinkela_wire_781)
    );

    bfr new_Jinkela_buffer_1588 (
        .din(new_Jinkela_wire_2591),
        .dout(new_Jinkela_wire_2592)
    );

    spl2 new_Jinkela_splitter_378 (
        .a(new_Jinkela_wire_2544),
        .b(new_Jinkela_wire_2545),
        .c(new_Jinkela_wire_2546)
    );

    bfr new_Jinkela_buffer_407 (
        .din(new_Jinkela_wire_760),
        .dout(new_Jinkela_wire_761)
    );

    bfr new_Jinkela_buffer_1568 (
        .din(new_Jinkela_wire_2546),
        .dout(new_Jinkela_wire_2547)
    );

    bfr new_Jinkela_buffer_411 (
        .din(new_Jinkela_wire_772),
        .dout(new_Jinkela_wire_773)
    );

    bfr new_Jinkela_buffer_408 (
        .din(new_Jinkela_wire_761),
        .dout(new_Jinkela_wire_762)
    );

    spl2 new_Jinkela_splitter_390 (
        .a(_0793_),
        .b(new_Jinkela_wire_2644),
        .c(new_Jinkela_wire_2645)
    );

    bfr new_Jinkela_buffer_417 (
        .din(G45),
        .dout(new_Jinkela_wire_786)
    );

    bfr new_Jinkela_buffer_1589 (
        .din(new_Jinkela_wire_2592),
        .dout(new_Jinkela_wire_2593)
    );

    bfr new_Jinkela_buffer_1569 (
        .din(new_Jinkela_wire_2547),
        .dout(new_Jinkela_wire_2548)
    );

    bfr new_Jinkela_buffer_409 (
        .din(new_Jinkela_wire_762),
        .dout(new_Jinkela_wire_763)
    );

    bfr new_Jinkela_buffer_418 (
        .din(new_Jinkela_wire_786),
        .dout(new_Jinkela_wire_787)
    );

    bfr new_Jinkela_buffer_1638 (
        .din(_0435_),
        .dout(new_Jinkela_wire_2649)
    );

    spl2 new_Jinkela_splitter_379 (
        .a(new_Jinkela_wire_2548),
        .b(new_Jinkela_wire_2549),
        .c(new_Jinkela_wire_2550)
    );

    spl2 new_Jinkela_splitter_136 (
        .a(new_Jinkela_wire_763),
        .b(new_Jinkela_wire_764),
        .c(new_Jinkela_wire_765)
    );

    bfr new_Jinkela_buffer_422 (
        .din(G15),
        .dout(new_Jinkela_wire_791)
    );

    bfr new_Jinkela_buffer_1636 (
        .din(new_Jinkela_wire_2641),
        .dout(new_Jinkela_wire_2642)
    );

    bfr new_Jinkela_buffer_412 (
        .din(new_Jinkela_wire_773),
        .dout(new_Jinkela_wire_774)
    );

    bfr new_Jinkela_buffer_1590 (
        .din(new_Jinkela_wire_2593),
        .dout(new_Jinkela_wire_2594)
    );

    spl2 new_Jinkela_splitter_139 (
        .a(new_Jinkela_wire_774),
        .b(new_Jinkela_wire_775),
        .c(new_Jinkela_wire_776)
    );

    bfr new_Jinkela_buffer_1591 (
        .din(new_Jinkela_wire_2594),
        .dout(new_Jinkela_wire_2595)
    );

    bfr new_Jinkela_buffer_420 (
        .din(new_Jinkela_wire_788),
        .dout(new_Jinkela_wire_789)
    );

    bfr new_Jinkela_buffer_413 (
        .din(new_Jinkela_wire_781),
        .dout(new_Jinkela_wire_782)
    );

    bfr new_Jinkela_buffer_414 (
        .din(new_Jinkela_wire_782),
        .dout(new_Jinkela_wire_783)
    );

    bfr new_Jinkela_buffer_1592 (
        .din(new_Jinkela_wire_2595),
        .dout(new_Jinkela_wire_2596)
    );

    bfr new_Jinkela_buffer_415 (
        .din(new_Jinkela_wire_783),
        .dout(new_Jinkela_wire_784)
    );

    bfr new_Jinkela_buffer_1637 (
        .din(new_Jinkela_wire_2642),
        .dout(new_Jinkela_wire_2643)
    );

    bfr new_Jinkela_buffer_318 (
        .din(new_Jinkela_wire_606),
        .dout(new_Jinkela_wire_607)
    );

    bfr new_Jinkela_buffer_344 (
        .din(new_Jinkela_wire_637),
        .dout(new_Jinkela_wire_638)
    );

    bfr new_Jinkela_buffer_319 (
        .din(new_Jinkela_wire_607),
        .dout(new_Jinkela_wire_608)
    );

    bfr new_Jinkela_buffer_320 (
        .din(new_Jinkela_wire_608),
        .dout(new_Jinkela_wire_609)
    );

    spl2 new_Jinkela_splitter_118 (
        .a(G44),
        .b(new_Jinkela_wire_689),
        .c(new_Jinkela_wire_690)
    );

    bfr new_Jinkela_buffer_345 (
        .din(new_Jinkela_wire_638),
        .dout(new_Jinkela_wire_639)
    );

    bfr new_Jinkela_buffer_321 (
        .din(new_Jinkela_wire_609),
        .dout(new_Jinkela_wire_610)
    );

    bfr new_Jinkela_buffer_359 (
        .din(new_Jinkela_wire_660),
        .dout(new_Jinkela_wire_661)
    );

    bfr new_Jinkela_buffer_322 (
        .din(new_Jinkela_wire_610),
        .dout(new_Jinkela_wire_611)
    );

    spl2 new_Jinkela_splitter_112 (
        .a(new_Jinkela_wire_648),
        .b(new_Jinkela_wire_649),
        .c(new_Jinkela_wire_650)
    );

    bfr new_Jinkela_buffer_346 (
        .din(new_Jinkela_wire_639),
        .dout(new_Jinkela_wire_640)
    );

    bfr new_Jinkela_buffer_323 (
        .din(new_Jinkela_wire_611),
        .dout(new_Jinkela_wire_612)
    );

    spl2 new_Jinkela_splitter_116 (
        .a(new_Jinkela_wire_677),
        .b(new_Jinkela_wire_678),
        .c(new_Jinkela_wire_679)
    );

    bfr new_Jinkela_buffer_324 (
        .din(new_Jinkela_wire_612),
        .dout(new_Jinkela_wire_613)
    );

    bfr new_Jinkela_buffer_347 (
        .din(new_Jinkela_wire_640),
        .dout(new_Jinkela_wire_641)
    );

    bfr new_Jinkela_buffer_325 (
        .din(new_Jinkela_wire_613),
        .dout(new_Jinkela_wire_614)
    );

    bfr new_Jinkela_buffer_326 (
        .din(new_Jinkela_wire_614),
        .dout(new_Jinkela_wire_615)
    );

    bfr new_Jinkela_buffer_351 (
        .din(new_Jinkela_wire_650),
        .dout(new_Jinkela_wire_651)
    );

    bfr new_Jinkela_buffer_348 (
        .din(new_Jinkela_wire_641),
        .dout(new_Jinkela_wire_642)
    );

    bfr new_Jinkela_buffer_327 (
        .din(new_Jinkela_wire_615),
        .dout(new_Jinkela_wire_616)
    );

    bfr new_Jinkela_buffer_328 (
        .din(new_Jinkela_wire_616),
        .dout(new_Jinkela_wire_617)
    );

    bfr new_Jinkela_buffer_349 (
        .din(new_Jinkela_wire_642),
        .dout(new_Jinkela_wire_643)
    );

    bfr new_Jinkela_buffer_329 (
        .din(new_Jinkela_wire_617),
        .dout(new_Jinkela_wire_618)
    );

    bfr new_Jinkela_buffer_360 (
        .din(new_Jinkela_wire_661),
        .dout(new_Jinkela_wire_662)
    );

    bfr new_Jinkela_buffer_330 (
        .din(new_Jinkela_wire_618),
        .dout(new_Jinkela_wire_619)
    );

    bfr new_Jinkela_buffer_350 (
        .din(new_Jinkela_wire_643),
        .dout(new_Jinkela_wire_644)
    );

    bfr new_Jinkela_buffer_331 (
        .din(new_Jinkela_wire_619),
        .dout(new_Jinkela_wire_620)
    );

    bfr new_Jinkela_buffer_370 (
        .din(new_Jinkela_wire_679),
        .dout(new_Jinkela_wire_680)
    );

    bfr new_Jinkela_buffer_332 (
        .din(new_Jinkela_wire_620),
        .dout(new_Jinkela_wire_621)
    );

    bfr new_Jinkela_buffer_352 (
        .din(new_Jinkela_wire_651),
        .dout(new_Jinkela_wire_652)
    );

    bfr new_Jinkela_buffer_333 (
        .din(new_Jinkela_wire_621),
        .dout(new_Jinkela_wire_622)
    );

    bfr new_Jinkela_buffer_361 (
        .din(new_Jinkela_wire_662),
        .dout(new_Jinkela_wire_663)
    );

    bfr new_Jinkela_buffer_334 (
        .din(new_Jinkela_wire_622),
        .dout(new_Jinkela_wire_623)
    );

    bfr new_Jinkela_buffer_353 (
        .din(new_Jinkela_wire_652),
        .dout(new_Jinkela_wire_653)
    );

    bfr new_Jinkela_buffer_335 (
        .din(new_Jinkela_wire_623),
        .dout(new_Jinkela_wire_624)
    );

    bfr new_Jinkela_buffer_336 (
        .din(new_Jinkela_wire_624),
        .dout(new_Jinkela_wire_625)
    );

    bfr new_Jinkela_buffer_362 (
        .din(new_Jinkela_wire_663),
        .dout(new_Jinkela_wire_664)
    );

    bfr new_Jinkela_buffer_354 (
        .din(new_Jinkela_wire_653),
        .dout(new_Jinkela_wire_654)
    );

    bfr new_Jinkela_buffer_337 (
        .din(new_Jinkela_wire_625),
        .dout(new_Jinkela_wire_626)
    );

    spl2 new_Jinkela_splitter_120 (
        .a(G12),
        .b(new_Jinkela_wire_701),
        .c(new_Jinkela_wire_704)
    );

    bfr new_Jinkela_buffer_355 (
        .din(new_Jinkela_wire_654),
        .dout(new_Jinkela_wire_655)
    );

    bfr new_Jinkela_buffer_377 (
        .din(new_Jinkela_wire_690),
        .dout(new_Jinkela_wire_691)
    );

    or_bb _0953_ (
        .a(_0124_),
        .b(new_Jinkela_wire_1727),
        .c(_0125_)
    );

    or_bi _0954_ (
        .a(_0125_),
        .b(_0119_),
        .c(_0126_)
    );

    or_bi _0955_ (
        .a(new_Jinkela_wire_3219),
        .b(new_Jinkela_wire_775),
        .c(_0127_)
    );

    and_bi _0956_ (
        .a(new_Jinkela_wire_176),
        .b(new_Jinkela_wire_3028),
        .c(_0128_)
    );

    or_bb _0957_ (
        .a(new_Jinkela_wire_439),
        .b(new_Jinkela_wire_222),
        .c(_0129_)
    );

    and_bi _0958_ (
        .a(new_Jinkela_wire_437),
        .b(new_Jinkela_wire_309),
        .c(_0130_)
    );

    and_bi _0959_ (
        .a(_0129_),
        .b(_0130_),
        .c(_0131_)
    );

    or_bb _0960_ (
        .a(new_Jinkela_wire_1179),
        .b(_0128_),
        .c(_0132_)
    );

    and_bi _0961_ (
        .a(new_Jinkela_wire_2065),
        .b(_0132_),
        .c(_0133_)
    );

    and_bi _0962_ (
        .a(new_Jinkela_wire_1048),
        .b(_0133_),
        .c(_0134_)
    );

    or_bb _0963_ (
        .a(new_Jinkela_wire_3043),
        .b(new_Jinkela_wire_839),
        .c(_0135_)
    );

    and_bi _0964_ (
        .a(new_Jinkela_wire_2568),
        .b(new_Jinkela_wire_2882),
        .c(_0136_)
    );

    or_bb _0965_ (
        .a(_0136_),
        .b(new_Jinkela_wire_1266),
        .c(_0137_)
    );

    or_bb _0966_ (
        .a(new_Jinkela_wire_2881),
        .b(new_Jinkela_wire_3066),
        .c(_0138_)
    );

    and_bi _0967_ (
        .a(new_Jinkela_wire_1265),
        .b(_0138_),
        .c(_0139_)
    );

    or_bi _0968_ (
        .a(new_Jinkela_wire_2878),
        .b(new_Jinkela_wire_2322),
        .c(_0140_)
    );

    inv _0969_ (
        .din(new_Jinkela_wire_3307),
        .dout(_0141_)
    );

    and_bi _0970_ (
        .a(new_Jinkela_wire_2874),
        .b(new_Jinkela_wire_3192),
        .c(_0142_)
    );

    or_bb _0971_ (
        .a(new_Jinkela_wire_934),
        .b(new_Jinkela_wire_208),
        .c(_0143_)
    );

    or_bb _0972_ (
        .a(new_Jinkela_wire_1282),
        .b(new_Jinkela_wire_1687),
        .c(_0144_)
    );

    and_bi _0973_ (
        .a(new_Jinkela_wire_747),
        .b(new_Jinkela_wire_3329),
        .c(_0145_)
    );

    and_bi _0974_ (
        .a(new_Jinkela_wire_3132),
        .b(_0145_),
        .c(_0146_)
    );

    and_bi _0975_ (
        .a(new_Jinkela_wire_3317),
        .b(_0146_),
        .c(_0147_)
    );

    and_bi _0976_ (
        .a(new_Jinkela_wire_2170),
        .b(new_Jinkela_wire_1944),
        .c(_0148_)
    );

    or_bb _0977_ (
        .a(_0148_),
        .b(_0147_),
        .c(_0149_)
    );

    and_bi _0978_ (
        .a(_0143_),
        .b(new_Jinkela_wire_2002),
        .c(_0150_)
    );

    inv _0979_ (
        .din(new_Jinkela_wire_305),
        .dout(_0151_)
    );

    or_bb _0980_ (
        .a(new_Jinkela_wire_3221),
        .b(new_Jinkela_wire_990),
        .c(_0152_)
    );

    and_bi _0981_ (
        .a(new_Jinkela_wire_44),
        .b(new_Jinkela_wire_3032),
        .c(_0153_)
    );

    or_bb _0982_ (
        .a(new_Jinkela_wire_443),
        .b(new_Jinkela_wire_712),
        .c(_0154_)
    );

    and_bi _0983_ (
        .a(new_Jinkela_wire_434),
        .b(new_Jinkela_wire_173),
        .c(_0155_)
    );

    and_bi _0984_ (
        .a(new_Jinkela_wire_2335),
        .b(new_Jinkela_wire_1403),
        .c(_0156_)
    );

    or_bb _0985_ (
        .a(_0156_),
        .b(_0153_),
        .c(_0157_)
    );

    and_bi _0986_ (
        .a(new_Jinkela_wire_2114),
        .b(_0157_),
        .c(_0158_)
    );

    and_bi _0987_ (
        .a(new_Jinkela_wire_1049),
        .b(_0158_),
        .c(_0159_)
    );

    or_bb _0988_ (
        .a(new_Jinkela_wire_1163),
        .b(new_Jinkela_wire_840),
        .c(_0160_)
    );

    and_bi _0989_ (
        .a(new_Jinkela_wire_2569),
        .b(new_Jinkela_wire_3255),
        .c(_0161_)
    );

    and_bi _0990_ (
        .a(new_Jinkela_wire_2447),
        .b(_0161_),
        .c(_0162_)
    );

    and_ii _0991_ (
        .a(new_Jinkela_wire_3254),
        .b(new_Jinkela_wire_3065),
        .c(_0163_)
    );

    and_bi _0992_ (
        .a(_0163_),
        .b(new_Jinkela_wire_2449),
        .c(_0164_)
    );

    or_bb _0993_ (
        .a(new_Jinkela_wire_3014),
        .b(new_Jinkela_wire_836),
        .c(_0165_)
    );

    or_bb _0994_ (
        .a(new_Jinkela_wire_1980),
        .b(new_Jinkela_wire_1628),
        .c(_0166_)
    );

    bfr new_Jinkela_buffer_304 (
        .din(new_Jinkela_wire_557),
        .dout(new_Jinkela_wire_558)
    );

    bfr new_Jinkela_buffer_1253 (
        .din(new_Jinkela_wire_2054),
        .dout(new_Jinkela_wire_2055)
    );

    bfr new_Jinkela_buffer_293 (
        .din(new_Jinkela_wire_544),
        .dout(new_Jinkela_wire_545)
    );

    spl3L new_Jinkela_splitter_314 (
        .a(new_Jinkela_wire_2071),
        .d(new_Jinkela_wire_2072),
        .b(new_Jinkela_wire_2073),
        .c(new_Jinkela_wire_2074)
    );

    spl3L new_Jinkela_splitter_104 (
        .a(new_Jinkela_wire_587),
        .d(new_Jinkela_wire_588),
        .b(new_Jinkela_wire_589),
        .c(new_Jinkela_wire_590)
    );

    bfr new_Jinkela_buffer_1261 (
        .din(new_Jinkela_wire_2068),
        .dout(new_Jinkela_wire_2069)
    );

    bfr new_Jinkela_buffer_1254 (
        .din(new_Jinkela_wire_2055),
        .dout(new_Jinkela_wire_2056)
    );

    bfr new_Jinkela_buffer_294 (
        .din(new_Jinkela_wire_545),
        .dout(new_Jinkela_wire_546)
    );

    spl2 new_Jinkela_splitter_103 (
        .a(G1),
        .b(new_Jinkela_wire_587),
        .c(new_Jinkela_wire_591)
    );

    bfr new_Jinkela_buffer_308 (
        .din(new_Jinkela_wire_563),
        .dout(new_Jinkela_wire_564)
    );

    bfr new_Jinkela_buffer_1255 (
        .din(new_Jinkela_wire_2056),
        .dout(new_Jinkela_wire_2057)
    );

    bfr new_Jinkela_buffer_295 (
        .din(new_Jinkela_wire_546),
        .dout(new_Jinkela_wire_547)
    );

    bfr new_Jinkela_buffer_1272 (
        .din(new_Jinkela_wire_2090),
        .dout(new_Jinkela_wire_2091)
    );

    bfr new_Jinkela_buffer_305 (
        .din(new_Jinkela_wire_558),
        .dout(new_Jinkela_wire_559)
    );

    bfr new_Jinkela_buffer_1262 (
        .din(new_Jinkela_wire_2069),
        .dout(new_Jinkela_wire_2070)
    );

    bfr new_Jinkela_buffer_1256 (
        .din(new_Jinkela_wire_2057),
        .dout(new_Jinkela_wire_2058)
    );

    bfr new_Jinkela_buffer_296 (
        .din(new_Jinkela_wire_547),
        .dout(new_Jinkela_wire_548)
    );

    bfr new_Jinkela_buffer_1271 (
        .din(_0356_),
        .dout(new_Jinkela_wire_2090)
    );

    bfr new_Jinkela_buffer_1257 (
        .din(new_Jinkela_wire_2058),
        .dout(new_Jinkela_wire_2059)
    );

    bfr new_Jinkela_buffer_297 (
        .din(new_Jinkela_wire_548),
        .dout(new_Jinkela_wire_549)
    );

    spl2 new_Jinkela_splitter_317 (
        .a(_0065_),
        .b(new_Jinkela_wire_2086),
        .c(new_Jinkela_wire_2087)
    );

    bfr new_Jinkela_buffer_306 (
        .din(new_Jinkela_wire_559),
        .dout(new_Jinkela_wire_560)
    );

    bfr new_Jinkela_buffer_1264 (
        .din(new_Jinkela_wire_2074),
        .dout(new_Jinkela_wire_2075)
    );

    bfr new_Jinkela_buffer_1258 (
        .din(new_Jinkela_wire_2059),
        .dout(new_Jinkela_wire_2060)
    );

    bfr new_Jinkela_buffer_298 (
        .din(new_Jinkela_wire_549),
        .dout(new_Jinkela_wire_550)
    );

    bfr new_Jinkela_buffer_1266 (
        .din(new_Jinkela_wire_2078),
        .dout(new_Jinkela_wire_2079)
    );

    spl2 new_Jinkela_splitter_96 (
        .a(new_Jinkela_wire_564),
        .b(new_Jinkela_wire_565),
        .c(new_Jinkela_wire_566)
    );

    spl2 new_Jinkela_splitter_318 (
        .a(new_Jinkela_wire_2087),
        .b(new_Jinkela_wire_2088),
        .c(new_Jinkela_wire_2089)
    );

    bfr new_Jinkela_buffer_299 (
        .din(new_Jinkela_wire_550),
        .dout(new_Jinkela_wire_551)
    );

    bfr new_Jinkela_buffer_1265 (
        .din(new_Jinkela_wire_2075),
        .dout(new_Jinkela_wire_2076)
    );

    spl4L new_Jinkela_splitter_105 (
        .a(new_Jinkela_wire_591),
        .d(new_Jinkela_wire_592),
        .e(new_Jinkela_wire_593),
        .b(new_Jinkela_wire_594),
        .c(new_Jinkela_wire_596)
    );

    bfr new_Jinkela_buffer_300 (
        .din(new_Jinkela_wire_551),
        .dout(new_Jinkela_wire_552)
    );

    bfr new_Jinkela_buffer_1295 (
        .din(_0452_),
        .dout(new_Jinkela_wire_2118)
    );

    bfr new_Jinkela_buffer_1267 (
        .din(new_Jinkela_wire_2079),
        .dout(new_Jinkela_wire_2080)
    );

    spl2 new_Jinkela_splitter_111 (
        .a(new_Jinkela_wire_646),
        .b(new_Jinkela_wire_647),
        .c(new_Jinkela_wire_648)
    );

    bfr new_Jinkela_buffer_1287 (
        .din(_0733_),
        .dout(new_Jinkela_wire_2110)
    );

    bfr new_Jinkela_buffer_309 (
        .din(new_Jinkela_wire_567),
        .dout(new_Jinkela_wire_568)
    );

    bfr new_Jinkela_buffer_1268 (
        .din(new_Jinkela_wire_2080),
        .dout(new_Jinkela_wire_2081)
    );

    bfr new_Jinkela_buffer_1288 (
        .din(new_Jinkela_wire_2110),
        .dout(new_Jinkela_wire_2111)
    );

    spl4L new_Jinkela_splitter_99 (
        .a(new_Jinkela_wire_573),
        .d(new_Jinkela_wire_574),
        .e(new_Jinkela_wire_575),
        .b(new_Jinkela_wire_576),
        .c(new_Jinkela_wire_577)
    );

    bfr new_Jinkela_buffer_1273 (
        .din(new_Jinkela_wire_2091),
        .dout(new_Jinkela_wire_2092)
    );

    spl2 new_Jinkela_splitter_100 (
        .a(new_Jinkela_wire_577),
        .b(new_Jinkela_wire_578),
        .c(new_Jinkela_wire_579)
    );

    bfr new_Jinkela_buffer_1269 (
        .din(new_Jinkela_wire_2081),
        .dout(new_Jinkela_wire_2082)
    );

    bfr new_Jinkela_buffer_1270 (
        .din(new_Jinkela_wire_2082),
        .dout(new_Jinkela_wire_2083)
    );

    bfr new_Jinkela_buffer_310 (
        .din(new_Jinkela_wire_579),
        .dout(new_Jinkela_wire_580)
    );

    bfr new_Jinkela_buffer_313 (
        .din(new_Jinkela_wire_594),
        .dout(new_Jinkela_wire_595)
    );

    spl2 new_Jinkela_splitter_108 (
        .a(G6),
        .b(new_Jinkela_wire_633),
        .c(new_Jinkela_wire_634)
    );

    spl2 new_Jinkela_splitter_316 (
        .a(new_Jinkela_wire_2083),
        .b(new_Jinkela_wire_2084),
        .c(new_Jinkela_wire_2085)
    );

    spl4L new_Jinkela_splitter_106 (
        .a(new_Jinkela_wire_596),
        .d(new_Jinkela_wire_597),
        .e(new_Jinkela_wire_598),
        .b(new_Jinkela_wire_599),
        .c(new_Jinkela_wire_600)
    );

    bfr new_Jinkela_buffer_340 (
        .din(new_Jinkela_wire_628),
        .dout(new_Jinkela_wire_629)
    );

    bfr new_Jinkela_buffer_311 (
        .din(new_Jinkela_wire_580),
        .dout(new_Jinkela_wire_581)
    );

    bfr new_Jinkela_buffer_1292 (
        .din(_0650_),
        .dout(new_Jinkela_wire_2115)
    );

    bfr new_Jinkela_buffer_1274 (
        .din(new_Jinkela_wire_2092),
        .dout(new_Jinkela_wire_2093)
    );

    bfr new_Jinkela_buffer_1289 (
        .din(new_Jinkela_wire_2111),
        .dout(new_Jinkela_wire_2112)
    );

    spl2 new_Jinkela_splitter_107 (
        .a(new_Jinkela_wire_600),
        .b(new_Jinkela_wire_601),
        .c(new_Jinkela_wire_602)
    );

    bfr new_Jinkela_buffer_1275 (
        .din(new_Jinkela_wire_2093),
        .dout(new_Jinkela_wire_2094)
    );

    spl2 new_Jinkela_splitter_101 (
        .a(new_Jinkela_wire_581),
        .b(new_Jinkela_wire_582),
        .c(new_Jinkela_wire_583)
    );

    bfr new_Jinkela_buffer_312 (
        .din(new_Jinkela_wire_583),
        .dout(new_Jinkela_wire_584)
    );

    bfr new_Jinkela_buffer_339 (
        .din(new_Jinkela_wire_627),
        .dout(new_Jinkela_wire_628)
    );

    bfr new_Jinkela_buffer_1290 (
        .din(new_Jinkela_wire_2112),
        .dout(new_Jinkela_wire_2113)
    );

    bfr new_Jinkela_buffer_338 (
        .din(G28),
        .dout(new_Jinkela_wire_627)
    );

    bfr new_Jinkela_buffer_1276 (
        .din(new_Jinkela_wire_2094),
        .dout(new_Jinkela_wire_2095)
    );

    spl2 new_Jinkela_splitter_102 (
        .a(new_Jinkela_wire_584),
        .b(new_Jinkela_wire_585),
        .c(new_Jinkela_wire_586)
    );

    bfr new_Jinkela_buffer_1291 (
        .din(_0152_),
        .dout(new_Jinkela_wire_2114)
    );

    bfr new_Jinkela_buffer_1277 (
        .din(new_Jinkela_wire_2095),
        .dout(new_Jinkela_wire_2096)
    );

    spl2 new_Jinkela_splitter_110 (
        .a(G24),
        .b(new_Jinkela_wire_645),
        .c(new_Jinkela_wire_646)
    );

    spl3L new_Jinkela_splitter_109 (
        .a(new_Jinkela_wire_634),
        .d(new_Jinkela_wire_635),
        .b(new_Jinkela_wire_636),
        .c(new_Jinkela_wire_637)
    );

    bfr new_Jinkela_buffer_1293 (
        .din(new_Jinkela_wire_2115),
        .dout(new_Jinkela_wire_2116)
    );

    bfr new_Jinkela_buffer_314 (
        .din(new_Jinkela_wire_602),
        .dout(new_Jinkela_wire_603)
    );

    bfr new_Jinkela_buffer_1278 (
        .din(new_Jinkela_wire_2096),
        .dout(new_Jinkela_wire_2097)
    );

    bfr new_Jinkela_buffer_341 (
        .din(new_Jinkela_wire_629),
        .dout(new_Jinkela_wire_630)
    );

    bfr new_Jinkela_buffer_1297 (
        .din(new_net_1477),
        .dout(new_Jinkela_wire_2120)
    );

    bfr new_Jinkela_buffer_315 (
        .din(new_Jinkela_wire_603),
        .dout(new_Jinkela_wire_604)
    );

    bfr new_Jinkela_buffer_1279 (
        .din(new_Jinkela_wire_2097),
        .dout(new_Jinkela_wire_2098)
    );

    bfr new_Jinkela_buffer_358 (
        .din(G20),
        .dout(new_Jinkela_wire_660)
    );

    bfr new_Jinkela_buffer_342 (
        .din(new_Jinkela_wire_630),
        .dout(new_Jinkela_wire_631)
    );

    bfr new_Jinkela_buffer_1294 (
        .din(new_Jinkela_wire_2116),
        .dout(new_Jinkela_wire_2117)
    );

    bfr new_Jinkela_buffer_316 (
        .din(new_Jinkela_wire_604),
        .dout(new_Jinkela_wire_605)
    );

    bfr new_Jinkela_buffer_1280 (
        .din(new_Jinkela_wire_2098),
        .dout(new_Jinkela_wire_2099)
    );

    bfr new_Jinkela_buffer_1296 (
        .din(new_Jinkela_wire_2118),
        .dout(new_Jinkela_wire_2119)
    );

    bfr new_Jinkela_buffer_317 (
        .din(new_Jinkela_wire_605),
        .dout(new_Jinkela_wire_606)
    );

    bfr new_Jinkela_buffer_1281 (
        .din(new_Jinkela_wire_2099),
        .dout(new_Jinkela_wire_2100)
    );

    bfr new_Jinkela_buffer_369 (
        .din(G43),
        .dout(new_Jinkela_wire_677)
    );

    bfr new_Jinkela_buffer_343 (
        .din(new_Jinkela_wire_631),
        .dout(new_Jinkela_wire_632)
    );

    spl2 new_Jinkela_splitter_320 (
        .a(_0071_),
        .b(new_Jinkela_wire_2165),
        .c(new_Jinkela_wire_2166)
    );

    bfr new_Jinkela_buffer_1593 (
        .din(new_Jinkela_wire_2596),
        .dout(new_Jinkela_wire_2597)
    );

    bfr new_Jinkela_buffer_1639 (
        .din(new_Jinkela_wire_2653),
        .dout(new_Jinkela_wire_2654)
    );

    spl3L new_Jinkela_splitter_393 (
        .a(new_net_5),
        .d(new_Jinkela_wire_2656),
        .b(new_Jinkela_wire_2657),
        .c(new_Jinkela_wire_2658)
    );

    bfr new_Jinkela_buffer_1594 (
        .din(new_Jinkela_wire_2597),
        .dout(new_Jinkela_wire_2598)
    );

    bfr new_Jinkela_buffer_1641 (
        .din(new_Jinkela_wire_2658),
        .dout(new_Jinkela_wire_2659)
    );

    bfr new_Jinkela_buffer_1595 (
        .din(new_Jinkela_wire_2598),
        .dout(new_Jinkela_wire_2599)
    );

    spl4L new_Jinkela_splitter_392 (
        .a(_0250_),
        .d(new_Jinkela_wire_2650),
        .e(new_Jinkela_wire_2651),
        .b(new_Jinkela_wire_2652),
        .c(new_Jinkela_wire_2653)
    );

    bfr new_Jinkela_buffer_1596 (
        .din(new_Jinkela_wire_2599),
        .dout(new_Jinkela_wire_2600)
    );

    bfr new_Jinkela_buffer_1657 (
        .din(new_net_1471),
        .dout(new_Jinkela_wire_2675)
    );

    bfr new_Jinkela_buffer_1597 (
        .din(new_Jinkela_wire_2600),
        .dout(new_Jinkela_wire_2601)
    );

    bfr new_Jinkela_buffer_1687 (
        .din(_0499_),
        .dout(new_Jinkela_wire_2705)
    );

    bfr new_Jinkela_buffer_1640 (
        .din(new_Jinkela_wire_2654),
        .dout(new_Jinkela_wire_2655)
    );

    bfr new_Jinkela_buffer_1598 (
        .din(new_Jinkela_wire_2601),
        .dout(new_Jinkela_wire_2602)
    );

    bfr new_Jinkela_buffer_1599 (
        .din(new_Jinkela_wire_2602),
        .dout(new_Jinkela_wire_2603)
    );

    bfr new_Jinkela_buffer_1658 (
        .din(new_Jinkela_wire_2675),
        .dout(new_Jinkela_wire_2676)
    );

    spl3L new_Jinkela_splitter_395 (
        .a(_0348_),
        .d(new_Jinkela_wire_2709),
        .b(new_Jinkela_wire_2710),
        .c(new_Jinkela_wire_2711)
    );

    bfr new_Jinkela_buffer_1600 (
        .din(new_Jinkela_wire_2603),
        .dout(new_Jinkela_wire_2604)
    );

    bfr new_Jinkela_buffer_1642 (
        .din(new_Jinkela_wire_2659),
        .dout(new_Jinkela_wire_2660)
    );

    bfr new_Jinkela_buffer_1601 (
        .din(new_Jinkela_wire_2604),
        .dout(new_Jinkela_wire_2605)
    );

    bfr new_Jinkela_buffer_1602 (
        .din(new_Jinkela_wire_2605),
        .dout(new_Jinkela_wire_2606)
    );

    bfr new_Jinkela_buffer_1688 (
        .din(new_Jinkela_wire_2705),
        .dout(new_Jinkela_wire_2706)
    );

    bfr new_Jinkela_buffer_1643 (
        .din(new_Jinkela_wire_2660),
        .dout(new_Jinkela_wire_2661)
    );

    bfr new_Jinkela_buffer_1603 (
        .din(new_Jinkela_wire_2606),
        .dout(new_Jinkela_wire_2607)
    );

    bfr new_Jinkela_buffer_1689 (
        .din(_0455_),
        .dout(new_Jinkela_wire_2712)
    );

    bfr new_Jinkela_buffer_1604 (
        .din(new_Jinkela_wire_2607),
        .dout(new_Jinkela_wire_2608)
    );

    bfr new_Jinkela_buffer_1659 (
        .din(new_Jinkela_wire_2676),
        .dout(new_Jinkela_wire_2677)
    );

    bfr new_Jinkela_buffer_1644 (
        .din(new_Jinkela_wire_2661),
        .dout(new_Jinkela_wire_2662)
    );

    bfr new_Jinkela_buffer_1605 (
        .din(new_Jinkela_wire_2608),
        .dout(new_Jinkela_wire_2609)
    );

    bfr new_Jinkela_buffer_1606 (
        .din(new_Jinkela_wire_2609),
        .dout(new_Jinkela_wire_2610)
    );

    bfr new_Jinkela_buffer_1645 (
        .din(new_Jinkela_wire_2662),
        .dout(new_Jinkela_wire_2663)
    );

    bfr new_Jinkela_buffer_1607 (
        .din(new_Jinkela_wire_2610),
        .dout(new_Jinkela_wire_2611)
    );

    bfr new_Jinkela_buffer_1608 (
        .din(new_Jinkela_wire_2611),
        .dout(new_Jinkela_wire_2612)
    );

    bfr new_Jinkela_buffer_1660 (
        .din(new_Jinkela_wire_2677),
        .dout(new_Jinkela_wire_2678)
    );

    bfr new_Jinkela_buffer_1646 (
        .din(new_Jinkela_wire_2663),
        .dout(new_Jinkela_wire_2664)
    );

    bfr new_Jinkela_buffer_1609 (
        .din(new_Jinkela_wire_2612),
        .dout(new_Jinkela_wire_2613)
    );

    bfr new_Jinkela_buffer_1610 (
        .din(new_Jinkela_wire_2613),
        .dout(new_Jinkela_wire_2614)
    );

    bfr new_Jinkela_buffer_1647 (
        .din(new_Jinkela_wire_2664),
        .dout(new_Jinkela_wire_2665)
    );

    bfr new_Jinkela_buffer_1611 (
        .din(new_Jinkela_wire_2614),
        .dout(new_Jinkela_wire_2615)
    );

    bfr new_Jinkela_buffer_1612 (
        .din(new_Jinkela_wire_2615),
        .dout(new_Jinkela_wire_2616)
    );

    bfr new_Jinkela_buffer_1661 (
        .din(new_Jinkela_wire_2678),
        .dout(new_Jinkela_wire_2679)
    );

    bfr new_Jinkela_buffer_1648 (
        .din(new_Jinkela_wire_2665),
        .dout(new_Jinkela_wire_2666)
    );

    bfr new_Jinkela_buffer_1613 (
        .din(new_Jinkela_wire_2616),
        .dout(new_Jinkela_wire_2617)
    );

    bfr new_Jinkela_buffer_1282 (
        .din(new_Jinkela_wire_2100),
        .dout(new_Jinkela_wire_2101)
    );

    spl4L new_Jinkela_splitter_321 (
        .a(_0052_),
        .d(new_Jinkela_wire_2167),
        .e(new_Jinkela_wire_2168),
        .b(new_Jinkela_wire_2169),
        .c(new_Jinkela_wire_2170)
    );

    bfr new_Jinkela_buffer_1298 (
        .din(new_Jinkela_wire_2120),
        .dout(new_Jinkela_wire_2121)
    );

    bfr new_Jinkela_buffer_1283 (
        .din(new_Jinkela_wire_2101),
        .dout(new_Jinkela_wire_2102)
    );

    bfr new_Jinkela_buffer_1284 (
        .din(new_Jinkela_wire_2102),
        .dout(new_Jinkela_wire_2103)
    );

    bfr new_Jinkela_buffer_1345 (
        .din(_0237_),
        .dout(new_Jinkela_wire_2183)
    );

    bfr new_Jinkela_buffer_1299 (
        .din(new_Jinkela_wire_2121),
        .dout(new_Jinkela_wire_2122)
    );

    bfr new_Jinkela_buffer_1285 (
        .din(new_Jinkela_wire_2103),
        .dout(new_Jinkela_wire_2104)
    );

    bfr new_Jinkela_buffer_1286 (
        .din(new_Jinkela_wire_2104),
        .dout(new_Jinkela_wire_2105)
    );

    spl3L new_Jinkela_splitter_322 (
        .a(_0212_),
        .d(new_Jinkela_wire_2171),
        .b(new_Jinkela_wire_2172),
        .c(new_Jinkela_wire_2173)
    );

    bfr new_Jinkela_buffer_1300 (
        .din(new_Jinkela_wire_2122),
        .dout(new_Jinkela_wire_2123)
    );

    spl4L new_Jinkela_splitter_319 (
        .a(new_Jinkela_wire_2105),
        .d(new_Jinkela_wire_2106),
        .e(new_Jinkela_wire_2107),
        .b(new_Jinkela_wire_2108),
        .c(new_Jinkela_wire_2109)
    );

    bfr new_Jinkela_buffer_1346 (
        .din(new_net_1473),
        .dout(new_Jinkela_wire_2184)
    );

    bfr new_Jinkela_buffer_1301 (
        .din(new_Jinkela_wire_2123),
        .dout(new_Jinkela_wire_2124)
    );

    spl4L new_Jinkela_splitter_324 (
        .a(_0213_),
        .d(new_Jinkela_wire_2176),
        .e(new_Jinkela_wire_2177),
        .b(new_Jinkela_wire_2178),
        .c(new_Jinkela_wire_2179)
    );

    spl2 new_Jinkela_splitter_323 (
        .a(_0430_),
        .b(new_Jinkela_wire_2174),
        .c(new_Jinkela_wire_2175)
    );

    bfr new_Jinkela_buffer_1302 (
        .din(new_Jinkela_wire_2124),
        .dout(new_Jinkela_wire_2125)
    );

    bfr new_Jinkela_buffer_1303 (
        .din(new_Jinkela_wire_2125),
        .dout(new_Jinkela_wire_2126)
    );

    bfr new_Jinkela_buffer_1343 (
        .din(new_Jinkela_wire_2180),
        .dout(new_Jinkela_wire_2181)
    );

    bfr new_Jinkela_buffer_1304 (
        .din(new_Jinkela_wire_2126),
        .dout(new_Jinkela_wire_2127)
    );

    bfr new_Jinkela_buffer_1342 (
        .din(new_Jinkela_wire_2179),
        .dout(new_Jinkela_wire_2180)
    );

    bfr new_Jinkela_buffer_1305 (
        .din(new_Jinkela_wire_2127),
        .dout(new_Jinkela_wire_2128)
    );

    bfr new_Jinkela_buffer_1350 (
        .din(_0198_),
        .dout(new_Jinkela_wire_2188)
    );

    bfr new_Jinkela_buffer_1306 (
        .din(new_Jinkela_wire_2128),
        .dout(new_Jinkela_wire_2129)
    );

    bfr new_Jinkela_buffer_1307 (
        .din(new_Jinkela_wire_2129),
        .dout(new_Jinkela_wire_2130)
    );

    bfr new_Jinkela_buffer_1347 (
        .din(new_Jinkela_wire_2184),
        .dout(new_Jinkela_wire_2185)
    );

    bfr new_Jinkela_buffer_1344 (
        .din(new_Jinkela_wire_2181),
        .dout(new_Jinkela_wire_2182)
    );

    bfr new_Jinkela_buffer_1308 (
        .din(new_Jinkela_wire_2130),
        .dout(new_Jinkela_wire_2131)
    );

    bfr new_Jinkela_buffer_1309 (
        .din(new_Jinkela_wire_2131),
        .dout(new_Jinkela_wire_2132)
    );

    spl2 new_Jinkela_splitter_325 (
        .a(_0286_),
        .b(new_Jinkela_wire_2190),
        .c(new_Jinkela_wire_2191)
    );

    bfr new_Jinkela_buffer_1366 (
        .din(_0193_),
        .dout(new_Jinkela_wire_2208)
    );

    bfr new_Jinkela_buffer_1310 (
        .din(new_Jinkela_wire_2132),
        .dout(new_Jinkela_wire_2133)
    );

    bfr new_Jinkela_buffer_1348 (
        .din(new_Jinkela_wire_2185),
        .dout(new_Jinkela_wire_2186)
    );

    bfr new_Jinkela_buffer_1311 (
        .din(new_Jinkela_wire_2133),
        .dout(new_Jinkela_wire_2134)
    );

    bfr new_Jinkela_buffer_1351 (
        .din(new_Jinkela_wire_2188),
        .dout(new_Jinkela_wire_2189)
    );

    bfr new_Jinkela_buffer_1312 (
        .din(new_Jinkela_wire_2134),
        .dout(new_Jinkela_wire_2135)
    );

    bfr new_Jinkela_buffer_1349 (
        .din(new_Jinkela_wire_2186),
        .dout(new_Jinkela_wire_2187)
    );

    bfr new_Jinkela_buffer_1313 (
        .din(new_Jinkela_wire_2135),
        .dout(new_Jinkela_wire_2136)
    );

    bfr new_Jinkela_buffer_1314 (
        .din(new_Jinkela_wire_2136),
        .dout(new_Jinkela_wire_2137)
    );

    bfr new_Jinkela_buffer_1368 (
        .din(_0210_),
        .dout(new_Jinkela_wire_2210)
    );

    bfr new_Jinkela_buffer_1315 (
        .din(new_Jinkela_wire_2137),
        .dout(new_Jinkela_wire_2138)
    );

    bfr new_Jinkela_buffer_1352 (
        .din(new_Jinkela_wire_2191),
        .dout(new_Jinkela_wire_2192)
    );

    and_bb _1331_ (
        .a(new_Jinkela_wire_2886),
        .b(new_Jinkela_wire_1640),
        .c(_0500_)
    );

    bfr new_Jinkela_buffer_270 (
        .din(new_Jinkela_wire_482),
        .dout(new_Jinkela_wire_483)
    );

    bfr new_Jinkela_buffer_859 (
        .din(new_Jinkela_wire_1457),
        .dout(new_Jinkela_wire_1458)
    );

    and_ii _1332_ (
        .a(new_Jinkela_wire_2007),
        .b(new_Jinkela_wire_898),
        .c(_0501_)
    );

    spl2 new_Jinkela_splitter_79 (
        .a(new_Jinkela_wire_489),
        .b(new_Jinkela_wire_490),
        .c(new_Jinkela_wire_491)
    );

    bfr new_Jinkela_buffer_879 (
        .din(_0531_),
        .dout(new_Jinkela_wire_1498)
    );

    or_bi _1333_ (
        .a(new_Jinkela_wire_2708),
        .b(new_Jinkela_wire_2213),
        .c(_0502_)
    );

    spl2 new_Jinkela_splitter_77 (
        .a(new_Jinkela_wire_483),
        .b(new_Jinkela_wire_484),
        .c(new_Jinkela_wire_485)
    );

    bfr new_Jinkela_buffer_860 (
        .din(new_Jinkela_wire_1458),
        .dout(new_Jinkela_wire_1459)
    );

    and_bi _1334_ (
        .a(new_Jinkela_wire_2707),
        .b(new_Jinkela_wire_2212),
        .c(_0503_)
    );

    bfr new_Jinkela_buffer_874 (
        .din(new_Jinkela_wire_1478),
        .dout(new_Jinkela_wire_1479)
    );

    bfr new_Jinkela_buffer_273 (
        .din(new_Jinkela_wire_491),
        .dout(new_Jinkela_wire_492)
    );

    or_bb _1335_ (
        .a(_0503_),
        .b(new_Jinkela_wire_1462),
        .c(_0504_)
    );

    bfr new_Jinkela_buffer_861 (
        .din(new_Jinkela_wire_1459),
        .dout(new_Jinkela_wire_1460)
    );

    spl2 new_Jinkela_splitter_85 (
        .a(new_Jinkela_wire_512),
        .b(new_Jinkela_wire_513),
        .c(new_Jinkela_wire_514)
    );

    and_bi _1336_ (
        .a(new_Jinkela_wire_3310),
        .b(_0504_),
        .c(_0505_)
    );

    bfr new_Jinkela_buffer_275 (
        .din(new_Jinkela_wire_493),
        .dout(new_Jinkela_wire_494)
    );

    bfr new_Jinkela_buffer_878 (
        .din(new_Jinkela_wire_1492),
        .dout(new_Jinkela_wire_1493)
    );

    spl2 new_Jinkela_splitter_86 (
        .a(new_Jinkela_wire_514),
        .b(new_Jinkela_wire_515),
        .c(new_Jinkela_wire_516)
    );

    or_bb _1337_ (
        .a(_0505_),
        .b(new_Jinkela_wire_1019),
        .c(new_net_3)
    );

    bfr new_Jinkela_buffer_862 (
        .din(new_Jinkela_wire_1460),
        .dout(new_Jinkela_wire_1461)
    );

    and_bi _1338_ (
        .a(new_Jinkela_wire_918),
        .b(new_Jinkela_wire_2461),
        .c(_0506_)
    );

    bfr new_Jinkela_buffer_875 (
        .din(new_Jinkela_wire_1479),
        .dout(new_Jinkela_wire_1480)
    );

    bfr new_Jinkela_buffer_274 (
        .din(new_Jinkela_wire_492),
        .dout(new_Jinkela_wire_493)
    );

    or_bb _1339_ (
        .a(new_Jinkela_wire_2108),
        .b(new_Jinkela_wire_1076),
        .c(_0507_)
    );

    spl2 new_Jinkela_splitter_95 (
        .a(G26),
        .b(new_Jinkela_wire_561),
        .c(new_Jinkela_wire_562)
    );

    bfr new_Jinkela_buffer_863 (
        .din(new_Jinkela_wire_1461),
        .dout(new_Jinkela_wire_1462)
    );

    bfr new_Jinkela_buffer_301 (
        .din(G38),
        .dout(new_Jinkela_wire_553)
    );

    and_bi _1340_ (
        .a(new_Jinkela_wire_245),
        .b(new_Jinkela_wire_1886),
        .c(_0508_)
    );

    spl2 new_Jinkela_splitter_97 (
        .a(G7),
        .b(new_Jinkela_wire_567),
        .c(new_Jinkela_wire_569)
    );

    spl2 new_Jinkela_splitter_241 (
        .a(_0197_),
        .b(new_Jinkela_wire_1499),
        .c(new_Jinkela_wire_1500)
    );

    spl3L new_Jinkela_splitter_242 (
        .a(_0346_),
        .d(new_Jinkela_wire_1502),
        .b(new_Jinkela_wire_1503),
        .c(new_Jinkela_wire_1504)
    );

    spl2 new_Jinkela_splitter_80 (
        .a(new_Jinkela_wire_494),
        .b(new_Jinkela_wire_495),
        .c(new_Jinkela_wire_496)
    );

    and_bi _1341_ (
        .a(new_Jinkela_wire_727),
        .b(new_Jinkela_wire_2362),
        .c(_0509_)
    );

    bfr new_Jinkela_buffer_289 (
        .din(new_Jinkela_wire_536),
        .dout(new_Jinkela_wire_537)
    );

    bfr new_Jinkela_buffer_876 (
        .din(new_Jinkela_wire_1480),
        .dout(new_Jinkela_wire_1481)
    );

    or_bb _1342_ (
        .a(_0509_),
        .b(new_Jinkela_wire_969),
        .c(_0510_)
    );

    spl2 new_Jinkela_splitter_239 (
        .a(new_Jinkela_wire_1493),
        .b(new_Jinkela_wire_1494),
        .c(new_Jinkela_wire_1495)
    );

    spl2 new_Jinkela_splitter_81 (
        .a(new_Jinkela_wire_496),
        .b(new_Jinkela_wire_497),
        .c(new_Jinkela_wire_498)
    );

    or_ii _1343_ (
        .a(new_Jinkela_wire_281),
        .b(new_Jinkela_wire_735),
        .c(_0511_)
    );

    spl2 new_Jinkela_splitter_235 (
        .a(new_Jinkela_wire_1481),
        .b(new_Jinkela_wire_1482),
        .c(new_Jinkela_wire_1483)
    );

    spl3L new_Jinkela_splitter_88 (
        .a(new_Jinkela_wire_521),
        .d(new_Jinkela_wire_522),
        .b(new_Jinkela_wire_523),
        .c(new_Jinkela_wire_524)
    );

    and_bi _1344_ (
        .a(new_Jinkela_wire_3253),
        .b(new_Jinkela_wire_2420),
        .c(_0512_)
    );

    bfr new_Jinkela_buffer_281 (
        .din(new_Jinkela_wire_516),
        .dout(new_Jinkela_wire_517)
    );

    bfr new_Jinkela_buffer_880 (
        .din(new_Jinkela_wire_1500),
        .dout(new_Jinkela_wire_1501)
    );

    bfr new_Jinkela_buffer_276 (
        .din(new_Jinkela_wire_498),
        .dout(new_Jinkela_wire_499)
    );

    and_bi _1345_ (
        .a(new_Jinkela_wire_2052),
        .b(new_Jinkela_wire_1744),
        .c(_0513_)
    );

    or_bb _1346_ (
        .a(new_Jinkela_wire_2773),
        .b(_0512_),
        .c(_0514_)
    );

    bfr new_Jinkela_buffer_881 (
        .din(_0632_),
        .dout(new_Jinkela_wire_1505)
    );

    bfr new_Jinkela_buffer_882 (
        .din(_0422_),
        .dout(new_Jinkela_wire_1506)
    );

    spl2 new_Jinkela_splitter_87 (
        .a(new_Jinkela_wire_519),
        .b(new_Jinkela_wire_520),
        .c(new_Jinkela_wire_521)
    );

    or_bb _1347_ (
        .a(new_Jinkela_wire_3047),
        .b(_0510_),
        .c(_0515_)
    );

    spl2 new_Jinkela_splitter_243 (
        .a(_0011_),
        .b(new_Jinkela_wire_1514),
        .c(new_Jinkela_wire_1515)
    );

    spl2 new_Jinkela_splitter_82 (
        .a(new_Jinkela_wire_499),
        .b(new_Jinkela_wire_500),
        .c(new_Jinkela_wire_501)
    );

    and_bi _1348_ (
        .a(new_Jinkela_wire_1723),
        .b(new_Jinkela_wire_3004),
        .c(_0516_)
    );

    bfr new_Jinkela_buffer_883 (
        .din(new_Jinkela_wire_1506),
        .dout(new_Jinkela_wire_1507)
    );

    bfr new_Jinkela_buffer_890 (
        .din(_0744_),
        .dout(new_Jinkela_wire_1516)
    );

    spl3L new_Jinkela_splitter_83 (
        .a(new_Jinkela_wire_501),
        .d(new_Jinkela_wire_502),
        .b(new_Jinkela_wire_503),
        .c(new_Jinkela_wire_504)
    );

    and_bi _1349_ (
        .a(new_Jinkela_wire_217),
        .b(new_Jinkela_wire_522),
        .c(_0517_)
    );

    spl2 new_Jinkela_splitter_89 (
        .a(new_Jinkela_wire_524),
        .b(new_Jinkela_wire_525),
        .c(new_Jinkela_wire_526)
    );

    and_ii _1350_ (
        .a(new_Jinkela_wire_2272),
        .b(new_Jinkela_wire_1131),
        .c(_0518_)
    );

    bfr new_Jinkela_buffer_892 (
        .din(new_Jinkela_wire_1517),
        .dout(new_Jinkela_wire_1518)
    );

    bfr new_Jinkela_buffer_898 (
        .din(_0337_),
        .dout(new_Jinkela_wire_1532)
    );

    bfr new_Jinkela_buffer_282 (
        .din(new_Jinkela_wire_517),
        .dout(new_Jinkela_wire_518)
    );

    or_bb _1351_ (
        .a(_0518_),
        .b(new_Jinkela_wire_3090),
        .c(_0519_)
    );

    bfr new_Jinkela_buffer_884 (
        .din(new_Jinkela_wire_1507),
        .dout(new_Jinkela_wire_1508)
    );

    bfr new_Jinkela_buffer_277 (
        .din(new_Jinkela_wire_504),
        .dout(new_Jinkela_wire_505)
    );

    or_bb _1352_ (
        .a(new_Jinkela_wire_3180),
        .b(_0516_),
        .c(_0520_)
    );

    spl2 new_Jinkela_splitter_93 (
        .a(new_Jinkela_wire_539),
        .b(new_Jinkela_wire_540),
        .c(new_Jinkela_wire_541)
    );

    or_bb _1353_ (
        .a(_0520_),
        .b(new_Jinkela_wire_2577),
        .c(_0521_)
    );

    bfr new_Jinkela_buffer_303 (
        .din(new_Jinkela_wire_554),
        .dout(new_Jinkela_wire_555)
    );

    bfr new_Jinkela_buffer_885 (
        .din(new_Jinkela_wire_1508),
        .dout(new_Jinkela_wire_1509)
    );

    bfr new_Jinkela_buffer_278 (
        .din(new_Jinkela_wire_505),
        .dout(new_Jinkela_wire_506)
    );

    or_bi _1354_ (
        .a(new_Jinkela_wire_1134),
        .b(new_Jinkela_wire_472),
        .c(_0522_)
    );

    spl2 new_Jinkela_splitter_245 (
        .a(_0554_),
        .b(new_Jinkela_wire_1523),
        .c(new_Jinkela_wire_1524)
    );

    bfr new_Jinkela_buffer_891 (
        .din(new_Jinkela_wire_1516),
        .dout(new_Jinkela_wire_1517)
    );

    and_bi _1355_ (
        .a(new_Jinkela_wire_188),
        .b(new_Jinkela_wire_1878),
        .c(_0523_)
    );

    bfr new_Jinkela_buffer_886 (
        .din(new_Jinkela_wire_1509),
        .dout(new_Jinkela_wire_1510)
    );

    bfr new_Jinkela_buffer_279 (
        .din(new_Jinkela_wire_506),
        .dout(new_Jinkela_wire_507)
    );

    and_bi _1356_ (
        .a(new_Jinkela_wire_503),
        .b(new_Jinkela_wire_1137),
        .c(_0524_)
    );

    or_bb _1357_ (
        .a(new_Jinkela_wire_2215),
        .b(new_Jinkela_wire_3290),
        .c(_0525_)
    );

    bfr new_Jinkela_buffer_284 (
        .din(new_Jinkela_wire_526),
        .dout(new_Jinkela_wire_527)
    );

    bfr new_Jinkela_buffer_887 (
        .din(new_Jinkela_wire_1510),
        .dout(new_Jinkela_wire_1511)
    );

    and_bi _1358_ (
        .a(new_Jinkela_wire_2410),
        .b(_0525_),
        .c(_0526_)
    );

    spl2 new_Jinkela_splitter_92 (
        .a(new_Jinkela_wire_537),
        .b(new_Jinkela_wire_538),
        .c(new_Jinkela_wire_539)
    );

    and_ii _1359_ (
        .a(new_Jinkela_wire_1178),
        .b(new_Jinkela_wire_2361),
        .c(_0527_)
    );

    bfr new_Jinkela_buffer_888 (
        .din(new_Jinkela_wire_1511),
        .dout(new_Jinkela_wire_1512)
    );

    or_bb _1360_ (
        .a(_0527_),
        .b(new_Jinkela_wire_829),
        .c(_0528_)
    );

    bfr new_Jinkela_buffer_285 (
        .din(new_Jinkela_wire_527),
        .dout(new_Jinkela_wire_528)
    );

    spl2 new_Jinkela_splitter_247 (
        .a(_0556_),
        .b(new_Jinkela_wire_1530),
        .c(new_Jinkela_wire_1531)
    );

    and_bi _1361_ (
        .a(new_Jinkela_wire_1689),
        .b(new_Jinkela_wire_1748),
        .c(_0529_)
    );

    bfr new_Jinkela_buffer_889 (
        .din(new_Jinkela_wire_1512),
        .dout(new_Jinkela_wire_1513)
    );

    and_bi _1362_ (
        .a(new_Jinkela_wire_668),
        .b(new_Jinkela_wire_2415),
        .c(_0530_)
    );

    bfr new_Jinkela_buffer_286 (
        .din(new_Jinkela_wire_528),
        .dout(new_Jinkela_wire_529)
    );

    bfr new_Jinkela_buffer_895 (
        .din(new_Jinkela_wire_1524),
        .dout(new_Jinkela_wire_1525)
    );

    bfr new_Jinkela_buffer_893 (
        .din(new_Jinkela_wire_1518),
        .dout(new_Jinkela_wire_1519)
    );

    or_bb _1363_ (
        .a(_0530_),
        .b(new_Jinkela_wire_1194),
        .c(_0531_)
    );

    bfr new_Jinkela_buffer_290 (
        .din(new_Jinkela_wire_541),
        .dout(new_Jinkela_wire_542)
    );

    or_bb _1364_ (
        .a(new_Jinkela_wire_1498),
        .b(_0528_),
        .c(_0532_)
    );

    bfr new_Jinkela_buffer_287 (
        .din(new_Jinkela_wire_529),
        .dout(new_Jinkela_wire_530)
    );

    bfr new_Jinkela_buffer_894 (
        .din(new_Jinkela_wire_1519),
        .dout(new_Jinkela_wire_1520)
    );

    or_bb _1365_ (
        .a(_0532_),
        .b(new_Jinkela_wire_1090),
        .c(_0533_)
    );

    bfr new_Jinkela_buffer_896 (
        .din(new_Jinkela_wire_1525),
        .dout(new_Jinkela_wire_1526)
    );

    and_bi _1366_ (
        .a(_0526_),
        .b(_0533_),
        .c(_0534_)
    );

    spl2 new_Jinkela_splitter_90 (
        .a(new_Jinkela_wire_530),
        .b(new_Jinkela_wire_531),
        .c(new_Jinkela_wire_532)
    );

    spl2 new_Jinkela_splitter_244 (
        .a(new_Jinkela_wire_1520),
        .b(new_Jinkela_wire_1521),
        .c(new_Jinkela_wire_1522)
    );

    and_bi _1367_ (
        .a(_0521_),
        .b(new_Jinkela_wire_1236),
        .c(_0535_)
    );

    bfr new_Jinkela_buffer_288 (
        .din(new_Jinkela_wire_532),
        .dout(new_Jinkela_wire_533)
    );

    bfr new_Jinkela_buffer_924 (
        .din(new_Jinkela_wire_1566),
        .dout(new_Jinkela_wire_1567)
    );

    and_bi _1368_ (
        .a(new_Jinkela_wire_1906),
        .b(_0535_),
        .c(_0536_)
    );

    bfr new_Jinkela_buffer_302 (
        .din(new_Jinkela_wire_553),
        .dout(new_Jinkela_wire_554)
    );

    bfr new_Jinkela_buffer_897 (
        .din(new_Jinkela_wire_1526),
        .dout(new_Jinkela_wire_1527)
    );

    bfr new_Jinkela_buffer_307 (
        .din(new_Jinkela_wire_562),
        .dout(new_Jinkela_wire_563)
    );

    or_bb _1369_ (
        .a(_0536_),
        .b(new_Jinkela_wire_1339),
        .c(_0537_)
    );

    spl4L new_Jinkela_splitter_98 (
        .a(new_Jinkela_wire_569),
        .d(new_Jinkela_wire_570),
        .e(new_Jinkela_wire_571),
        .b(new_Jinkela_wire_572),
        .c(new_Jinkela_wire_573)
    );

    bfr new_Jinkela_buffer_925 (
        .din(_0171_),
        .dout(new_Jinkela_wire_1568)
    );

    bfr new_Jinkela_buffer_291 (
        .din(new_Jinkela_wire_542),
        .dout(new_Jinkela_wire_543)
    );

    and_bi _1370_ (
        .a(_0507_),
        .b(new_Jinkela_wire_1159),
        .c(_0538_)
    );

    bfr new_Jinkela_buffer_923 (
        .din(_0693_),
        .dout(new_Jinkela_wire_1566)
    );

    and_ii _0844_ (
        .a(new_Jinkela_wire_768),
        .b(new_Jinkela_wire_303),
        .c(_0018_)
    );

    spl2 new_Jinkela_splitter_94 (
        .a(new_Jinkela_wire_555),
        .b(new_Jinkela_wire_556),
        .c(new_Jinkela_wire_557)
    );

    and_bi _1371_ (
        .a(new_Jinkela_wire_2545),
        .b(new_Jinkela_wire_1504),
        .c(_0539_)
    );

    spl2 new_Jinkela_splitter_246 (
        .a(new_Jinkela_wire_1527),
        .b(new_Jinkela_wire_1528),
        .c(new_Jinkela_wire_1529)
    );

    bfr new_Jinkela_buffer_292 (
        .din(new_Jinkela_wire_543),
        .dout(new_Jinkela_wire_544)
    );

    or_bb _1372_ (
        .a(_0539_),
        .b(new_Jinkela_wire_1323),
        .c(_0540_)
    );

    bfr new_Jinkela_buffer_899 (
        .din(new_Jinkela_wire_1532),
        .dout(new_Jinkela_wire_1533)
    );

    bfr new_Jinkela_buffer_1614 (
        .din(new_Jinkela_wire_2617),
        .dout(new_Jinkela_wire_2618)
    );

    bfr new_Jinkela_buffer_1690 (
        .din(new_Jinkela_wire_2712),
        .dout(new_Jinkela_wire_2713)
    );

    bfr new_Jinkela_buffer_1649 (
        .din(new_Jinkela_wire_2666),
        .dout(new_Jinkela_wire_2667)
    );

    bfr new_Jinkela_buffer_1615 (
        .din(new_Jinkela_wire_2618),
        .dout(new_Jinkela_wire_2619)
    );

    spl2 new_Jinkela_splitter_394 (
        .a(new_Jinkela_wire_2706),
        .b(new_Jinkela_wire_2707),
        .c(new_Jinkela_wire_2708)
    );

    bfr new_Jinkela_buffer_1616 (
        .din(new_Jinkela_wire_2619),
        .dout(new_Jinkela_wire_2620)
    );

    bfr new_Jinkela_buffer_1662 (
        .din(new_Jinkela_wire_2679),
        .dout(new_Jinkela_wire_2680)
    );

    bfr new_Jinkela_buffer_1650 (
        .din(new_Jinkela_wire_2667),
        .dout(new_Jinkela_wire_2668)
    );

    bfr new_Jinkela_buffer_1617 (
        .din(new_Jinkela_wire_2620),
        .dout(new_Jinkela_wire_2621)
    );

    bfr new_Jinkela_buffer_1618 (
        .din(new_Jinkela_wire_2621),
        .dout(new_Jinkela_wire_2622)
    );

    bfr new_Jinkela_buffer_1651 (
        .din(new_Jinkela_wire_2668),
        .dout(new_Jinkela_wire_2669)
    );

    bfr new_Jinkela_buffer_1619 (
        .din(new_Jinkela_wire_2622),
        .dout(new_Jinkela_wire_2623)
    );

    bfr new_Jinkela_buffer_1620 (
        .din(new_Jinkela_wire_2623),
        .dout(new_Jinkela_wire_2624)
    );

    bfr new_Jinkela_buffer_1663 (
        .din(new_Jinkela_wire_2680),
        .dout(new_Jinkela_wire_2681)
    );

    bfr new_Jinkela_buffer_1652 (
        .din(new_Jinkela_wire_2669),
        .dout(new_Jinkela_wire_2670)
    );

    bfr new_Jinkela_buffer_1621 (
        .din(new_Jinkela_wire_2624),
        .dout(new_Jinkela_wire_2625)
    );

    bfr new_Jinkela_buffer_1622 (
        .din(new_Jinkela_wire_2625),
        .dout(new_Jinkela_wire_2626)
    );

    and_bi _0823_ (
        .a(new_Jinkela_wire_1684),
        .b(new_Jinkela_wire_2305),
        .c(_0796_)
    );

    spl2 new_Jinkela_splitter_396 (
        .a(_0008_),
        .b(new_Jinkela_wire_2722),
        .c(new_Jinkela_wire_2723)
    );

    and_ii _0801_ (
        .a(new_Jinkela_wire_595),
        .b(new_Jinkela_wire_156),
        .c(_0652_)
    );

    bfr new_Jinkela_buffer_1653 (
        .din(new_Jinkela_wire_2670),
        .dout(new_Jinkela_wire_2671)
    );

    and_ii _0799_ (
        .a(new_Jinkela_wire_709),
        .b(new_Jinkela_wire_218),
        .c(_0631_)
    );

    bfr new_Jinkela_buffer_1623 (
        .din(new_Jinkela_wire_2626),
        .dout(new_Jinkela_wire_2627)
    );

    or_bb _0800_ (
        .a(new_Jinkela_wire_3285),
        .b(new_Jinkela_wire_2049),
        .c(new_net_1475)
    );

    bfr new_Jinkela_buffer_1698 (
        .din(_0649_),
        .dout(new_Jinkela_wire_2721)
    );

    inv _0798_ (
        .din(new_Jinkela_wire_323),
        .dout(_0620_)
    );

    bfr new_Jinkela_buffer_1624 (
        .din(new_Jinkela_wire_2627),
        .dout(new_Jinkela_wire_2628)
    );

    and_bi _0802_ (
        .a(new_Jinkela_wire_307),
        .b(new_Jinkela_wire_198),
        .c(_0662_)
    );

    bfr new_Jinkela_buffer_1664 (
        .din(new_Jinkela_wire_2681),
        .dout(new_Jinkela_wire_2682)
    );

    and_bi _0806_ (
        .a(new_Jinkela_wire_777),
        .b(new_Jinkela_wire_275),
        .c(_0705_)
    );

    bfr new_Jinkela_buffer_1654 (
        .din(new_Jinkela_wire_2671),
        .dout(new_Jinkela_wire_2672)
    );

    bfr new_Jinkela_buffer_1625 (
        .din(new_Jinkela_wire_2628),
        .dout(new_Jinkela_wire_2629)
    );

    or_bi _0805_ (
        .a(new_Jinkela_wire_215),
        .b(new_Jinkela_wire_513),
        .c(_0695_)
    );

    and_bi _0803_ (
        .a(new_Jinkela_wire_168),
        .b(new_Jinkela_wire_266),
        .c(_0673_)
    );

    bfr new_Jinkela_buffer_1626 (
        .din(new_Jinkela_wire_2629),
        .dout(new_Jinkela_wire_2630)
    );

    or_bb _0815_ (
        .a(_0785_),
        .b(_0756_),
        .c(_0788_)
    );

    and_ii _0804_ (
        .a(new_Jinkela_wire_2842),
        .b(_0662_),
        .c(_0684_)
    );

    bfr new_Jinkela_buffer_1655 (
        .din(new_Jinkela_wire_2672),
        .dout(new_Jinkela_wire_2673)
    );

    or_bi _0807_ (
        .a(new_Jinkela_wire_1202),
        .b(_0695_),
        .c(_0716_)
    );

    bfr new_Jinkela_buffer_1627 (
        .din(new_Jinkela_wire_2630),
        .dout(new_Jinkela_wire_2631)
    );

    and_bi _0808_ (
        .a(_0684_),
        .b(_0716_),
        .c(_0727_)
    );

    bfr new_Jinkela_buffer_1699 (
        .din(_0639_),
        .dout(new_Jinkela_wire_2724)
    );

    and_bi _0809_ (
        .a(new_Jinkela_wire_257),
        .b(new_Jinkela_wire_325),
        .c(_0736_)
    );

    bfr new_Jinkela_buffer_1628 (
        .din(new_Jinkela_wire_2631),
        .dout(new_Jinkela_wire_2632)
    );

    and_bi _0810_ (
        .a(new_Jinkela_wire_476),
        .b(new_Jinkela_wire_703),
        .c(_0746_)
    );

    bfr new_Jinkela_buffer_1665 (
        .din(new_Jinkela_wire_2682),
        .dout(new_Jinkela_wire_2683)
    );

    bfr new_Jinkela_buffer_1656 (
        .din(new_Jinkela_wire_2673),
        .dout(new_Jinkela_wire_2674)
    );

    or_bb _0811_ (
        .a(_0746_),
        .b(_0736_),
        .c(_0756_)
    );

    bfr new_Jinkela_buffer_1629 (
        .din(new_Jinkela_wire_2632),
        .dout(new_Jinkela_wire_2633)
    );

    and_bi _0812_ (
        .a(new_Jinkela_wire_767),
        .b(new_Jinkela_wire_733),
        .c(_0764_)
    );

    and_bi _0813_ (
        .a(new_Jinkela_wire_36),
        .b(new_Jinkela_wire_570),
        .c(_0775_)
    );

    bfr new_Jinkela_buffer_1630 (
        .din(new_Jinkela_wire_2633),
        .dout(new_Jinkela_wire_2634)
    );

    or_bb _0814_ (
        .a(_0775_),
        .b(_0764_),
        .c(_0785_)
    );

    bfr new_Jinkela_buffer_1691 (
        .din(new_Jinkela_wire_2713),
        .dout(new_Jinkela_wire_2714)
    );

    bfr new_Jinkela_buffer_1631 (
        .din(new_Jinkela_wire_2634),
        .dout(new_Jinkela_wire_2635)
    );

    and_bi _0816_ (
        .a(_0727_),
        .b(new_Jinkela_wire_2790),
        .c(_0789_)
    );

    bfr new_Jinkela_buffer_1666 (
        .din(new_Jinkela_wire_2683),
        .dout(new_Jinkela_wire_2684)
    );

    or_bb _0817_ (
        .a(_0789_),
        .b(new_Jinkela_wire_3326),
        .c(_0790_)
    );

    bfr new_Jinkela_buffer_1632 (
        .din(new_Jinkela_wire_2635),
        .dout(new_Jinkela_wire_2636)
    );

    inv _0818_ (
        .din(new_Jinkela_wire_149),
        .dout(_0791_)
    );

    or_bi _0819_ (
        .a(new_Jinkela_wire_590),
        .b(new_Jinkela_wire_794),
        .c(_0792_)
    );

    bfr new_Jinkela_buffer_1701 (
        .din(_0418_),
        .dout(new_Jinkela_wire_2726)
    );

    bfr new_Jinkela_buffer_1667 (
        .din(new_Jinkela_wire_2684),
        .dout(new_Jinkela_wire_2685)
    );

    and_bi _0820_ (
        .a(new_Jinkela_wire_2944),
        .b(new_Jinkela_wire_2507),
        .c(_0793_)
    );

    bfr new_Jinkela_buffer_1692 (
        .din(new_Jinkela_wire_2714),
        .dout(new_Jinkela_wire_2715)
    );

    inv _0821_ (
        .din(new_Jinkela_wire_572),
        .dout(_0794_)
    );

    bfr new_Jinkela_buffer_1668 (
        .din(new_Jinkela_wire_2685),
        .dout(new_Jinkela_wire_2686)
    );

    and_ii _0822_ (
        .a(new_Jinkela_wire_195),
        .b(new_Jinkela_wire_267),
        .c(_0795_)
    );

    bfr new_Jinkela_buffer_829 (
        .din(new_Jinkela_wire_1423),
        .dout(new_Jinkela_wire_1424)
    );

    bfr new_Jinkela_buffer_1316 (
        .din(new_Jinkela_wire_2138),
        .dout(new_Jinkela_wire_2139)
    );

    spl2 new_Jinkela_splitter_234 (
        .a(_0622_),
        .b(new_Jinkela_wire_1473),
        .c(new_Jinkela_wire_1474)
    );

    bfr new_Jinkela_buffer_845 (
        .din(new_Jinkela_wire_1441),
        .dout(new_Jinkela_wire_1442)
    );

    bfr new_Jinkela_buffer_1367 (
        .din(new_Jinkela_wire_2208),
        .dout(new_Jinkela_wire_2209)
    );

    bfr new_Jinkela_buffer_830 (
        .din(new_Jinkela_wire_1424),
        .dout(new_Jinkela_wire_1425)
    );

    bfr new_Jinkela_buffer_1317 (
        .din(new_Jinkela_wire_2139),
        .dout(new_Jinkela_wire_2140)
    );

    bfr new_Jinkela_buffer_1353 (
        .din(new_Jinkela_wire_2192),
        .dout(new_Jinkela_wire_2193)
    );

    bfr new_Jinkela_buffer_831 (
        .din(new_Jinkela_wire_1425),
        .dout(new_Jinkela_wire_1426)
    );

    bfr new_Jinkela_buffer_1318 (
        .din(new_Jinkela_wire_2140),
        .dout(new_Jinkela_wire_2141)
    );

    bfr new_Jinkela_buffer_846 (
        .din(new_Jinkela_wire_1442),
        .dout(new_Jinkela_wire_1443)
    );

    spl2 new_Jinkela_splitter_327 (
        .a(_0501_),
        .b(new_Jinkela_wire_2212),
        .c(new_Jinkela_wire_2213)
    );

    bfr new_Jinkela_buffer_832 (
        .din(new_Jinkela_wire_1426),
        .dout(new_Jinkela_wire_1427)
    );

    spl2 new_Jinkela_splitter_328 (
        .a(_0524_),
        .b(new_Jinkela_wire_2214),
        .c(new_Jinkela_wire_2215)
    );

    bfr new_Jinkela_buffer_1319 (
        .din(new_Jinkela_wire_2141),
        .dout(new_Jinkela_wire_2142)
    );

    spl2 new_Jinkela_splitter_240 (
        .a(_0747_),
        .b(new_Jinkela_wire_1496),
        .c(new_Jinkela_wire_1497)
    );

    bfr new_Jinkela_buffer_1354 (
        .din(new_Jinkela_wire_2193),
        .dout(new_Jinkela_wire_2194)
    );

    bfr new_Jinkela_buffer_833 (
        .din(new_Jinkela_wire_1427),
        .dout(new_Jinkela_wire_1428)
    );

    bfr new_Jinkela_buffer_1320 (
        .din(new_Jinkela_wire_2142),
        .dout(new_Jinkela_wire_2143)
    );

    spl3L new_Jinkela_splitter_236 (
        .a(_0572_),
        .d(new_Jinkela_wire_1484),
        .b(new_Jinkela_wire_1485),
        .c(new_Jinkela_wire_1486)
    );

    bfr new_Jinkela_buffer_847 (
        .din(new_Jinkela_wire_1443),
        .dout(new_Jinkela_wire_1444)
    );

    bfr new_Jinkela_buffer_1369 (
        .din(new_Jinkela_wire_2210),
        .dout(new_Jinkela_wire_2211)
    );

    bfr new_Jinkela_buffer_834 (
        .din(new_Jinkela_wire_1428),
        .dout(new_Jinkela_wire_1429)
    );

    bfr new_Jinkela_buffer_1321 (
        .din(new_Jinkela_wire_2143),
        .dout(new_Jinkela_wire_2144)
    );

    bfr new_Jinkela_buffer_865 (
        .din(new_Jinkela_wire_1467),
        .dout(new_Jinkela_wire_1468)
    );

    bfr new_Jinkela_buffer_1355 (
        .din(new_Jinkela_wire_2194),
        .dout(new_Jinkela_wire_2195)
    );

    bfr new_Jinkela_buffer_835 (
        .din(new_Jinkela_wire_1429),
        .dout(new_Jinkela_wire_1430)
    );

    bfr new_Jinkela_buffer_1322 (
        .din(new_Jinkela_wire_2144),
        .dout(new_Jinkela_wire_2145)
    );

    bfr new_Jinkela_buffer_848 (
        .din(new_Jinkela_wire_1444),
        .dout(new_Jinkela_wire_1445)
    );

    bfr new_Jinkela_buffer_1418 (
        .din(_0517_),
        .dout(new_Jinkela_wire_2266)
    );

    bfr new_Jinkela_buffer_836 (
        .din(new_Jinkela_wire_1430),
        .dout(new_Jinkela_wire_1431)
    );

    bfr new_Jinkela_buffer_1323 (
        .din(new_Jinkela_wire_2145),
        .dout(new_Jinkela_wire_2146)
    );

    bfr new_Jinkela_buffer_866 (
        .din(new_Jinkela_wire_1468),
        .dout(new_Jinkela_wire_1469)
    );

    bfr new_Jinkela_buffer_1356 (
        .din(new_Jinkela_wire_2195),
        .dout(new_Jinkela_wire_2196)
    );

    bfr new_Jinkela_buffer_837 (
        .din(new_Jinkela_wire_1431),
        .dout(new_Jinkela_wire_1432)
    );

    bfr new_Jinkela_buffer_1324 (
        .din(new_Jinkela_wire_2146),
        .dout(new_Jinkela_wire_2147)
    );

    bfr new_Jinkela_buffer_849 (
        .din(new_Jinkela_wire_1445),
        .dout(new_Jinkela_wire_1446)
    );

    bfr new_Jinkela_buffer_838 (
        .din(new_Jinkela_wire_1432),
        .dout(new_Jinkela_wire_1433)
    );

    bfr new_Jinkela_buffer_1370 (
        .din(_0285_),
        .dout(new_Jinkela_wire_2216)
    );

    bfr new_Jinkela_buffer_1325 (
        .din(new_Jinkela_wire_2147),
        .dout(new_Jinkela_wire_2148)
    );

    bfr new_Jinkela_buffer_1357 (
        .din(new_Jinkela_wire_2196),
        .dout(new_Jinkela_wire_2197)
    );

    bfr new_Jinkela_buffer_839 (
        .din(new_Jinkela_wire_1433),
        .dout(new_Jinkela_wire_1434)
    );

    bfr new_Jinkela_buffer_1326 (
        .din(new_Jinkela_wire_2148),
        .dout(new_Jinkela_wire_2149)
    );

    spl3L new_Jinkela_splitter_238 (
        .a(_0753_),
        .d(new_Jinkela_wire_1490),
        .b(new_Jinkela_wire_1491),
        .c(new_Jinkela_wire_1492)
    );

    bfr new_Jinkela_buffer_850 (
        .din(new_Jinkela_wire_1446),
        .dout(new_Jinkela_wire_1447)
    );

    bfr new_Jinkela_buffer_840 (
        .din(new_Jinkela_wire_1434),
        .dout(new_Jinkela_wire_1435)
    );

    bfr new_Jinkela_buffer_1327 (
        .din(new_Jinkela_wire_2149),
        .dout(new_Jinkela_wire_2150)
    );

    bfr new_Jinkela_buffer_867 (
        .din(new_Jinkela_wire_1469),
        .dout(new_Jinkela_wire_1470)
    );

    spl2 new_Jinkela_splitter_326 (
        .a(new_Jinkela_wire_2197),
        .b(new_Jinkela_wire_2198),
        .c(new_Jinkela_wire_2199)
    );

    bfr new_Jinkela_buffer_851 (
        .din(new_Jinkela_wire_1447),
        .dout(new_Jinkela_wire_1448)
    );

    bfr new_Jinkela_buffer_1328 (
        .din(new_Jinkela_wire_2150),
        .dout(new_Jinkela_wire_2151)
    );

    bfr new_Jinkela_buffer_870 (
        .din(new_Jinkela_wire_1474),
        .dout(new_Jinkela_wire_1475)
    );

    bfr new_Jinkela_buffer_1358 (
        .din(new_Jinkela_wire_2199),
        .dout(new_Jinkela_wire_2200)
    );

    spl2 new_Jinkela_splitter_237 (
        .a(_0323_),
        .b(new_Jinkela_wire_1488),
        .c(new_Jinkela_wire_1489)
    );

    bfr new_Jinkela_buffer_852 (
        .din(new_Jinkela_wire_1448),
        .dout(new_Jinkela_wire_1449)
    );

    bfr new_Jinkela_buffer_1329 (
        .din(new_Jinkela_wire_2151),
        .dout(new_Jinkela_wire_2152)
    );

    bfr new_Jinkela_buffer_868 (
        .din(new_Jinkela_wire_1470),
        .dout(new_Jinkela_wire_1471)
    );

    bfr new_Jinkela_buffer_1417 (
        .din(_0222_),
        .dout(new_Jinkela_wire_2265)
    );

    bfr new_Jinkela_buffer_1371 (
        .din(new_Jinkela_wire_2216),
        .dout(new_Jinkela_wire_2217)
    );

    bfr new_Jinkela_buffer_853 (
        .din(new_Jinkela_wire_1449),
        .dout(new_Jinkela_wire_1450)
    );

    bfr new_Jinkela_buffer_1330 (
        .din(new_Jinkela_wire_2152),
        .dout(new_Jinkela_wire_2153)
    );

    bfr new_Jinkela_buffer_877 (
        .din(new_Jinkela_wire_1486),
        .dout(new_Jinkela_wire_1487)
    );

    bfr new_Jinkela_buffer_1423 (
        .din(_0741_),
        .dout(new_Jinkela_wire_2273)
    );

    spl2 new_Jinkela_splitter_231 (
        .a(new_Jinkela_wire_1450),
        .b(new_Jinkela_wire_1451),
        .c(new_Jinkela_wire_1452)
    );

    bfr new_Jinkela_buffer_1331 (
        .din(new_Jinkela_wire_2153),
        .dout(new_Jinkela_wire_2154)
    );

    bfr new_Jinkela_buffer_854 (
        .din(new_Jinkela_wire_1452),
        .dout(new_Jinkela_wire_1453)
    );

    bfr new_Jinkela_buffer_1359 (
        .din(new_Jinkela_wire_2200),
        .dout(new_Jinkela_wire_2201)
    );

    bfr new_Jinkela_buffer_869 (
        .din(new_Jinkela_wire_1471),
        .dout(new_Jinkela_wire_1472)
    );

    bfr new_Jinkela_buffer_1332 (
        .din(new_Jinkela_wire_2154),
        .dout(new_Jinkela_wire_2155)
    );

    bfr new_Jinkela_buffer_871 (
        .din(new_Jinkela_wire_1475),
        .dout(new_Jinkela_wire_1476)
    );

    bfr new_Jinkela_buffer_1372 (
        .din(new_Jinkela_wire_2217),
        .dout(new_Jinkela_wire_2218)
    );

    bfr new_Jinkela_buffer_855 (
        .din(new_Jinkela_wire_1453),
        .dout(new_Jinkela_wire_1454)
    );

    bfr new_Jinkela_buffer_1333 (
        .din(new_Jinkela_wire_2155),
        .dout(new_Jinkela_wire_2156)
    );

    bfr new_Jinkela_buffer_1360 (
        .din(new_Jinkela_wire_2201),
        .dout(new_Jinkela_wire_2202)
    );

    bfr new_Jinkela_buffer_872 (
        .din(new_Jinkela_wire_1476),
        .dout(new_Jinkela_wire_1477)
    );

    bfr new_Jinkela_buffer_856 (
        .din(new_Jinkela_wire_1454),
        .dout(new_Jinkela_wire_1455)
    );

    bfr new_Jinkela_buffer_1334 (
        .din(new_Jinkela_wire_2156),
        .dout(new_Jinkela_wire_2157)
    );

    bfr new_Jinkela_buffer_857 (
        .din(new_Jinkela_wire_1455),
        .dout(new_Jinkela_wire_1456)
    );

    bfr new_Jinkela_buffer_1335 (
        .din(new_Jinkela_wire_2157),
        .dout(new_Jinkela_wire_2158)
    );

    bfr new_Jinkela_buffer_1361 (
        .din(new_Jinkela_wire_2202),
        .dout(new_Jinkela_wire_2203)
    );

    bfr new_Jinkela_buffer_858 (
        .din(new_Jinkela_wire_1456),
        .dout(new_Jinkela_wire_1457)
    );

    bfr new_Jinkela_buffer_1336 (
        .din(new_Jinkela_wire_2158),
        .dout(new_Jinkela_wire_2159)
    );

    bfr new_Jinkela_buffer_873 (
        .din(new_Jinkela_wire_1477),
        .dout(new_Jinkela_wire_1478)
    );

    spl3L new_Jinkela_splitter_331 (
        .a(_0269_),
        .d(new_Jinkela_wire_2274),
        .b(new_Jinkela_wire_2275),
        .c(new_Jinkela_wire_2276)
    );

    and_bi _0995_ (
        .a(new_Jinkela_wire_2877),
        .b(new_Jinkela_wire_1237),
        .c(_0167_)
    );

    inv _0996_ (
        .din(new_Jinkela_wire_2310),
        .dout(_0168_)
    );

    and_bi _0997_ (
        .a(new_Jinkela_wire_3286),
        .b(new_Jinkela_wire_335),
        .c(_0169_)
    );

    or_bb _0998_ (
        .a(_0169_),
        .b(new_Jinkela_wire_2950),
        .c(_0170_)
    );

    and_bi _0999_ (
        .a(new_Jinkela_wire_1937),
        .b(new_Jinkela_wire_1283),
        .c(_0171_)
    );

    inv _1000_ (
        .din(new_Jinkela_wire_702),
        .dout(_0172_)
    );

    and_bi _1001_ (
        .a(new_Jinkela_wire_1712),
        .b(new_Jinkela_wire_3331),
        .c(_0173_)
    );

    or_bb _1002_ (
        .a(_0173_),
        .b(new_Jinkela_wire_1568),
        .c(_0174_)
    );

    and_bi _1003_ (
        .a(new_Jinkela_wire_2730),
        .b(_0174_),
        .c(_0175_)
    );

    or_bi _1004_ (
        .a(_0175_),
        .b(new_Jinkela_wire_3321),
        .c(_0176_)
    );

    and_bi _1005_ (
        .a(new_Jinkela_wire_442),
        .b(new_Jinkela_wire_601),
        .c(_0177_)
    );

    or_bb _1006_ (
        .a(new_Jinkela_wire_2046),
        .b(new_Jinkela_wire_3301),
        .c(_0178_)
    );

    or_bb _1007_ (
        .a(_0178_),
        .b(new_Jinkela_wire_3314),
        .c(_0179_)
    );

    and_bi _1008_ (
        .a(new_Jinkela_wire_342),
        .b(new_Jinkela_wire_2441),
        .c(_0180_)
    );

    and_bi _1009_ (
        .a(new_Jinkela_wire_3299),
        .b(new_Jinkela_wire_338),
        .c(_0181_)
    );

    or_bb _1010_ (
        .a(new_Jinkela_wire_1765),
        .b(_0180_),
        .c(_0182_)
    );

    or_bi _1011_ (
        .a(_0182_),
        .b(new_Jinkela_wire_2321),
        .c(_0183_)
    );

    or_bb _1012_ (
        .a(new_Jinkela_wire_3030),
        .b(new_Jinkela_wire_989),
        .c(_0184_)
    );

    or_bb _1013_ (
        .a(new_Jinkela_wire_412),
        .b(new_Jinkela_wire_283),
        .c(_0185_)
    );

    and_bi _1014_ (
        .a(new_Jinkela_wire_418),
        .b(new_Jinkela_wire_771),
        .c(_0186_)
    );

    and_bi _1015_ (
        .a(_0185_),
        .b(_0186_),
        .c(_0187_)
    );

    and_bi _1016_ (
        .a(_0184_),
        .b(new_Jinkela_wire_1333),
        .c(_0188_)
    );

    or_bb _1017_ (
        .a(new_Jinkela_wire_593),
        .b(new_Jinkela_wire_636),
        .c(_0189_)
    );

    or_bb _1018_ (
        .a(new_Jinkela_wire_2382),
        .b(new_Jinkela_wire_556),
        .c(_0190_)
    );

    and_ii _1019_ (
        .a(new_Jinkela_wire_592),
        .b(new_Jinkela_wire_635),
        .c(_0191_)
    );

    and_bi _1020_ (
        .a(new_Jinkela_wire_1140),
        .b(new_Jinkela_wire_1400),
        .c(_0192_)
    );

    and_bi _1021_ (
        .a(_0190_),
        .b(_0192_),
        .c(_0193_)
    );

    and_bi _1022_ (
        .a(_0188_),
        .b(new_Jinkela_wire_2209),
        .c(_0194_)
    );

    and_bi _1023_ (
        .a(new_Jinkela_wire_1050),
        .b(_0194_),
        .c(_0195_)
    );

    or_bb _1024_ (
        .a(new_Jinkela_wire_1203),
        .b(new_Jinkela_wire_3056),
        .c(_0196_)
    );

    and_bi _1025_ (
        .a(new_Jinkela_wire_1167),
        .b(new_Jinkela_wire_2992),
        .c(_0197_)
    );

    or_bi _1026_ (
        .a(new_Jinkela_wire_1204),
        .b(new_Jinkela_wire_2560),
        .c(_0198_)
    );

    and_bi _1027_ (
        .a(new_Jinkela_wire_2189),
        .b(new_Jinkela_wire_1168),
        .c(_0199_)
    );

    and_ii _1028_ (
        .a(new_Jinkela_wire_1279),
        .b(new_Jinkela_wire_1499),
        .c(_0200_)
    );

    and_bi _1029_ (
        .a(new_Jinkela_wire_1713),
        .b(new_Jinkela_wire_3306),
        .c(_0201_)
    );

    and_bi _1030_ (
        .a(new_Jinkela_wire_2442),
        .b(new_Jinkela_wire_1719),
        .c(_0202_)
    );

    or_bb _1031_ (
        .a(_0202_),
        .b(new_Jinkela_wire_916),
        .c(_0203_)
    );

    and_bb _1032_ (
        .a(new_Jinkela_wire_710),
        .b(new_Jinkela_wire_219),
        .c(_0204_)
    );

    or_bb _1033_ (
        .a(new_Jinkela_wire_3042),
        .b(new_Jinkela_wire_3287),
        .c(_0205_)
    );

    and_bi _1034_ (
        .a(new_Jinkela_wire_3191),
        .b(new_Jinkela_wire_809),
        .c(_0206_)
    );

    and_bi _1035_ (
        .a(new_Jinkela_wire_2945),
        .b(new_Jinkela_wire_1463),
        .c(_0207_)
    );

    and_bb _1036_ (
        .a(new_Jinkela_wire_440),
        .b(new_Jinkela_wire_221),
        .c(_0208_)
    );

    spl2 new_Jinkela_splitter_252 (
        .a(_0370_),
        .b(new_Jinkela_wire_1569),
        .c(new_Jinkela_wire_1570)
    );

    bfr new_Jinkela_buffer_926 (
        .din(_0417_),
        .dout(new_Jinkela_wire_1571)
    );

    and_bb _0845_ (
        .a(new_Jinkela_wire_769),
        .b(new_Jinkela_wire_304),
        .c(_0019_)
    );

    bfr new_Jinkela_buffer_900 (
        .din(new_Jinkela_wire_1533),
        .dout(new_Jinkela_wire_1534)
    );

    bfr new_Jinkela_buffer_927 (
        .din(new_Jinkela_wire_1571),
        .dout(new_Jinkela_wire_1572)
    );

    bfr new_Jinkela_buffer_901 (
        .din(new_Jinkela_wire_1534),
        .dout(new_Jinkela_wire_1535)
    );

    bfr new_Jinkela_buffer_902 (
        .din(new_Jinkela_wire_1535),
        .dout(new_Jinkela_wire_1536)
    );

    bfr new_Jinkela_buffer_932 (
        .din(new_net_1463),
        .dout(new_Jinkela_wire_1577)
    );

    bfr new_Jinkela_buffer_903 (
        .din(new_Jinkela_wire_1536),
        .dout(new_Jinkela_wire_1537)
    );

    bfr new_Jinkela_buffer_975 (
        .din(_0211_),
        .dout(new_Jinkela_wire_1620)
    );

    bfr new_Jinkela_buffer_904 (
        .din(new_Jinkela_wire_1537),
        .dout(new_Jinkela_wire_1538)
    );

    bfr new_Jinkela_buffer_928 (
        .din(new_Jinkela_wire_1572),
        .dout(new_Jinkela_wire_1573)
    );

    bfr new_Jinkela_buffer_905 (
        .din(new_Jinkela_wire_1538),
        .dout(new_Jinkela_wire_1539)
    );

    bfr new_Jinkela_buffer_933 (
        .din(new_Jinkela_wire_1577),
        .dout(new_Jinkela_wire_1578)
    );

    bfr new_Jinkela_buffer_906 (
        .din(new_Jinkela_wire_1539),
        .dout(new_Jinkela_wire_1540)
    );

    bfr new_Jinkela_buffer_929 (
        .din(new_Jinkela_wire_1573),
        .dout(new_Jinkela_wire_1574)
    );

    bfr new_Jinkela_buffer_907 (
        .din(new_Jinkela_wire_1540),
        .dout(new_Jinkela_wire_1541)
    );

    bfr new_Jinkela_buffer_976 (
        .din(_0551_),
        .dout(new_Jinkela_wire_1621)
    );

    spl2 new_Jinkela_splitter_254 (
        .a(_0033_),
        .b(new_Jinkela_wire_1625),
        .c(new_Jinkela_wire_1626)
    );

    bfr new_Jinkela_buffer_908 (
        .din(new_Jinkela_wire_1541),
        .dout(new_Jinkela_wire_1542)
    );

    bfr new_Jinkela_buffer_930 (
        .din(new_Jinkela_wire_1574),
        .dout(new_Jinkela_wire_1575)
    );

    bfr new_Jinkela_buffer_909 (
        .din(new_Jinkela_wire_1542),
        .dout(new_Jinkela_wire_1543)
    );

    bfr new_Jinkela_buffer_934 (
        .din(new_Jinkela_wire_1578),
        .dout(new_Jinkela_wire_1579)
    );

    bfr new_Jinkela_buffer_910 (
        .din(new_Jinkela_wire_1543),
        .dout(new_Jinkela_wire_1544)
    );

    bfr new_Jinkela_buffer_931 (
        .din(new_Jinkela_wire_1575),
        .dout(new_Jinkela_wire_1576)
    );

    bfr new_Jinkela_buffer_911 (
        .din(new_Jinkela_wire_1544),
        .dout(new_Jinkela_wire_1545)
    );

    bfr new_Jinkela_buffer_977 (
        .din(new_Jinkela_wire_1621),
        .dout(new_Jinkela_wire_1622)
    );

    bfr new_Jinkela_buffer_978 (
        .din(_0276_),
        .dout(new_Jinkela_wire_1627)
    );

    bfr new_Jinkela_buffer_912 (
        .din(new_Jinkela_wire_1545),
        .dout(new_Jinkela_wire_1546)
    );

    bfr new_Jinkela_buffer_935 (
        .din(new_Jinkela_wire_1579),
        .dout(new_Jinkela_wire_1580)
    );

    bfr new_Jinkela_buffer_913 (
        .din(new_Jinkela_wire_1546),
        .dout(new_Jinkela_wire_1547)
    );

    spl4L new_Jinkela_splitter_255 (
        .a(_0140_),
        .d(new_Jinkela_wire_1628),
        .e(new_Jinkela_wire_1629),
        .b(new_Jinkela_wire_1630),
        .c(new_Jinkela_wire_1631)
    );

    bfr new_Jinkela_buffer_914 (
        .din(new_Jinkela_wire_1547),
        .dout(new_Jinkela_wire_1548)
    );

    bfr new_Jinkela_buffer_936 (
        .din(new_Jinkela_wire_1580),
        .dout(new_Jinkela_wire_1581)
    );

    bfr new_Jinkela_buffer_915 (
        .din(new_Jinkela_wire_1548),
        .dout(new_Jinkela_wire_1549)
    );

    spl2 new_Jinkela_splitter_256 (
        .a(_0568_),
        .b(new_Jinkela_wire_1641),
        .c(new_Jinkela_wire_1642)
    );

    spl2 new_Jinkela_splitter_248 (
        .a(new_Jinkela_wire_1549),
        .b(new_Jinkela_wire_1550),
        .c(new_Jinkela_wire_1551)
    );

    spl3L new_Jinkela_splitter_249 (
        .a(new_Jinkela_wire_1551),
        .d(new_Jinkela_wire_1552),
        .b(new_Jinkela_wire_1553),
        .c(new_Jinkela_wire_1554)
    );

    bfr new_Jinkela_buffer_937 (
        .din(new_Jinkela_wire_1581),
        .dout(new_Jinkela_wire_1582)
    );

    spl2 new_Jinkela_splitter_253 (
        .a(new_Jinkela_wire_1622),
        .b(new_Jinkela_wire_1623),
        .c(new_Jinkela_wire_1624)
    );

    bfr new_Jinkela_buffer_916 (
        .din(new_Jinkela_wire_1554),
        .dout(new_Jinkela_wire_1555)
    );

    bfr new_Jinkela_buffer_938 (
        .din(new_Jinkela_wire_1582),
        .dout(new_Jinkela_wire_1583)
    );

    bfr new_Jinkela_buffer_917 (
        .din(new_Jinkela_wire_1555),
        .dout(new_Jinkela_wire_1556)
    );

    bfr new_Jinkela_buffer_918 (
        .din(new_Jinkela_wire_1556),
        .dout(new_Jinkela_wire_1557)
    );

    bfr new_Jinkela_buffer_1373 (
        .din(new_Jinkela_wire_2218),
        .dout(new_Jinkela_wire_2219)
    );

    bfr new_Jinkela_buffer_1337 (
        .din(new_Jinkela_wire_2159),
        .dout(new_Jinkela_wire_2160)
    );

    bfr new_Jinkela_buffer_1669 (
        .din(new_Jinkela_wire_2686),
        .dout(new_Jinkela_wire_2687)
    );

    bfr new_Jinkela_buffer_795 (
        .din(new_Jinkela_wire_1377),
        .dout(new_Jinkela_wire_1378)
    );

    bfr new_Jinkela_buffer_1362 (
        .din(new_Jinkela_wire_2203),
        .dout(new_Jinkela_wire_2204)
    );

    bfr new_Jinkela_buffer_1693 (
        .din(new_Jinkela_wire_2715),
        .dout(new_Jinkela_wire_2716)
    );

    spl2 new_Jinkela_splitter_226 (
        .a(_0625_),
        .b(new_Jinkela_wire_1404),
        .c(new_Jinkela_wire_1405)
    );

    bfr new_Jinkela_buffer_1338 (
        .din(new_Jinkela_wire_2160),
        .dout(new_Jinkela_wire_2161)
    );

    bfr new_Jinkela_buffer_1670 (
        .din(new_Jinkela_wire_2687),
        .dout(new_Jinkela_wire_2688)
    );

    spl3L new_Jinkela_splitter_227 (
        .a(_0247_),
        .d(new_Jinkela_wire_1406),
        .b(new_Jinkela_wire_1407),
        .c(new_Jinkela_wire_1408)
    );

    bfr new_Jinkela_buffer_796 (
        .din(new_Jinkela_wire_1378),
        .dout(new_Jinkela_wire_1379)
    );

    bfr new_Jinkela_buffer_1700 (
        .din(new_Jinkela_wire_2724),
        .dout(new_Jinkela_wire_2725)
    );

    bfr new_Jinkela_buffer_1419 (
        .din(new_Jinkela_wire_2266),
        .dout(new_Jinkela_wire_2267)
    );

    bfr new_Jinkela_buffer_1339 (
        .din(new_Jinkela_wire_2161),
        .dout(new_Jinkela_wire_2162)
    );

    bfr new_Jinkela_buffer_1671 (
        .din(new_Jinkela_wire_2688),
        .dout(new_Jinkela_wire_2689)
    );

    bfr new_Jinkela_buffer_819 (
        .din(new_Jinkela_wire_1408),
        .dout(new_Jinkela_wire_1409)
    );

    bfr new_Jinkela_buffer_797 (
        .din(new_Jinkela_wire_1379),
        .dout(new_Jinkela_wire_1380)
    );

    bfr new_Jinkela_buffer_1363 (
        .din(new_Jinkela_wire_2204),
        .dout(new_Jinkela_wire_2205)
    );

    bfr new_Jinkela_buffer_1694 (
        .din(new_Jinkela_wire_2716),
        .dout(new_Jinkela_wire_2717)
    );

    bfr new_Jinkela_buffer_1340 (
        .din(new_Jinkela_wire_2162),
        .dout(new_Jinkela_wire_2163)
    );

    bfr new_Jinkela_buffer_1672 (
        .din(new_Jinkela_wire_2689),
        .dout(new_Jinkela_wire_2690)
    );

    spl2 new_Jinkela_splitter_228 (
        .a(_0541_),
        .b(new_Jinkela_wire_1413),
        .c(new_Jinkela_wire_1414)
    );

    bfr new_Jinkela_buffer_798 (
        .din(new_Jinkela_wire_1380),
        .dout(new_Jinkela_wire_1381)
    );

    bfr new_Jinkela_buffer_1704 (
        .din(_0170_),
        .dout(new_Jinkela_wire_2729)
    );

    spl2 new_Jinkela_splitter_329 (
        .a(new_Jinkela_wire_2219),
        .b(new_Jinkela_wire_2220),
        .c(new_Jinkela_wire_2221)
    );

    bfr new_Jinkela_buffer_823 (
        .din(new_net_6),
        .dout(new_Jinkela_wire_1415)
    );

    bfr new_Jinkela_buffer_1341 (
        .din(new_Jinkela_wire_2163),
        .dout(new_Jinkela_wire_2164)
    );

    bfr new_Jinkela_buffer_1673 (
        .din(new_Jinkela_wire_2690),
        .dout(new_Jinkela_wire_2691)
    );

    spl2 new_Jinkela_splitter_230 (
        .a(_0406_),
        .b(new_Jinkela_wire_1439),
        .c(new_Jinkela_wire_1440)
    );

    bfr new_Jinkela_buffer_799 (
        .din(new_Jinkela_wire_1381),
        .dout(new_Jinkela_wire_1382)
    );

    bfr new_Jinkela_buffer_1364 (
        .din(new_Jinkela_wire_2205),
        .dout(new_Jinkela_wire_2206)
    );

    bfr new_Jinkela_buffer_1695 (
        .din(new_Jinkela_wire_2717),
        .dout(new_Jinkela_wire_2718)
    );

    bfr new_Jinkela_buffer_1674 (
        .din(new_Jinkela_wire_2691),
        .dout(new_Jinkela_wire_2692)
    );

    bfr new_Jinkela_buffer_1374 (
        .din(new_Jinkela_wire_2221),
        .dout(new_Jinkela_wire_2222)
    );

    bfr new_Jinkela_buffer_800 (
        .din(new_Jinkela_wire_1382),
        .dout(new_Jinkela_wire_1383)
    );

    bfr new_Jinkela_buffer_1365 (
        .din(new_Jinkela_wire_2206),
        .dout(new_Jinkela_wire_2207)
    );

    bfr new_Jinkela_buffer_1702 (
        .din(new_Jinkela_wire_2726),
        .dout(new_Jinkela_wire_2727)
    );

    bfr new_Jinkela_buffer_1675 (
        .din(new_Jinkela_wire_2692),
        .dout(new_Jinkela_wire_2693)
    );

    spl2 new_Jinkela_splitter_332 (
        .a(_0561_),
        .b(new_Jinkela_wire_2277),
        .c(new_Jinkela_wire_2278)
    );

    bfr new_Jinkela_buffer_820 (
        .din(new_Jinkela_wire_1409),
        .dout(new_Jinkela_wire_1410)
    );

    bfr new_Jinkela_buffer_801 (
        .din(new_Jinkela_wire_1383),
        .dout(new_Jinkela_wire_1384)
    );

    bfr new_Jinkela_buffer_1696 (
        .din(new_Jinkela_wire_2718),
        .dout(new_Jinkela_wire_2719)
    );

    bfr new_Jinkela_buffer_1420 (
        .din(new_Jinkela_wire_2267),
        .dout(new_Jinkela_wire_2268)
    );

    bfr new_Jinkela_buffer_1676 (
        .din(new_Jinkela_wire_2693),
        .dout(new_Jinkela_wire_2694)
    );

    bfr new_Jinkela_buffer_1375 (
        .din(new_Jinkela_wire_2222),
        .dout(new_Jinkela_wire_2223)
    );

    bfr new_Jinkela_buffer_802 (
        .din(new_Jinkela_wire_1384),
        .dout(new_Jinkela_wire_1385)
    );

    bfr new_Jinkela_buffer_1706 (
        .din(_0056_),
        .dout(new_Jinkela_wire_2731)
    );

    spl2 new_Jinkela_splitter_333 (
        .a(_0565_),
        .b(new_Jinkela_wire_2279),
        .c(new_Jinkela_wire_2280)
    );

    bfr new_Jinkela_buffer_841 (
        .din(_0721_),
        .dout(new_Jinkela_wire_1436)
    );

    bfr new_Jinkela_buffer_1677 (
        .din(new_Jinkela_wire_2694),
        .dout(new_Jinkela_wire_2695)
    );

    bfr new_Jinkela_buffer_1376 (
        .din(new_Jinkela_wire_2223),
        .dout(new_Jinkela_wire_2224)
    );

    bfr new_Jinkela_buffer_821 (
        .din(new_Jinkela_wire_1410),
        .dout(new_Jinkela_wire_1411)
    );

    bfr new_Jinkela_buffer_803 (
        .din(new_Jinkela_wire_1385),
        .dout(new_Jinkela_wire_1386)
    );

    bfr new_Jinkela_buffer_1697 (
        .din(new_Jinkela_wire_2719),
        .dout(new_Jinkela_wire_2720)
    );

    bfr new_Jinkela_buffer_1421 (
        .din(new_Jinkela_wire_2268),
        .dout(new_Jinkela_wire_2269)
    );

    bfr new_Jinkela_buffer_1678 (
        .din(new_Jinkela_wire_2695),
        .dout(new_Jinkela_wire_2696)
    );

    bfr new_Jinkela_buffer_1377 (
        .din(new_Jinkela_wire_2224),
        .dout(new_Jinkela_wire_2225)
    );

    bfr new_Jinkela_buffer_824 (
        .din(new_Jinkela_wire_1415),
        .dout(new_Jinkela_wire_1416)
    );

    bfr new_Jinkela_buffer_804 (
        .din(new_Jinkela_wire_1386),
        .dout(new_Jinkela_wire_1387)
    );

    bfr new_Jinkela_buffer_1703 (
        .din(new_Jinkela_wire_2727),
        .dout(new_Jinkela_wire_2728)
    );

    bfr new_Jinkela_buffer_842 (
        .din(new_Jinkela_wire_1436),
        .dout(new_Jinkela_wire_1437)
    );

    spl3L new_Jinkela_splitter_334 (
        .a(_0113_),
        .d(new_Jinkela_wire_2283),
        .b(new_Jinkela_wire_2284),
        .c(new_Jinkela_wire_2285)
    );

    bfr new_Jinkela_buffer_1679 (
        .din(new_Jinkela_wire_2696),
        .dout(new_Jinkela_wire_2697)
    );

    bfr new_Jinkela_buffer_1378 (
        .din(new_Jinkela_wire_2225),
        .dout(new_Jinkela_wire_2226)
    );

    bfr new_Jinkela_buffer_822 (
        .din(new_Jinkela_wire_1411),
        .dout(new_Jinkela_wire_1412)
    );

    bfr new_Jinkela_buffer_805 (
        .din(new_Jinkela_wire_1387),
        .dout(new_Jinkela_wire_1388)
    );

    bfr new_Jinkela_buffer_1705 (
        .din(new_Jinkela_wire_2729),
        .dout(new_Jinkela_wire_2730)
    );

    spl2 new_Jinkela_splitter_330 (
        .a(new_Jinkela_wire_2269),
        .b(new_Jinkela_wire_2270),
        .c(new_Jinkela_wire_2271)
    );

    bfr new_Jinkela_buffer_1680 (
        .din(new_Jinkela_wire_2697),
        .dout(new_Jinkela_wire_2698)
    );

    bfr new_Jinkela_buffer_1379 (
        .din(new_Jinkela_wire_2226),
        .dout(new_Jinkela_wire_2227)
    );

    bfr new_Jinkela_buffer_806 (
        .din(new_Jinkela_wire_1388),
        .dout(new_Jinkela_wire_1389)
    );

    bfr new_Jinkela_buffer_1709 (
        .din(_0440_),
        .dout(new_Jinkela_wire_2734)
    );

    bfr new_Jinkela_buffer_1422 (
        .din(new_Jinkela_wire_2271),
        .dout(new_Jinkela_wire_2272)
    );

    bfr new_Jinkela_buffer_1681 (
        .din(new_Jinkela_wire_2698),
        .dout(new_Jinkela_wire_2699)
    );

    bfr new_Jinkela_buffer_1380 (
        .din(new_Jinkela_wire_2227),
        .dout(new_Jinkela_wire_2228)
    );

    spl3L new_Jinkela_splitter_229 (
        .a(new_Jinkela_wire_1416),
        .d(new_Jinkela_wire_1417),
        .b(new_Jinkela_wire_1418),
        .c(new_Jinkela_wire_1419)
    );

    bfr new_Jinkela_buffer_807 (
        .din(new_Jinkela_wire_1389),
        .dout(new_Jinkela_wire_1390)
    );

    bfr new_Jinkela_buffer_1707 (
        .din(new_Jinkela_wire_2731),
        .dout(new_Jinkela_wire_2732)
    );

    spl2 new_Jinkela_splitter_232 (
        .a(_0048_),
        .b(new_Jinkela_wire_1463),
        .c(new_Jinkela_wire_1464)
    );

    bfr new_Jinkela_buffer_1424 (
        .din(new_Jinkela_wire_2280),
        .dout(new_Jinkela_wire_2281)
    );

    bfr new_Jinkela_buffer_1682 (
        .din(new_Jinkela_wire_2699),
        .dout(new_Jinkela_wire_2700)
    );

    bfr new_Jinkela_buffer_1381 (
        .din(new_Jinkela_wire_2228),
        .dout(new_Jinkela_wire_2229)
    );

    bfr new_Jinkela_buffer_808 (
        .din(new_Jinkela_wire_1390),
        .dout(new_Jinkela_wire_1391)
    );

    spl3L new_Jinkela_splitter_397 (
        .a(_0322_),
        .d(new_Jinkela_wire_2735),
        .b(new_Jinkela_wire_2736),
        .c(new_Jinkela_wire_2737)
    );

    bfr new_Jinkela_buffer_1711 (
        .din(_0476_),
        .dout(new_Jinkela_wire_2739)
    );

    bfr new_Jinkela_buffer_1426 (
        .din(_0208_),
        .dout(new_Jinkela_wire_2286)
    );

    bfr new_Jinkela_buffer_1683 (
        .din(new_Jinkela_wire_2700),
        .dout(new_Jinkela_wire_2701)
    );

    bfr new_Jinkela_buffer_1382 (
        .din(new_Jinkela_wire_2229),
        .dout(new_Jinkela_wire_2230)
    );

    bfr new_Jinkela_buffer_825 (
        .din(new_Jinkela_wire_1419),
        .dout(new_Jinkela_wire_1420)
    );

    bfr new_Jinkela_buffer_809 (
        .din(new_Jinkela_wire_1391),
        .dout(new_Jinkela_wire_1392)
    );

    bfr new_Jinkela_buffer_1708 (
        .din(new_Jinkela_wire_2732),
        .dout(new_Jinkela_wire_2733)
    );

    bfr new_Jinkela_buffer_1427 (
        .din(new_net_0),
        .dout(new_Jinkela_wire_2287)
    );

    bfr new_Jinkela_buffer_1438 (
        .din(_0477_),
        .dout(new_Jinkela_wire_2301)
    );

    bfr new_Jinkela_buffer_1684 (
        .din(new_Jinkela_wire_2701),
        .dout(new_Jinkela_wire_2702)
    );

    bfr new_Jinkela_buffer_1383 (
        .din(new_Jinkela_wire_2230),
        .dout(new_Jinkela_wire_2231)
    );

    bfr new_Jinkela_buffer_810 (
        .din(new_Jinkela_wire_1392),
        .dout(new_Jinkela_wire_1393)
    );

    bfr new_Jinkela_buffer_1712 (
        .din(_0489_),
        .dout(new_Jinkela_wire_2740)
    );

    bfr new_Jinkela_buffer_1425 (
        .din(new_Jinkela_wire_2281),
        .dout(new_Jinkela_wire_2282)
    );

    bfr new_Jinkela_buffer_843 (
        .din(new_Jinkela_wire_1437),
        .dout(new_Jinkela_wire_1438)
    );

    bfr new_Jinkela_buffer_1685 (
        .din(new_Jinkela_wire_2702),
        .dout(new_Jinkela_wire_2703)
    );

    bfr new_Jinkela_buffer_1384 (
        .din(new_Jinkela_wire_2231),
        .dout(new_Jinkela_wire_2232)
    );

    bfr new_Jinkela_buffer_826 (
        .din(new_Jinkela_wire_1420),
        .dout(new_Jinkela_wire_1421)
    );

    bfr new_Jinkela_buffer_811 (
        .din(new_Jinkela_wire_1393),
        .dout(new_Jinkela_wire_1394)
    );

    bfr new_Jinkela_buffer_1710 (
        .din(new_Jinkela_wire_2737),
        .dout(new_Jinkela_wire_2738)
    );

    bfr new_Jinkela_buffer_1719 (
        .din(_0761_),
        .dout(new_Jinkela_wire_2749)
    );

    bfr new_Jinkela_buffer_1686 (
        .din(new_Jinkela_wire_2703),
        .dout(new_Jinkela_wire_2704)
    );

    bfr new_Jinkela_buffer_1385 (
        .din(new_Jinkela_wire_2232),
        .dout(new_Jinkela_wire_2233)
    );

    bfr new_Jinkela_buffer_812 (
        .din(new_Jinkela_wire_1394),
        .dout(new_Jinkela_wire_1395)
    );

    spl3L new_Jinkela_splitter_336 (
        .a(_0200_),
        .d(new_Jinkela_wire_2302),
        .b(new_Jinkela_wire_2303),
        .c(new_Jinkela_wire_2304)
    );

    bfr new_Jinkela_buffer_1714 (
        .din(new_Jinkela_wire_2741),
        .dout(new_Jinkela_wire_2742)
    );

    bfr new_Jinkela_buffer_1386 (
        .din(new_Jinkela_wire_2233),
        .dout(new_Jinkela_wire_2234)
    );

    bfr new_Jinkela_buffer_827 (
        .din(new_Jinkela_wire_1421),
        .dout(new_Jinkela_wire_1422)
    );

    bfr new_Jinkela_buffer_813 (
        .din(new_Jinkela_wire_1395),
        .dout(new_Jinkela_wire_1396)
    );

    bfr new_Jinkela_buffer_1722 (
        .din(new_net_1469),
        .dout(new_Jinkela_wire_2752)
    );

    bfr new_Jinkela_buffer_1713 (
        .din(new_Jinkela_wire_2740),
        .dout(new_Jinkela_wire_2741)
    );

    bfr new_Jinkela_buffer_1387 (
        .din(new_Jinkela_wire_2234),
        .dout(new_Jinkela_wire_2235)
    );

    spl2 new_Jinkela_splitter_233 (
        .a(new_Jinkela_wire_1464),
        .b(new_Jinkela_wire_1465),
        .c(new_Jinkela_wire_1466)
    );

    bfr new_Jinkela_buffer_844 (
        .din(new_Jinkela_wire_1440),
        .dout(new_Jinkela_wire_1441)
    );

    bfr new_Jinkela_buffer_1720 (
        .din(new_Jinkela_wire_2749),
        .dout(new_Jinkela_wire_2750)
    );

    spl4L new_Jinkela_splitter_337 (
        .a(_0795_),
        .d(new_Jinkela_wire_2305),
        .e(new_Jinkela_wire_2306),
        .b(new_Jinkela_wire_2307),
        .c(new_Jinkela_wire_2308)
    );

    bfr new_Jinkela_buffer_828 (
        .din(new_Jinkela_wire_1422),
        .dout(new_Jinkela_wire_1423)
    );

    spl3L new_Jinkela_splitter_335 (
        .a(new_Jinkela_wire_2287),
        .d(new_Jinkela_wire_2288),
        .b(new_Jinkela_wire_2289),
        .c(new_Jinkela_wire_2290)
    );

    bfr new_Jinkela_buffer_1388 (
        .din(new_Jinkela_wire_2235),
        .dout(new_Jinkela_wire_2236)
    );

    bfr new_Jinkela_buffer_864 (
        .din(_0475_),
        .dout(new_Jinkela_wire_1467)
    );

    bfr new_Jinkela_buffer_1724 (
        .din(_0723_),
        .dout(new_Jinkela_wire_2754)
    );

    or_bb _1373_ (
        .a(new_Jinkela_wire_1073),
        .b(_0506_),
        .c(new_net_2)
    );

    or_bb _1374_ (
        .a(new_Jinkela_wire_2900),
        .b(new_Jinkela_wire_3271),
        .c(_0541_)
    );

    or_bb _1375_ (
        .a(new_Jinkela_wire_2972),
        .b(new_Jinkela_wire_1155),
        .c(_0542_)
    );

    and_bi _1376_ (
        .a(new_Jinkela_wire_2833),
        .b(new_Jinkela_wire_2651),
        .c(_0543_)
    );

    and_bi _1377_ (
        .a(new_Jinkela_wire_2650),
        .b(new_Jinkela_wire_2832),
        .c(_0544_)
    );

    or_bb _1378_ (
        .a(_0544_),
        .b(_0543_),
        .c(_0545_)
    );

    and_ii _1379_ (
        .a(new_Jinkela_wire_2971),
        .b(new_Jinkela_wire_1891),
        .c(_0546_)
    );

    or_bb _1380_ (
        .a(new_Jinkela_wire_1934),
        .b(new_Jinkela_wire_1146),
        .c(_0547_)
    );

    and_bb _1381_ (
        .a(new_Jinkela_wire_1933),
        .b(new_Jinkela_wire_1145),
        .c(_0548_)
    );

    and_bi _1382_ (
        .a(_0547_),
        .b(_0548_),
        .c(_0549_)
    );

    or_ii _1383_ (
        .a(new_Jinkela_wire_2061),
        .b(new_Jinkela_wire_26),
        .c(_0550_)
    );

    and_bi _1384_ (
        .a(new_Jinkela_wire_3203),
        .b(_0550_),
        .c(new_net_4)
    );

    and_ii _1385_ (
        .a(new_Jinkela_wire_2970),
        .b(new_Jinkela_wire_2173),
        .c(_0551_)
    );

    or_bi _1386_ (
        .a(new_Jinkela_wire_1624),
        .b(new_Jinkela_wire_908),
        .c(_0552_)
    );

    and_bi _1387_ (
        .a(new_Jinkela_wire_1623),
        .b(new_Jinkela_wire_907),
        .c(_0553_)
    );

    or_bi _1388_ (
        .a(_0553_),
        .b(_0552_),
        .c(_0554_)
    );

    and_bi _1389_ (
        .a(new_Jinkela_wire_2978),
        .b(new_Jinkela_wire_1752),
        .c(_0555_)
    );

    or_bi _1390_ (
        .a(new_Jinkela_wire_3041),
        .b(new_Jinkela_wire_3201),
        .c(_0556_)
    );

    and_bi _1391_ (
        .a(new_Jinkela_wire_2979),
        .b(new_Jinkela_wire_1407),
        .c(_0557_)
    );

    and_bi _1392_ (
        .a(new_Jinkela_wire_1531),
        .b(new_Jinkela_wire_897),
        .c(_0558_)
    );

    and_bi _1393_ (
        .a(new_Jinkela_wire_1529),
        .b(new_Jinkela_wire_2013),
        .c(_0559_)
    );

    and_bi _1394_ (
        .a(new_Jinkela_wire_2012),
        .b(new_Jinkela_wire_1528),
        .c(_0560_)
    );

    and_ii _1395_ (
        .a(new_Jinkela_wire_2957),
        .b(new_Jinkela_wire_2004),
        .c(_0561_)
    );

    and_bi _1396_ (
        .a(new_Jinkela_wire_2278),
        .b(new_Jinkela_wire_2467),
        .c(_0562_)
    );

    and_bi _1397_ (
        .a(new_Jinkela_wire_2468),
        .b(new_Jinkela_wire_2277),
        .c(_0563_)
    );

    or_bb _1398_ (
        .a(new_Jinkela_wire_2571),
        .b(new_Jinkela_wire_3215),
        .c(_0564_)
    );

    and_bi _1399_ (
        .a(new_Jinkela_wire_25),
        .b(new_Jinkela_wire_2062),
        .c(_0565_)
    );

    inv _1400_ (
        .din(new_Jinkela_wire_2279),
        .dout(_0566_)
    );

    and_bb _1401_ (
        .a(new_Jinkela_wire_3037),
        .b(new_Jinkela_wire_2652),
        .c(_0567_)
    );

    or_bi _1402_ (
        .a(new_Jinkela_wire_3207),
        .b(new_Jinkela_wire_1530),
        .c(_0568_)
    );

    or_ii _1403_ (
        .a(new_Jinkela_wire_1642),
        .b(new_Jinkela_wire_2783),
        .c(_0569_)
    );

    and_bi _1404_ (
        .a(new_Jinkela_wire_2282),
        .b(new_Jinkela_wire_1641),
        .c(_0570_)
    );

    and_bi _1405_ (
        .a(_0569_),
        .b(_0570_),
        .c(_0571_)
    );

    or_bb _1406_ (
        .a(new_Jinkela_wire_830),
        .b(new_Jinkela_wire_2892),
        .c(_0572_)
    );

    or_ii _1407_ (
        .a(new_Jinkela_wire_1484),
        .b(new_Jinkela_wire_1553),
        .c(_0573_)
    );

    and_ii _1408_ (
        .a(new_Jinkela_wire_1680),
        .b(new_Jinkela_wire_1734),
        .c(_0574_)
    );

    or_bb _1409_ (
        .a(new_Jinkela_wire_3334),
        .b(new_Jinkela_wire_803),
        .c(_0575_)
    );

    or_bb _1410_ (
        .a(new_Jinkela_wire_1663),
        .b(new_Jinkela_wire_1523),
        .c(_0576_)
    );

    and_bi _1411_ (
        .a(new_Jinkela_wire_502),
        .b(new_Jinkela_wire_2364),
        .c(_0577_)
    );

    and_bi _1412_ (
        .a(new_Jinkela_wire_1064),
        .b(new_Jinkela_wire_1124),
        .c(_0578_)
    );

    or_ii _1413_ (
        .a(new_Jinkela_wire_571),
        .b(new_Jinkela_wire_330),
        .c(_0579_)
    );

    and_bi _1414_ (
        .a(new_Jinkela_wire_3024),
        .b(new_Jinkela_wire_2419),
        .c(_0580_)
    );

    bfr new_Jinkela_buffer_939 (
        .din(new_Jinkela_wire_1583),
        .dout(new_Jinkela_wire_1584)
    );

    bfr new_Jinkela_buffer_919 (
        .din(new_Jinkela_wire_1557),
        .dout(new_Jinkela_wire_1558)
    );

    bfr new_Jinkela_buffer_920 (
        .din(new_Jinkela_wire_1558),
        .dout(new_Jinkela_wire_1559)
    );

    bfr new_Jinkela_buffer_940 (
        .din(new_Jinkela_wire_1584),
        .dout(new_Jinkela_wire_1585)
    );

    spl2 new_Jinkela_splitter_250 (
        .a(new_Jinkela_wire_1559),
        .b(new_Jinkela_wire_1560),
        .c(new_Jinkela_wire_1561)
    );

    bfr new_Jinkela_buffer_921 (
        .din(new_Jinkela_wire_1561),
        .dout(new_Jinkela_wire_1562)
    );

    bfr new_Jinkela_buffer_979 (
        .din(new_Jinkela_wire_1631),
        .dout(new_Jinkela_wire_1632)
    );

    bfr new_Jinkela_buffer_941 (
        .din(new_Jinkela_wire_1585),
        .dout(new_Jinkela_wire_1586)
    );

    bfr new_Jinkela_buffer_922 (
        .din(new_Jinkela_wire_1562),
        .dout(new_Jinkela_wire_1563)
    );

    spl2 new_Jinkela_splitter_258 (
        .a(_0277_),
        .b(new_Jinkela_wire_1645),
        .c(new_Jinkela_wire_1646)
    );

    spl2 new_Jinkela_splitter_257 (
        .a(_0473_),
        .b(new_Jinkela_wire_1643),
        .c(new_Jinkela_wire_1644)
    );

    spl2 new_Jinkela_splitter_251 (
        .a(new_Jinkela_wire_1563),
        .b(new_Jinkela_wire_1564),
        .c(new_Jinkela_wire_1565)
    );

    bfr new_Jinkela_buffer_980 (
        .din(new_Jinkela_wire_1632),
        .dout(new_Jinkela_wire_1633)
    );

    bfr new_Jinkela_buffer_942 (
        .din(new_Jinkela_wire_1586),
        .dout(new_Jinkela_wire_1587)
    );

    bfr new_Jinkela_buffer_943 (
        .din(new_Jinkela_wire_1587),
        .dout(new_Jinkela_wire_1588)
    );

    bfr new_Jinkela_buffer_944 (
        .din(new_Jinkela_wire_1588),
        .dout(new_Jinkela_wire_1589)
    );

    bfr new_Jinkela_buffer_992 (
        .din(_0575_),
        .dout(new_Jinkela_wire_1651)
    );

    bfr new_Jinkela_buffer_981 (
        .din(new_Jinkela_wire_1633),
        .dout(new_Jinkela_wire_1634)
    );

    bfr new_Jinkela_buffer_945 (
        .din(new_Jinkela_wire_1589),
        .dout(new_Jinkela_wire_1590)
    );

    bfr new_Jinkela_buffer_988 (
        .din(_0689_),
        .dout(new_Jinkela_wire_1647)
    );

    bfr new_Jinkela_buffer_946 (
        .din(new_Jinkela_wire_1590),
        .dout(new_Jinkela_wire_1591)
    );

    bfr new_Jinkela_buffer_982 (
        .din(new_Jinkela_wire_1634),
        .dout(new_Jinkela_wire_1635)
    );

    bfr new_Jinkela_buffer_947 (
        .din(new_Jinkela_wire_1591),
        .dout(new_Jinkela_wire_1592)
    );

    bfr new_Jinkela_buffer_948 (
        .din(new_Jinkela_wire_1592),
        .dout(new_Jinkela_wire_1593)
    );

    bfr new_Jinkela_buffer_989 (
        .din(_0599_),
        .dout(new_Jinkela_wire_1648)
    );

    bfr new_Jinkela_buffer_983 (
        .din(new_Jinkela_wire_1635),
        .dout(new_Jinkela_wire_1636)
    );

    bfr new_Jinkela_buffer_949 (
        .din(new_Jinkela_wire_1593),
        .dout(new_Jinkela_wire_1594)
    );

    spl3L new_Jinkela_splitter_260 (
        .a(_0740_),
        .d(new_Jinkela_wire_1667),
        .b(new_Jinkela_wire_1668),
        .c(new_Jinkela_wire_1669)
    );

    bfr new_Jinkela_buffer_950 (
        .din(new_Jinkela_wire_1594),
        .dout(new_Jinkela_wire_1595)
    );

    bfr new_Jinkela_buffer_990 (
        .din(new_Jinkela_wire_1648),
        .dout(new_Jinkela_wire_1649)
    );

    bfr new_Jinkela_buffer_984 (
        .din(new_Jinkela_wire_1636),
        .dout(new_Jinkela_wire_1637)
    );

    bfr new_Jinkela_buffer_951 (
        .din(new_Jinkela_wire_1595),
        .dout(new_Jinkela_wire_1596)
    );

    bfr new_Jinkela_buffer_952 (
        .din(new_Jinkela_wire_1596),
        .dout(new_Jinkela_wire_1597)
    );

    bfr new_Jinkela_buffer_985 (
        .din(new_Jinkela_wire_1637),
        .dout(new_Jinkela_wire_1638)
    );

    bfr new_Jinkela_buffer_953 (
        .din(new_Jinkela_wire_1597),
        .dout(new_Jinkela_wire_1598)
    );

    spl2 new_Jinkela_splitter_262 (
        .a(_0039_),
        .b(new_Jinkela_wire_1673),
        .c(new_Jinkela_wire_1674)
    );

    bfr new_Jinkela_buffer_954 (
        .din(new_Jinkela_wire_1598),
        .dout(new_Jinkela_wire_1599)
    );

    bfr new_Jinkela_buffer_991 (
        .din(new_Jinkela_wire_1649),
        .dout(new_Jinkela_wire_1650)
    );

    bfr new_Jinkela_buffer_986 (
        .din(new_Jinkela_wire_1638),
        .dout(new_Jinkela_wire_1639)
    );

    bfr new_Jinkela_buffer_955 (
        .din(new_Jinkela_wire_1599),
        .dout(new_Jinkela_wire_1600)
    );

    bfr new_Jinkela_buffer_956 (
        .din(new_Jinkela_wire_1600),
        .dout(new_Jinkela_wire_1601)
    );

    bfr new_Jinkela_buffer_1005 (
        .din(_0105_),
        .dout(new_Jinkela_wire_1675)
    );

    bfr new_Jinkela_buffer_1428 (
        .din(new_Jinkela_wire_2290),
        .dout(new_Jinkela_wire_2291)
    );

    bfr new_Jinkela_buffer_1715 (
        .din(new_Jinkela_wire_2742),
        .dout(new_Jinkela_wire_2743)
    );

    and_bi _1037_ (
        .a(new_Jinkela_wire_2638),
        .b(new_Jinkela_wire_2286),
        .c(_0209_)
    );

    bfr new_Jinkela_buffer_758 (
        .din(new_Jinkela_wire_1317),
        .dout(new_Jinkela_wire_1318)
    );

    bfr new_Jinkela_buffer_1389 (
        .din(new_Jinkela_wire_2236),
        .dout(new_Jinkela_wire_2237)
    );

    and_bi _1038_ (
        .a(new_Jinkela_wire_1034),
        .b(_0209_),
        .c(_0210_)
    );

    bfr new_Jinkela_buffer_771 (
        .din(new_Jinkela_wire_1332),
        .dout(new_Jinkela_wire_1333)
    );

    bfr new_Jinkela_buffer_1721 (
        .din(new_Jinkela_wire_2750),
        .dout(new_Jinkela_wire_2751)
    );

    bfr new_Jinkela_buffer_1716 (
        .din(new_Jinkela_wire_2743),
        .dout(new_Jinkela_wire_2744)
    );

    or_bb _1039_ (
        .a(new_Jinkela_wire_2211),
        .b(_0206_),
        .c(_0211_)
    );

    bfr new_Jinkela_buffer_759 (
        .din(new_Jinkela_wire_1318),
        .dout(new_Jinkela_wire_1319)
    );

    spl2 new_Jinkela_splitter_338 (
        .a(_0167_),
        .b(new_Jinkela_wire_2310),
        .c(new_Jinkela_wire_2311)
    );

    bfr new_Jinkela_buffer_1390 (
        .din(new_Jinkela_wire_2237),
        .dout(new_Jinkela_wire_2238)
    );

    and_bi _1040_ (
        .a(_0203_),
        .b(new_Jinkela_wire_1620),
        .c(_0212_)
    );

    bfr new_Jinkela_buffer_1723 (
        .din(new_Jinkela_wire_2752),
        .dout(new_Jinkela_wire_2753)
    );

    spl2 new_Jinkela_splitter_220 (
        .a(_0030_),
        .b(new_Jinkela_wire_1352),
        .c(new_Jinkela_wire_1353)
    );

    bfr new_Jinkela_buffer_1429 (
        .din(new_Jinkela_wire_2291),
        .dout(new_Jinkela_wire_2292)
    );

    bfr new_Jinkela_buffer_1717 (
        .din(new_Jinkela_wire_2744),
        .dout(new_Jinkela_wire_2745)
    );

    or_bb _1041_ (
        .a(new_Jinkela_wire_2381),
        .b(new_Jinkela_wire_540),
        .c(_0213_)
    );

    bfr new_Jinkela_buffer_760 (
        .din(new_Jinkela_wire_1319),
        .dout(new_Jinkela_wire_1320)
    );

    bfr new_Jinkela_buffer_1391 (
        .din(new_Jinkela_wire_2238),
        .dout(new_Jinkela_wire_2239)
    );

    and_ii _1042_ (
        .a(new_Jinkela_wire_2182),
        .b(new_Jinkela_wire_2165),
        .c(_0214_)
    );

    bfr new_Jinkela_buffer_1725 (
        .din(_0729_),
        .dout(new_Jinkela_wire_2755)
    );

    bfr new_Jinkela_buffer_1444 (
        .din(_0137_),
        .dout(new_Jinkela_wire_2322)
    );

    spl2 new_Jinkela_splitter_221 (
        .a(_0268_),
        .b(new_Jinkela_wire_1354),
        .c(new_Jinkela_wire_1355)
    );

    spl2 new_Jinkela_splitter_398 (
        .a(new_Jinkela_wire_2745),
        .b(new_Jinkela_wire_2746),
        .c(new_Jinkela_wire_2747)
    );

    or_ii _1043_ (
        .a(new_Jinkela_wire_2176),
        .b(new_Jinkela_wire_484),
        .c(_0215_)
    );

    bfr new_Jinkela_buffer_761 (
        .din(new_Jinkela_wire_1320),
        .dout(new_Jinkela_wire_1321)
    );

    spl2 new_Jinkela_splitter_341 (
        .a(_0304_),
        .b(new_Jinkela_wire_2318),
        .c(new_Jinkela_wire_2319)
    );

    bfr new_Jinkela_buffer_1392 (
        .din(new_Jinkela_wire_2239),
        .dout(new_Jinkela_wire_2240)
    );

    bfr new_Jinkela_buffer_1718 (
        .din(new_Jinkela_wire_2747),
        .dout(new_Jinkela_wire_2748)
    );

    and_bi _1044_ (
        .a(new_Jinkela_wire_776),
        .b(new_Jinkela_wire_3029),
        .c(_0216_)
    );

    bfr new_Jinkela_buffer_779 (
        .din(new_Jinkela_wire_1350),
        .dout(new_Jinkela_wire_1351)
    );

    bfr new_Jinkela_buffer_1430 (
        .din(new_Jinkela_wire_2292),
        .dout(new_Jinkela_wire_2293)
    );

    bfr new_Jinkela_buffer_773 (
        .din(new_Jinkela_wire_1334),
        .dout(new_Jinkela_wire_1335)
    );

    or_bb _1045_ (
        .a(new_Jinkela_wire_237),
        .b(new_Jinkela_wire_438),
        .c(_0217_)
    );

    bfr new_Jinkela_buffer_762 (
        .din(new_Jinkela_wire_1321),
        .dout(new_Jinkela_wire_1322)
    );

    bfr new_Jinkela_buffer_1727 (
        .din(_0116_),
        .dout(new_Jinkela_wire_2757)
    );

    bfr new_Jinkela_buffer_1393 (
        .din(new_Jinkela_wire_2240),
        .dout(new_Jinkela_wire_2241)
    );

    and_bi _1046_ (
        .a(new_Jinkela_wire_422),
        .b(new_Jinkela_wire_259),
        .c(_0218_)
    );

    bfr new_Jinkela_buffer_774 (
        .din(new_Jinkela_wire_1335),
        .dout(new_Jinkela_wire_1336)
    );

    bfr new_Jinkela_buffer_1726 (
        .din(new_Jinkela_wire_2755),
        .dout(new_Jinkela_wire_2756)
    );

    and_bi _1047_ (
        .a(_0217_),
        .b(new_Jinkela_wire_3128),
        .c(_0219_)
    );

    bfr new_Jinkela_buffer_763 (
        .din(new_Jinkela_wire_1322),
        .dout(new_Jinkela_wire_1323)
    );

    spl2 new_Jinkela_splitter_340 (
        .a(_0436_),
        .b(new_Jinkela_wire_2316),
        .c(new_Jinkela_wire_2317)
    );

    bfr new_Jinkela_buffer_1394 (
        .din(new_Jinkela_wire_2241),
        .dout(new_Jinkela_wire_2242)
    );

    spl2 new_Jinkela_splitter_402 (
        .a(_0027_),
        .b(new_Jinkela_wire_2777),
        .c(new_Jinkela_wire_2778)
    );

    or_bb _1048_ (
        .a(new_Jinkela_wire_2320),
        .b(_0216_),
        .c(_0220_)
    );

    bfr new_Jinkela_buffer_1728 (
        .din(new_Jinkela_wire_2757),
        .dout(new_Jinkela_wire_2758)
    );

    bfr new_Jinkela_buffer_780 (
        .din(_0574_),
        .dout(new_Jinkela_wire_1356)
    );

    bfr new_Jinkela_buffer_1431 (
        .din(new_Jinkela_wire_2293),
        .dout(new_Jinkela_wire_2294)
    );

    and_bi _1049_ (
        .a(new_Jinkela_wire_1273),
        .b(_0220_),
        .c(_0221_)
    );

    bfr new_Jinkela_buffer_784 (
        .din(_0585_),
        .dout(new_Jinkela_wire_1367)
    );

    bfr new_Jinkela_buffer_1395 (
        .din(new_Jinkela_wire_2242),
        .dout(new_Jinkela_wire_2243)
    );

    bfr new_Jinkela_buffer_775 (
        .din(new_Jinkela_wire_1336),
        .dout(new_Jinkela_wire_1337)
    );

    bfr new_Jinkela_buffer_1737 (
        .din(_0513_),
        .dout(new_Jinkela_wire_2772)
    );

    and_bi _1050_ (
        .a(new_Jinkela_wire_1043),
        .b(_0221_),
        .c(_0222_)
    );

    bfr new_Jinkela_buffer_1729 (
        .din(new_Jinkela_wire_2758),
        .dout(new_Jinkela_wire_2759)
    );

    bfr new_Jinkela_buffer_1439 (
        .din(new_Jinkela_wire_2308),
        .dout(new_Jinkela_wire_2309)
    );

    or_bb _1051_ (
        .a(new_Jinkela_wire_2265),
        .b(new_Jinkela_wire_962),
        .c(_0223_)
    );

    bfr new_Jinkela_buffer_1735 (
        .din(_0487_),
        .dout(new_Jinkela_wire_2770)
    );

    bfr new_Jinkela_buffer_1396 (
        .din(new_Jinkela_wire_2243),
        .dout(new_Jinkela_wire_2244)
    );

    bfr new_Jinkela_buffer_781 (
        .din(_0316_),
        .dout(new_Jinkela_wire_1359)
    );

    or_bb _1052_ (
        .a(new_Jinkela_wire_2584),
        .b(new_Jinkela_wire_3064),
        .c(_0224_)
    );

    bfr new_Jinkela_buffer_1736 (
        .din(new_Jinkela_wire_2770),
        .dout(new_Jinkela_wire_2771)
    );

    spl2 new_Jinkela_splitter_217 (
        .a(new_Jinkela_wire_1337),
        .b(new_Jinkela_wire_1338),
        .c(new_Jinkela_wire_1340)
    );

    bfr new_Jinkela_buffer_1432 (
        .din(new_Jinkela_wire_2294),
        .dout(new_Jinkela_wire_2295)
    );

    and_ii _1053_ (
        .a(_0224_),
        .b(new_Jinkela_wire_2171),
        .c(_0225_)
    );

    spl2 new_Jinkela_splitter_399 (
        .a(new_Jinkela_wire_2759),
        .b(new_Jinkela_wire_2760),
        .c(new_Jinkela_wire_2761)
    );

    spl4L new_Jinkela_splitter_218 (
        .a(new_Jinkela_wire_1340),
        .d(new_Jinkela_wire_1341),
        .e(new_Jinkela_wire_1342),
        .b(new_Jinkela_wire_1343),
        .c(new_Jinkela_wire_1345)
    );

    bfr new_Jinkela_buffer_1397 (
        .din(new_Jinkela_wire_2244),
        .dout(new_Jinkela_wire_2245)
    );

    spl3L new_Jinkela_splitter_403 (
        .a(new_Jinkela_wire_2778),
        .d(new_Jinkela_wire_2779),
        .b(new_Jinkela_wire_2780),
        .c(new_Jinkela_wire_2781)
    );

    and_bi _1054_ (
        .a(new_Jinkela_wire_2567),
        .b(new_Jinkela_wire_2585),
        .c(_0226_)
    );

    bfr new_Jinkela_buffer_1730 (
        .din(new_Jinkela_wire_2761),
        .dout(new_Jinkela_wire_2762)
    );

    bfr new_Jinkela_buffer_776 (
        .din(new_Jinkela_wire_1338),
        .dout(new_Jinkela_wire_1339)
    );

    and_bi _1055_ (
        .a(new_Jinkela_wire_2172),
        .b(_0226_),
        .c(_0227_)
    );

    bfr new_Jinkela_buffer_1440 (
        .din(new_Jinkela_wire_2311),
        .dout(new_Jinkela_wire_2312)
    );

    spl2 new_Jinkela_splitter_401 (
        .a(new_Jinkela_wire_2772),
        .b(new_Jinkela_wire_2773),
        .c(new_Jinkela_wire_2774)
    );

    bfr new_Jinkela_buffer_1398 (
        .din(new_Jinkela_wire_2245),
        .dout(new_Jinkela_wire_2246)
    );

    or_bb _1056_ (
        .a(new_Jinkela_wire_1767),
        .b(new_Jinkela_wire_1198),
        .c(_0228_)
    );

    spl2 new_Jinkela_splitter_222 (
        .a(_0362_),
        .b(new_Jinkela_wire_1357),
        .c(new_Jinkela_wire_1358)
    );

    bfr new_Jinkela_buffer_1738 (
        .din(new_Jinkela_wire_2774),
        .dout(new_Jinkela_wire_2775)
    );

    spl4L new_Jinkela_splitter_219 (
        .a(new_Jinkela_wire_1345),
        .d(new_Jinkela_wire_1346),
        .e(new_Jinkela_wire_1347),
        .b(new_Jinkela_wire_1348),
        .c(new_Jinkela_wire_1349)
    );

    bfr new_Jinkela_buffer_1433 (
        .din(new_Jinkela_wire_2295),
        .dout(new_Jinkela_wire_2296)
    );

    and_bi _1057_ (
        .a(new_Jinkela_wire_2302),
        .b(new_Jinkela_wire_906),
        .c(_0229_)
    );

    bfr new_Jinkela_buffer_1731 (
        .din(new_Jinkela_wire_2762),
        .dout(new_Jinkela_wire_2763)
    );

    bfr new_Jinkela_buffer_777 (
        .din(new_Jinkela_wire_1343),
        .dout(new_Jinkela_wire_1344)
    );

    bfr new_Jinkela_buffer_1399 (
        .din(new_Jinkela_wire_2246),
        .dout(new_Jinkela_wire_2247)
    );

    or_bb _1058_ (
        .a(new_Jinkela_wire_933),
        .b(new_Jinkela_wire_231),
        .c(_0230_)
    );

    bfr new_Jinkela_buffer_1740 (
        .din(_0393_),
        .dout(new_Jinkela_wire_2784)
    );

    and_bi _1059_ (
        .a(new_Jinkela_wire_229),
        .b(new_Jinkela_wire_2443),
        .c(_0231_)
    );

    spl3L new_Jinkela_splitter_400 (
        .a(new_Jinkela_wire_2763),
        .d(new_Jinkela_wire_2764),
        .b(new_Jinkela_wire_2765),
        .c(new_Jinkela_wire_2766)
    );

    bfr new_Jinkela_buffer_1400 (
        .din(new_Jinkela_wire_2247),
        .dout(new_Jinkela_wire_2248)
    );

    bfr new_Jinkela_buffer_782 (
        .din(new_Jinkela_wire_1359),
        .dout(new_Jinkela_wire_1360)
    );

    and_bb _1060_ (
        .a(new_Jinkela_wire_417),
        .b(new_Jinkela_wire_284),
        .c(_0232_)
    );

    bfr new_Jinkela_buffer_786 (
        .din(_0773_),
        .dout(new_Jinkela_wire_1369)
    );

    spl3L new_Jinkela_splitter_224 (
        .a(_0114_),
        .d(new_Jinkela_wire_1364),
        .b(new_Jinkela_wire_1365),
        .c(new_Jinkela_wire_1366)
    );

    bfr new_Jinkela_buffer_1434 (
        .din(new_Jinkela_wire_2296),
        .dout(new_Jinkela_wire_2297)
    );

    and_bi _1061_ (
        .a(new_Jinkela_wire_3176),
        .b(new_Jinkela_wire_2005),
        .c(_0233_)
    );

    bfr new_Jinkela_buffer_1732 (
        .din(new_Jinkela_wire_2766),
        .dout(new_Jinkela_wire_2767)
    );

    bfr new_Jinkela_buffer_1401 (
        .din(new_Jinkela_wire_2248),
        .dout(new_Jinkela_wire_2249)
    );

    and_bi _1062_ (
        .a(new_Jinkela_wire_1031),
        .b(_0233_),
        .c(_0234_)
    );

    spl2 new_Jinkela_splitter_404 (
        .a(_0566_),
        .b(new_Jinkela_wire_2782),
        .c(new_Jinkela_wire_2783)
    );

    bfr new_Jinkela_buffer_1739 (
        .din(new_Jinkela_wire_2775),
        .dout(new_Jinkela_wire_2776)
    );

    bfr new_Jinkela_buffer_783 (
        .din(new_Jinkela_wire_1360),
        .dout(new_Jinkela_wire_1361)
    );

    or_bb _1063_ (
        .a(new_Jinkela_wire_2017),
        .b(_0231_),
        .c(_0235_)
    );

    spl2 new_Jinkela_splitter_339 (
        .a(new_Jinkela_wire_2312),
        .b(new_Jinkela_wire_2313),
        .c(new_Jinkela_wire_2314)
    );

    bfr new_Jinkela_buffer_1733 (
        .din(new_Jinkela_wire_2767),
        .dout(new_Jinkela_wire_2768)
    );

    bfr new_Jinkela_buffer_1402 (
        .din(new_Jinkela_wire_2249),
        .dout(new_Jinkela_wire_2250)
    );

    and_bi _1064_ (
        .a(_0230_),
        .b(_0235_),
        .c(_0236_)
    );

    bfr new_Jinkela_buffer_785 (
        .din(new_Jinkela_wire_1367),
        .dout(new_Jinkela_wire_1368)
    );

    bfr new_Jinkela_buffer_1435 (
        .din(new_Jinkela_wire_2297),
        .dout(new_Jinkela_wire_2298)
    );

    spl2 new_Jinkela_splitter_223 (
        .a(new_Jinkela_wire_1361),
        .b(new_Jinkela_wire_1362),
        .c(new_Jinkela_wire_1363)
    );

    or_ii _1065_ (
        .a(new_Jinkela_wire_2178),
        .b(new_Jinkela_wire_518),
        .c(_0237_)
    );

    bfr new_Jinkela_buffer_1734 (
        .din(new_Jinkela_wire_2768),
        .dout(new_Jinkela_wire_2769)
    );

    bfr new_Jinkela_buffer_1403 (
        .din(new_Jinkela_wire_2250),
        .dout(new_Jinkela_wire_2251)
    );

    and_bb _1066_ (
        .a(new_Jinkela_wire_415),
        .b(new_Jinkela_wire_480),
        .c(_0238_)
    );

    bfr new_Jinkela_buffer_787 (
        .din(new_Jinkela_wire_1369),
        .dout(new_Jinkela_wire_1370)
    );

    bfr new_Jinkela_buffer_1743 (
        .din(_0259_),
        .dout(new_Jinkela_wire_2787)
    );

    and_bi _1067_ (
        .a(new_Jinkela_wire_717),
        .b(new_Jinkela_wire_424),
        .c(_0239_)
    );

    bfr new_Jinkela_buffer_789 (
        .din(new_net_1483),
        .dout(new_Jinkela_wire_1372)
    );

    bfr new_Jinkela_buffer_1441 (
        .din(new_Jinkela_wire_2314),
        .dout(new_Jinkela_wire_2315)
    );

    bfr new_Jinkela_buffer_1404 (
        .din(new_Jinkela_wire_2251),
        .dout(new_Jinkela_wire_2252)
    );

    bfr new_Jinkela_buffer_1741 (
        .din(new_Jinkela_wire_2784),
        .dout(new_Jinkela_wire_2785)
    );

    or_bb _1068_ (
        .a(_0239_),
        .b(_0238_),
        .c(_0240_)
    );

    bfr new_Jinkela_buffer_814 (
        .din(_0077_),
        .dout(new_Jinkela_wire_1397)
    );

    bfr new_Jinkela_buffer_1746 (
        .din(_0788_),
        .dout(new_Jinkela_wire_2790)
    );

    bfr new_Jinkela_buffer_1436 (
        .din(new_Jinkela_wire_2298),
        .dout(new_Jinkela_wire_2299)
    );

    and_bi _1069_ (
        .a(new_Jinkela_wire_263),
        .b(new_Jinkela_wire_3027),
        .c(_0241_)
    );

    bfr new_Jinkela_buffer_788 (
        .din(new_Jinkela_wire_1370),
        .dout(new_Jinkela_wire_1371)
    );

    bfr new_Jinkela_buffer_1742 (
        .din(new_Jinkela_wire_2785),
        .dout(new_Jinkela_wire_2786)
    );

    bfr new_Jinkela_buffer_1405 (
        .din(new_Jinkela_wire_2252),
        .dout(new_Jinkela_wire_2253)
    );

    or_bb _1070_ (
        .a(_0241_),
        .b(new_Jinkela_wire_1239),
        .c(_0242_)
    );

    bfr new_Jinkela_buffer_790 (
        .din(new_Jinkela_wire_1372),
        .dout(new_Jinkela_wire_1373)
    );

    bfr new_Jinkela_buffer_1744 (
        .din(new_Jinkela_wire_2787),
        .dout(new_Jinkela_wire_2788)
    );

    bfr new_Jinkela_buffer_1747 (
        .din(new_net_8),
        .dout(new_Jinkela_wire_2791)
    );

    and_bi _1071_ (
        .a(new_Jinkela_wire_2183),
        .b(_0242_),
        .c(_0243_)
    );

    bfr new_Jinkela_buffer_816 (
        .din(_0743_),
        .dout(new_Jinkela_wire_1399)
    );

    bfr new_Jinkela_buffer_1406 (
        .din(new_Jinkela_wire_2253),
        .dout(new_Jinkela_wire_2254)
    );

    bfr new_Jinkela_buffer_1442 (
        .din(_0219_),
        .dout(new_Jinkela_wire_2320)
    );

    bfr new_Jinkela_buffer_1774 (
        .din(_0712_),
        .dout(new_Jinkela_wire_2821)
    );

    and_bi _1072_ (
        .a(new_Jinkela_wire_1045),
        .b(_0243_),
        .c(_0244_)
    );

    bfr new_Jinkela_buffer_791 (
        .din(new_Jinkela_wire_1373),
        .dout(new_Jinkela_wire_1374)
    );

    bfr new_Jinkela_buffer_1745 (
        .din(new_Jinkela_wire_2788),
        .dout(new_Jinkela_wire_2789)
    );

    bfr new_Jinkela_buffer_1437 (
        .din(new_Jinkela_wire_2299),
        .dout(new_Jinkela_wire_2300)
    );

    or_bb _1073_ (
        .a(new_Jinkela_wire_2011),
        .b(new_Jinkela_wire_963),
        .c(_0245_)
    );

    bfr new_Jinkela_buffer_815 (
        .din(new_Jinkela_wire_1397),
        .dout(new_Jinkela_wire_1398)
    );

    bfr new_Jinkela_buffer_1749 (
        .din(new_Jinkela_wire_2792),
        .dout(new_Jinkela_wire_2793)
    );

    bfr new_Jinkela_buffer_1407 (
        .din(new_Jinkela_wire_2254),
        .dout(new_Jinkela_wire_2255)
    );

    or_bb _1074_ (
        .a(new_Jinkela_wire_1036),
        .b(new_Jinkela_wire_3059),
        .c(_0246_)
    );

    bfr new_Jinkela_buffer_792 (
        .din(new_Jinkela_wire_1374),
        .dout(new_Jinkela_wire_1375)
    );

    bfr new_Jinkela_buffer_1748 (
        .din(new_Jinkela_wire_2791),
        .dout(new_Jinkela_wire_2792)
    );

    or_bb _1075_ (
        .a(_0246_),
        .b(new_Jinkela_wire_1154),
        .c(_0247_)
    );

    spl2 new_Jinkela_splitter_225 (
        .a(_0191_),
        .b(new_Jinkela_wire_1400),
        .c(new_Jinkela_wire_1401)
    );

    bfr new_Jinkela_buffer_1443 (
        .din(_0176_),
        .dout(new_Jinkela_wire_2321)
    );

    bfr new_Jinkela_buffer_1408 (
        .din(new_Jinkela_wire_2255),
        .dout(new_Jinkela_wire_2256)
    );

    bfr new_Jinkela_buffer_818 (
        .din(_0155_),
        .dout(new_Jinkela_wire_1403)
    );

    and_bi _1076_ (
        .a(new_Jinkela_wire_2564),
        .b(new_Jinkela_wire_1037),
        .c(_0248_)
    );

    bfr new_Jinkela_buffer_793 (
        .din(new_Jinkela_wire_1375),
        .dout(new_Jinkela_wire_1376)
    );

    bfr new_Jinkela_buffer_1777 (
        .din(_0104_),
        .dout(new_Jinkela_wire_2824)
    );

    and_bi _1077_ (
        .a(new_Jinkela_wire_1156),
        .b(_0248_),
        .c(_0249_)
    );

    bfr new_Jinkela_buffer_817 (
        .din(new_Jinkela_wire_1401),
        .dout(new_Jinkela_wire_1402)
    );

    spl2 new_Jinkela_splitter_342 (
        .a(_0314_),
        .b(new_Jinkela_wire_2323),
        .c(new_Jinkela_wire_2324)
    );

    bfr new_Jinkela_buffer_1409 (
        .din(new_Jinkela_wire_2256),
        .dout(new_Jinkela_wire_2257)
    );

    bfr new_Jinkela_buffer_1775 (
        .din(new_Jinkela_wire_2821),
        .dout(new_Jinkela_wire_2822)
    );

    and_bi _1078_ (
        .a(new_Jinkela_wire_1406),
        .b(new_Jinkela_wire_935),
        .c(_0250_)
    );

    bfr new_Jinkela_buffer_794 (
        .din(new_Jinkela_wire_1376),
        .dout(new_Jinkela_wire_1377)
    );

    bfr new_Jinkela_buffer_1778 (
        .din(_0750_),
        .dout(new_Jinkela_wire_2825)
    );

    bfr new_Jinkela_buffer_7 (
        .din(new_Jinkela_wire_10),
        .dout(new_Jinkela_wire_11)
    );

    bfr new_Jinkela_buffer_31 (
        .din(new_Jinkela_wire_46),
        .dout(new_Jinkela_wire_47)
    );

    bfr new_Jinkela_buffer_8 (
        .din(new_Jinkela_wire_11),
        .dout(new_Jinkela_wire_12)
    );

    bfr new_Jinkela_buffer_28 (
        .din(new_Jinkela_wire_41),
        .dout(new_Jinkela_wire_42)
    );

    bfr new_Jinkela_buffer_9 (
        .din(new_Jinkela_wire_12),
        .dout(new_Jinkela_wire_13)
    );

    bfr new_Jinkela_buffer_10 (
        .din(new_Jinkela_wire_13),
        .dout(new_Jinkela_wire_14)
    );

    spl2 new_Jinkela_splitter_5 (
        .a(new_Jinkela_wire_42),
        .b(new_Jinkela_wire_43),
        .c(new_Jinkela_wire_44)
    );

    bfr new_Jinkela_buffer_11 (
        .din(new_Jinkela_wire_14),
        .dout(new_Jinkela_wire_15)
    );

    bfr new_Jinkela_buffer_77 (
        .din(new_Jinkela_wire_96),
        .dout(new_Jinkela_wire_97)
    );

    bfr new_Jinkela_buffer_12 (
        .din(new_Jinkela_wire_15),
        .dout(new_Jinkela_wire_16)
    );

    bfr new_Jinkela_buffer_32 (
        .din(new_Jinkela_wire_47),
        .dout(new_Jinkela_wire_48)
    );

    bfr new_Jinkela_buffer_13 (
        .din(new_Jinkela_wire_16),
        .dout(new_Jinkela_wire_17)
    );

    bfr new_Jinkela_buffer_33 (
        .din(new_Jinkela_wire_48),
        .dout(new_Jinkela_wire_49)
    );

    bfr new_Jinkela_buffer_14 (
        .din(new_Jinkela_wire_17),
        .dout(new_Jinkela_wire_18)
    );

    and_ii _0846_ (
        .a(_0019_),
        .b(_0018_),
        .c(_0020_)
    );

    bfr new_Jinkela_buffer_128 (
        .din(G31),
        .dout(new_Jinkela_wire_167)
    );

    bfr new_Jinkela_buffer_15 (
        .din(new_Jinkela_wire_18),
        .dout(new_Jinkela_wire_19)
    );

    bfr new_Jinkela_buffer_78 (
        .din(new_Jinkela_wire_97),
        .dout(new_Jinkela_wire_98)
    );

    bfr new_Jinkela_buffer_34 (
        .din(new_Jinkela_wire_49),
        .dout(new_Jinkela_wire_50)
    );

    bfr new_Jinkela_buffer_16 (
        .din(new_Jinkela_wire_19),
        .dout(new_Jinkela_wire_20)
    );

    bfr new_Jinkela_buffer_17 (
        .din(new_Jinkela_wire_20),
        .dout(new_Jinkela_wire_21)
    );

    spl3L new_Jinkela_splitter_10 (
        .a(new_Jinkela_wire_146),
        .d(new_Jinkela_wire_147),
        .b(new_Jinkela_wire_148),
        .c(new_Jinkela_wire_149)
    );

    bfr new_Jinkela_buffer_35 (
        .din(new_Jinkela_wire_50),
        .dout(new_Jinkela_wire_51)
    );

    bfr new_Jinkela_buffer_18 (
        .din(new_Jinkela_wire_21),
        .dout(new_Jinkela_wire_22)
    );

    spl4L new_Jinkela_splitter_11 (
        .a(new_Jinkela_wire_150),
        .d(new_Jinkela_wire_151),
        .e(new_Jinkela_wire_152),
        .b(new_Jinkela_wire_153),
        .c(new_Jinkela_wire_155)
    );

    bfr new_Jinkela_buffer_19 (
        .din(new_Jinkela_wire_22),
        .dout(new_Jinkela_wire_23)
    );

    bfr new_Jinkela_buffer_79 (
        .din(new_Jinkela_wire_98),
        .dout(new_Jinkela_wire_99)
    );

    bfr new_Jinkela_buffer_36 (
        .din(new_Jinkela_wire_51),
        .dout(new_Jinkela_wire_52)
    );

    spl4L new_Jinkela_splitter_2 (
        .a(new_Jinkela_wire_23),
        .d(new_Jinkela_wire_24),
        .e(new_Jinkela_wire_25),
        .b(new_Jinkela_wire_26),
        .c(new_Jinkela_wire_27)
    );

    bfr new_Jinkela_buffer_20 (
        .din(new_Jinkela_wire_27),
        .dout(new_Jinkela_wire_28)
    );

    bfr new_Jinkela_buffer_37 (
        .din(new_Jinkela_wire_52),
        .dout(new_Jinkela_wire_53)
    );

    bfr new_Jinkela_buffer_21 (
        .din(new_Jinkela_wire_28),
        .dout(new_Jinkela_wire_29)
    );

    bfr new_Jinkela_buffer_22 (
        .din(new_Jinkela_wire_29),
        .dout(new_Jinkela_wire_30)
    );

    bfr new_Jinkela_buffer_80 (
        .din(new_Jinkela_wire_99),
        .dout(new_Jinkela_wire_100)
    );

    bfr new_Jinkela_buffer_38 (
        .din(new_Jinkela_wire_53),
        .dout(new_Jinkela_wire_54)
    );

    bfr new_Jinkela_buffer_23 (
        .din(new_Jinkela_wire_30),
        .dout(new_Jinkela_wire_31)
    );

    bfr new_Jinkela_buffer_24 (
        .din(new_Jinkela_wire_31),
        .dout(new_Jinkela_wire_32)
    );

    spl2 new_Jinkela_splitter_23 (
        .a(G13),
        .b(new_Jinkela_wire_209),
        .c(new_Jinkela_wire_211)
    );

    bfr new_Jinkela_buffer_39 (
        .din(new_Jinkela_wire_54),
        .dout(new_Jinkela_wire_55)
    );

    bfr new_Jinkela_buffer_25 (
        .din(new_Jinkela_wire_32),
        .dout(new_Jinkela_wire_33)
    );

    spl4L new_Jinkela_splitter_14 (
        .a(new_Jinkela_wire_167),
        .d(new_Jinkela_wire_168),
        .e(new_Jinkela_wire_169),
        .b(new_Jinkela_wire_170),
        .c(new_Jinkela_wire_171)
    );

    bfr new_Jinkela_buffer_81 (
        .din(new_Jinkela_wire_100),
        .dout(new_Jinkela_wire_101)
    );

    bfr new_Jinkela_buffer_40 (
        .din(new_Jinkela_wire_55),
        .dout(new_Jinkela_wire_56)
    );

    spl2 new_Jinkela_splitter_213 (
        .a(_0100_),
        .b(new_Jinkela_wire_1290),
        .c(new_Jinkela_wire_1291)
    );

    bfr new_Jinkela_buffer_987 (
        .din(new_Jinkela_wire_1639),
        .dout(new_Jinkela_wire_1640)
    );

    bfr new_Jinkela_buffer_722 (
        .din(new_Jinkela_wire_1257),
        .dout(new_Jinkela_wire_1258)
    );

    bfr new_Jinkela_buffer_957 (
        .din(new_Jinkela_wire_1601),
        .dout(new_Jinkela_wire_1602)
    );

    bfr new_Jinkela_buffer_993 (
        .din(new_Jinkela_wire_1651),
        .dout(new_Jinkela_wire_1652)
    );

    bfr new_Jinkela_buffer_723 (
        .din(new_Jinkela_wire_1258),
        .dout(new_Jinkela_wire_1259)
    );

    bfr new_Jinkela_buffer_958 (
        .din(new_Jinkela_wire_1602),
        .dout(new_Jinkela_wire_1603)
    );

    bfr new_Jinkela_buffer_732 (
        .din(new_Jinkela_wire_1285),
        .dout(new_Jinkela_wire_1286)
    );

    bfr new_Jinkela_buffer_736 (
        .din(_0672_),
        .dout(new_Jinkela_wire_1294)
    );

    bfr new_Jinkela_buffer_1007 (
        .din(_0573_),
        .dout(new_Jinkela_wire_1679)
    );

    bfr new_Jinkela_buffer_724 (
        .din(new_Jinkela_wire_1259),
        .dout(new_Jinkela_wire_1260)
    );

    bfr new_Jinkela_buffer_959 (
        .din(new_Jinkela_wire_1603),
        .dout(new_Jinkela_wire_1604)
    );

    bfr new_Jinkela_buffer_742 (
        .din(_0462_),
        .dout(new_Jinkela_wire_1302)
    );

    bfr new_Jinkela_buffer_733 (
        .din(new_Jinkela_wire_1286),
        .dout(new_Jinkela_wire_1287)
    );

    bfr new_Jinkela_buffer_994 (
        .din(new_Jinkela_wire_1652),
        .dout(new_Jinkela_wire_1653)
    );

    bfr new_Jinkela_buffer_725 (
        .din(new_Jinkela_wire_1260),
        .dout(new_Jinkela_wire_1261)
    );

    bfr new_Jinkela_buffer_960 (
        .din(new_Jinkela_wire_1604),
        .dout(new_Jinkela_wire_1605)
    );

    spl2 new_Jinkela_splitter_214 (
        .a(new_Jinkela_wire_1291),
        .b(new_Jinkela_wire_1292),
        .c(new_Jinkela_wire_1293)
    );

    bfr new_Jinkela_buffer_726 (
        .din(new_Jinkela_wire_1261),
        .dout(new_Jinkela_wire_1262)
    );

    bfr new_Jinkela_buffer_961 (
        .din(new_Jinkela_wire_1605),
        .dout(new_Jinkela_wire_1606)
    );

    bfr new_Jinkela_buffer_734 (
        .din(new_Jinkela_wire_1287),
        .dout(new_Jinkela_wire_1288)
    );

    bfr new_Jinkela_buffer_995 (
        .din(new_Jinkela_wire_1653),
        .dout(new_Jinkela_wire_1654)
    );

    bfr new_Jinkela_buffer_962 (
        .din(new_Jinkela_wire_1606),
        .dout(new_Jinkela_wire_1607)
    );

    bfr new_Jinkela_buffer_738 (
        .din(new_Jinkela_wire_1295),
        .dout(new_Jinkela_wire_1296)
    );

    bfr new_Jinkela_buffer_1009 (
        .din(_0604_),
        .dout(new_Jinkela_wire_1681)
    );

    bfr new_Jinkela_buffer_963 (
        .din(new_Jinkela_wire_1607),
        .dout(new_Jinkela_wire_1608)
    );

    bfr new_Jinkela_buffer_749 (
        .din(_0538_),
        .dout(new_Jinkela_wire_1309)
    );

    bfr new_Jinkela_buffer_737 (
        .din(new_Jinkela_wire_1294),
        .dout(new_Jinkela_wire_1295)
    );

    bfr new_Jinkela_buffer_743 (
        .din(new_Jinkela_wire_1302),
        .dout(new_Jinkela_wire_1303)
    );

    bfr new_Jinkela_buffer_964 (
        .din(new_Jinkela_wire_1608),
        .dout(new_Jinkela_wire_1609)
    );

    spl2 new_Jinkela_splitter_261 (
        .a(new_Jinkela_wire_1670),
        .b(new_Jinkela_wire_1671),
        .c(new_Jinkela_wire_1672)
    );

    bfr new_Jinkela_buffer_996 (
        .din(new_Jinkela_wire_1654),
        .dout(new_Jinkela_wire_1655)
    );

    bfr new_Jinkela_buffer_764 (
        .din(_0330_),
        .dout(new_Jinkela_wire_1324)
    );

    bfr new_Jinkela_buffer_965 (
        .din(new_Jinkela_wire_1609),
        .dout(new_Jinkela_wire_1610)
    );

    bfr new_Jinkela_buffer_739 (
        .din(new_Jinkela_wire_1296),
        .dout(new_Jinkela_wire_1297)
    );

    bfr new_Jinkela_buffer_1004 (
        .din(new_Jinkela_wire_1669),
        .dout(new_Jinkela_wire_1670)
    );

    bfr new_Jinkela_buffer_997 (
        .din(new_Jinkela_wire_1655),
        .dout(new_Jinkela_wire_1656)
    );

    bfr new_Jinkela_buffer_744 (
        .din(new_Jinkela_wire_1303),
        .dout(new_Jinkela_wire_1304)
    );

    bfr new_Jinkela_buffer_966 (
        .din(new_Jinkela_wire_1610),
        .dout(new_Jinkela_wire_1611)
    );

    bfr new_Jinkela_buffer_740 (
        .din(new_Jinkela_wire_1297),
        .dout(new_Jinkela_wire_1298)
    );

    bfr new_Jinkela_buffer_750 (
        .din(new_Jinkela_wire_1309),
        .dout(new_Jinkela_wire_1310)
    );

    bfr new_Jinkela_buffer_967 (
        .din(new_Jinkela_wire_1611),
        .dout(new_Jinkela_wire_1612)
    );

    bfr new_Jinkela_buffer_741 (
        .din(new_Jinkela_wire_1298),
        .dout(new_Jinkela_wire_1299)
    );

    spl2 new_Jinkela_splitter_263 (
        .a(new_Jinkela_wire_1676),
        .b(new_Jinkela_wire_1677),
        .c(new_Jinkela_wire_1678)
    );

    bfr new_Jinkela_buffer_998 (
        .din(new_Jinkela_wire_1656),
        .dout(new_Jinkela_wire_1657)
    );

    bfr new_Jinkela_buffer_745 (
        .din(new_Jinkela_wire_1304),
        .dout(new_Jinkela_wire_1305)
    );

    bfr new_Jinkela_buffer_968 (
        .din(new_Jinkela_wire_1612),
        .dout(new_Jinkela_wire_1613)
    );

    spl2 new_Jinkela_splitter_215 (
        .a(new_Jinkela_wire_1299),
        .b(new_Jinkela_wire_1300),
        .c(new_Jinkela_wire_1301)
    );

    bfr new_Jinkela_buffer_746 (
        .din(new_Jinkela_wire_1305),
        .dout(new_Jinkela_wire_1306)
    );

    bfr new_Jinkela_buffer_969 (
        .din(new_Jinkela_wire_1613),
        .dout(new_Jinkela_wire_1614)
    );

    bfr new_Jinkela_buffer_769 (
        .din(_0073_),
        .dout(new_Jinkela_wire_1329)
    );

    bfr new_Jinkela_buffer_1006 (
        .din(_0459_),
        .dout(new_Jinkela_wire_1676)
    );

    bfr new_Jinkela_buffer_999 (
        .din(new_Jinkela_wire_1657),
        .dout(new_Jinkela_wire_1658)
    );

    bfr new_Jinkela_buffer_751 (
        .din(new_Jinkela_wire_1310),
        .dout(new_Jinkela_wire_1311)
    );

    bfr new_Jinkela_buffer_970 (
        .din(new_Jinkela_wire_1614),
        .dout(new_Jinkela_wire_1615)
    );

    bfr new_Jinkela_buffer_747 (
        .din(new_Jinkela_wire_1306),
        .dout(new_Jinkela_wire_1307)
    );

    bfr new_Jinkela_buffer_765 (
        .din(new_Jinkela_wire_1324),
        .dout(new_Jinkela_wire_1325)
    );

    bfr new_Jinkela_buffer_971 (
        .din(new_Jinkela_wire_1615),
        .dout(new_Jinkela_wire_1616)
    );

    bfr new_Jinkela_buffer_748 (
        .din(new_Jinkela_wire_1307),
        .dout(new_Jinkela_wire_1308)
    );

    bfr new_Jinkela_buffer_1000 (
        .din(new_Jinkela_wire_1658),
        .dout(new_Jinkela_wire_1659)
    );

    bfr new_Jinkela_buffer_752 (
        .din(new_Jinkela_wire_1311),
        .dout(new_Jinkela_wire_1312)
    );

    bfr new_Jinkela_buffer_972 (
        .din(new_Jinkela_wire_1616),
        .dout(new_Jinkela_wire_1617)
    );

    spl2 new_Jinkela_splitter_216 (
        .a(_0023_),
        .b(new_Jinkela_wire_1330),
        .c(new_Jinkela_wire_1331)
    );

    bfr new_Jinkela_buffer_770 (
        .din(_0187_),
        .dout(new_Jinkela_wire_1332)
    );

    bfr new_Jinkela_buffer_753 (
        .din(new_Jinkela_wire_1312),
        .dout(new_Jinkela_wire_1313)
    );

    bfr new_Jinkela_buffer_973 (
        .din(new_Jinkela_wire_1617),
        .dout(new_Jinkela_wire_1618)
    );

    bfr new_Jinkela_buffer_766 (
        .din(new_Jinkela_wire_1325),
        .dout(new_Jinkela_wire_1326)
    );

    spl2 new_Jinkela_splitter_264 (
        .a(_0794_),
        .b(new_Jinkela_wire_1684),
        .c(new_Jinkela_wire_1685)
    );

    bfr new_Jinkela_buffer_1001 (
        .din(new_Jinkela_wire_1659),
        .dout(new_Jinkela_wire_1660)
    );

    bfr new_Jinkela_buffer_754 (
        .din(new_Jinkela_wire_1313),
        .dout(new_Jinkela_wire_1314)
    );

    bfr new_Jinkela_buffer_974 (
        .din(new_Jinkela_wire_1618),
        .dout(new_Jinkela_wire_1619)
    );

    bfr new_Jinkela_buffer_772 (
        .din(_0407_),
        .dout(new_Jinkela_wire_1334)
    );

    bfr new_Jinkela_buffer_778 (
        .din(_0731_),
        .dout(new_Jinkela_wire_1350)
    );

    bfr new_Jinkela_buffer_755 (
        .din(new_Jinkela_wire_1314),
        .dout(new_Jinkela_wire_1315)
    );

    bfr new_Jinkela_buffer_1008 (
        .din(new_Jinkela_wire_1679),
        .dout(new_Jinkela_wire_1680)
    );

    bfr new_Jinkela_buffer_1002 (
        .din(new_Jinkela_wire_1660),
        .dout(new_Jinkela_wire_1661)
    );

    bfr new_Jinkela_buffer_767 (
        .din(new_Jinkela_wire_1326),
        .dout(new_Jinkela_wire_1327)
    );

    bfr new_Jinkela_buffer_1018 (
        .din(_0590_),
        .dout(new_Jinkela_wire_1698)
    );

    bfr new_Jinkela_buffer_756 (
        .din(new_Jinkela_wire_1315),
        .dout(new_Jinkela_wire_1316)
    );

    bfr new_Jinkela_buffer_1010 (
        .din(new_Jinkela_wire_1681),
        .dout(new_Jinkela_wire_1682)
    );

    bfr new_Jinkela_buffer_1003 (
        .din(new_Jinkela_wire_1661),
        .dout(new_Jinkela_wire_1662)
    );

    bfr new_Jinkela_buffer_757 (
        .din(new_Jinkela_wire_1316),
        .dout(new_Jinkela_wire_1317)
    );

    spl4L new_Jinkela_splitter_259 (
        .a(new_Jinkela_wire_1662),
        .d(new_Jinkela_wire_1663),
        .e(new_Jinkela_wire_1664),
        .b(new_Jinkela_wire_1665),
        .c(new_Jinkela_wire_1666)
    );

    bfr new_Jinkela_buffer_768 (
        .din(new_Jinkela_wire_1327),
        .dout(new_Jinkela_wire_1328)
    );

    spl2 new_Jinkela_splitter_343 (
        .a(_0361_),
        .b(new_Jinkela_wire_2332),
        .c(new_Jinkela_wire_2333)
    );

    bfr new_Jinkela_buffer_1750 (
        .din(new_Jinkela_wire_2793),
        .dout(new_Jinkela_wire_2794)
    );

    or_bb _1415_ (
        .a(new_Jinkela_wire_1983),
        .b(_0578_),
        .c(_0581_)
    );

    bfr new_Jinkela_buffer_1445 (
        .din(new_Jinkela_wire_2324),
        .dout(new_Jinkela_wire_2325)
    );

    bfr new_Jinkela_buffer_1410 (
        .din(new_Jinkela_wire_2257),
        .dout(new_Jinkela_wire_2258)
    );

    bfr new_Jinkela_buffer_1780 (
        .din(_0291_),
        .dout(new_Jinkela_wire_2829)
    );

    or_bb _1416_ (
        .a(_0581_),
        .b(new_Jinkela_wire_2583),
        .c(_0582_)
    );

    bfr new_Jinkela_buffer_1776 (
        .din(new_Jinkela_wire_2822),
        .dout(new_Jinkela_wire_2823)
    );

    bfr new_Jinkela_buffer_1751 (
        .din(new_Jinkela_wire_2794),
        .dout(new_Jinkela_wire_2795)
    );

    and_bi _1417_ (
        .a(new_Jinkela_wire_1950),
        .b(new_Jinkela_wire_3000),
        .c(_0583_)
    );

    bfr new_Jinkela_buffer_1411 (
        .din(new_Jinkela_wire_2258),
        .dout(new_Jinkela_wire_2259)
    );

    and_bi _1418_ (
        .a(new_Jinkela_wire_403),
        .b(new_Jinkela_wire_1887),
        .c(_0584_)
    );

    bfr new_Jinkela_buffer_1779 (
        .din(new_Jinkela_wire_2825),
        .dout(new_Jinkela_wire_2826)
    );

    spl2 new_Jinkela_splitter_344 (
        .a(_0154_),
        .b(new_Jinkela_wire_2334),
        .c(new_Jinkela_wire_2335)
    );

    bfr new_Jinkela_buffer_1752 (
        .din(new_Jinkela_wire_2795),
        .dout(new_Jinkela_wire_2796)
    );

    or_bb _1419_ (
        .a(_0584_),
        .b(new_Jinkela_wire_1241),
        .c(_0585_)
    );

    bfr new_Jinkela_buffer_1453 (
        .din(new_Jinkela_wire_2336),
        .dout(new_Jinkela_wire_2337)
    );

    bfr new_Jinkela_buffer_1412 (
        .din(new_Jinkela_wire_2259),
        .dout(new_Jinkela_wire_2260)
    );

    or_bb _1420_ (
        .a(new_Jinkela_wire_1368),
        .b(new_Jinkela_wire_842),
        .c(_0586_)
    );

    bfr new_Jinkela_buffer_1781 (
        .din(_0542_),
        .dout(new_Jinkela_wire_2830)
    );

    spl3L new_Jinkela_splitter_405 (
        .a(new_Jinkela_wire_2796),
        .d(new_Jinkela_wire_2797),
        .b(new_Jinkela_wire_2798),
        .c(new_Jinkela_wire_2799)
    );

    or_bb _1421_ (
        .a(_0586_),
        .b(_0583_),
        .c(_0587_)
    );

    bfr new_Jinkela_buffer_1413 (
        .din(new_Jinkela_wire_2260),
        .dout(new_Jinkela_wire_2261)
    );

    or_bb _1422_ (
        .a(_0587_),
        .b(new_Jinkela_wire_2406),
        .c(_0588_)
    );

    bfr new_Jinkela_buffer_1446 (
        .din(new_Jinkela_wire_2325),
        .dout(new_Jinkela_wire_2326)
    );

    bfr new_Jinkela_buffer_1753 (
        .din(new_Jinkela_wire_2799),
        .dout(new_Jinkela_wire_2800)
    );

    or_bi _1423_ (
        .a(new_Jinkela_wire_1874),
        .b(new_Jinkela_wire_320),
        .c(_0589_)
    );

    bfr new_Jinkela_buffer_1414 (
        .din(new_Jinkela_wire_2261),
        .dout(new_Jinkela_wire_2262)
    );

    bfr new_Jinkela_buffer_1783 (
        .din(_0297_),
        .dout(new_Jinkela_wire_2834)
    );

    or_bb _1424_ (
        .a(new_Jinkela_wire_689),
        .b(new_Jinkela_wire_713),
        .c(_0590_)
    );

    bfr new_Jinkela_buffer_1782 (
        .din(new_Jinkela_wire_2830),
        .dout(new_Jinkela_wire_2831)
    );

    bfr new_Jinkela_buffer_1452 (
        .din(_0275_),
        .dout(new_Jinkela_wire_2336)
    );

    bfr new_Jinkela_buffer_1754 (
        .din(new_Jinkela_wire_2800),
        .dout(new_Jinkela_wire_2801)
    );

    and_bi _1425_ (
        .a(new_Jinkela_wire_1705),
        .b(new_Jinkela_wire_1138),
        .c(_0591_)
    );

    spl2 new_Jinkela_splitter_346 (
        .a(_0368_),
        .b(new_Jinkela_wire_2346),
        .c(new_Jinkela_wire_2349)
    );

    bfr new_Jinkela_buffer_1415 (
        .din(new_Jinkela_wire_2262),
        .dout(new_Jinkela_wire_2263)
    );

    spl2 new_Jinkela_splitter_406 (
        .a(new_Jinkela_wire_2826),
        .b(new_Jinkela_wire_2827),
        .c(new_Jinkela_wire_2828)
    );

    and_bi _1426_ (
        .a(new_Jinkela_wire_3018),
        .b(_0591_),
        .c(_0592_)
    );

    bfr new_Jinkela_buffer_1447 (
        .din(new_Jinkela_wire_2326),
        .dout(new_Jinkela_wire_2327)
    );

    bfr new_Jinkela_buffer_1755 (
        .din(new_Jinkela_wire_2801),
        .dout(new_Jinkela_wire_2802)
    );

    and_bi _1427_ (
        .a(new_Jinkela_wire_688),
        .b(new_Jinkela_wire_2363),
        .c(_0593_)
    );

    bfr new_Jinkela_buffer_1416 (
        .din(new_Jinkela_wire_2263),
        .dout(new_Jinkela_wire_2264)
    );

    and_bi _1428_ (
        .a(new_Jinkela_wire_2394),
        .b(new_Jinkela_wire_1743),
        .c(_0594_)
    );

    bfr new_Jinkela_buffer_1756 (
        .din(new_Jinkela_wire_2802),
        .dout(new_Jinkela_wire_2803)
    );

    or_bb _1429_ (
        .a(new_Jinkela_wire_2582),
        .b(_0593_),
        .c(_0595_)
    );

    bfr new_Jinkela_buffer_1455 (
        .din(_0284_),
        .dout(new_Jinkela_wire_2339)
    );

    bfr new_Jinkela_buffer_1448 (
        .din(new_Jinkela_wire_2327),
        .dout(new_Jinkela_wire_2328)
    );

    and_bi _1430_ (
        .a(_0592_),
        .b(_0595_),
        .c(_0596_)
    );

    bfr new_Jinkela_buffer_1791 (
        .din(_0673_),
        .dout(new_Jinkela_wire_2842)
    );

    bfr new_Jinkela_buffer_1757 (
        .din(new_Jinkela_wire_2803),
        .dout(new_Jinkela_wire_2804)
    );

    and_bi _1431_ (
        .a(new_Jinkela_wire_251),
        .b(new_Jinkela_wire_3001),
        .c(_0597_)
    );

    bfr new_Jinkela_buffer_1449 (
        .din(new_Jinkela_wire_2328),
        .dout(new_Jinkela_wire_2329)
    );

    and_ii _1432_ (
        .a(new_Jinkela_wire_2270),
        .b(new_Jinkela_wire_2412),
        .c(_0598_)
    );

    bfr new_Jinkela_buffer_1784 (
        .din(new_Jinkela_wire_2834),
        .dout(new_Jinkela_wire_2835)
    );

    bfr new_Jinkela_buffer_1758 (
        .din(new_Jinkela_wire_2804),
        .dout(new_Jinkela_wire_2805)
    );

    or_bb _1433_ (
        .a(_0598_),
        .b(new_Jinkela_wire_3088),
        .c(_0599_)
    );

    bfr new_Jinkela_buffer_1454 (
        .din(new_Jinkela_wire_2337),
        .dout(new_Jinkela_wire_2338)
    );

    bfr new_Jinkela_buffer_1450 (
        .din(new_Jinkela_wire_2329),
        .dout(new_Jinkela_wire_2330)
    );

    spl2 new_Jinkela_splitter_407 (
        .a(new_Jinkela_wire_2831),
        .b(new_Jinkela_wire_2832),
        .c(new_Jinkela_wire_2833)
    );

    or_bb _1434_ (
        .a(new_Jinkela_wire_1650),
        .b(_0597_),
        .c(_0600_)
    );

    bfr new_Jinkela_buffer_1759 (
        .din(new_Jinkela_wire_2805),
        .dout(new_Jinkela_wire_2806)
    );

    and_bi _1435_ (
        .a(new_Jinkela_wire_3189),
        .b(_0600_),
        .c(_0601_)
    );

    bfr new_Jinkela_buffer_1451 (
        .din(new_Jinkela_wire_2330),
        .dout(new_Jinkela_wire_2331)
    );

    and_bi _1436_ (
        .a(_0588_),
        .b(_0601_),
        .c(_0602_)
    );

    bfr new_Jinkela_buffer_1785 (
        .din(new_Jinkela_wire_2835),
        .dout(new_Jinkela_wire_2836)
    );

    bfr new_Jinkela_buffer_1456 (
        .din(new_Jinkela_wire_2339),
        .dout(new_Jinkela_wire_2340)
    );

    bfr new_Jinkela_buffer_1760 (
        .din(new_Jinkela_wire_2806),
        .dout(new_Jinkela_wire_2807)
    );

    and_bi _1437_ (
        .a(new_Jinkela_wire_1908),
        .b(_0602_),
        .c(_0603_)
    );

    bfr new_Jinkela_buffer_1463 (
        .din(_0481_),
        .dout(new_Jinkela_wire_2373)
    );

    or_bb _1438_ (
        .a(_0603_),
        .b(new_Jinkela_wire_1341),
        .c(_0604_)
    );

    spl4L new_Jinkela_splitter_347 (
        .a(new_Jinkela_wire_2349),
        .d(new_Jinkela_wire_2350),
        .e(new_Jinkela_wire_2355),
        .b(new_Jinkela_wire_2360),
        .c(new_Jinkela_wire_2365)
    );

    bfr new_Jinkela_buffer_1792 (
        .din(_0780_),
        .dout(new_Jinkela_wire_2843)
    );

    bfr new_Jinkela_buffer_1457 (
        .din(new_Jinkela_wire_2340),
        .dout(new_Jinkela_wire_2341)
    );

    bfr new_Jinkela_buffer_1761 (
        .din(new_Jinkela_wire_2807),
        .dout(new_Jinkela_wire_2808)
    );

    and_bi _1439_ (
        .a(_0576_),
        .b(new_Jinkela_wire_1683),
        .c(_0605_)
    );

    and_bi _1440_ (
        .a(new_Jinkela_wire_1552),
        .b(new_Jinkela_wire_1485),
        .c(_0606_)
    );

    bfr new_Jinkela_buffer_1460 (
        .din(new_Jinkela_wire_2346),
        .dout(new_Jinkela_wire_2347)
    );

    bfr new_Jinkela_buffer_1818 (
        .din(_0335_),
        .dout(new_Jinkela_wire_2869)
    );

    spl2 new_Jinkela_splitter_345 (
        .a(new_Jinkela_wire_2341),
        .b(new_Jinkela_wire_2342),
        .c(new_Jinkela_wire_2343)
    );

    bfr new_Jinkela_buffer_1762 (
        .din(new_Jinkela_wire_2808),
        .dout(new_Jinkela_wire_2809)
    );

    and_ii _1441_ (
        .a(_0606_),
        .b(new_Jinkela_wire_2537),
        .c(_0607_)
    );

    bfr new_Jinkela_buffer_1458 (
        .din(new_Jinkela_wire_2343),
        .dout(new_Jinkela_wire_2344)
    );

    and_bi _1442_ (
        .a(new_Jinkela_wire_1736),
        .b(new_Jinkela_wire_1182),
        .c(_0608_)
    );

    bfr new_Jinkela_buffer_1786 (
        .din(new_Jinkela_wire_2836),
        .dout(new_Jinkela_wire_2837)
    );

    bfr new_Jinkela_buffer_1462 (
        .din(new_Jinkela_wire_2371),
        .dout(new_Jinkela_wire_2372)
    );

    bfr new_Jinkela_buffer_1763 (
        .din(new_Jinkela_wire_2809),
        .dout(new_Jinkela_wire_2810)
    );

    or_bb _1443_ (
        .a(_0608_),
        .b(new_Jinkela_wire_820),
        .c(_0609_)
    );

    spl2 new_Jinkela_splitter_352 (
        .a(_0087_),
        .b(new_Jinkela_wire_2370),
        .c(new_Jinkela_wire_2371)
    );

    or_bb _1444_ (
        .a(_0609_),
        .b(new_Jinkela_wire_1356),
        .c(new_net_6)
    );

    bfr new_Jinkela_buffer_1793 (
        .din(new_Jinkela_wire_2843),
        .dout(new_Jinkela_wire_2844)
    );

    bfr new_Jinkela_buffer_1459 (
        .din(new_Jinkela_wire_2344),
        .dout(new_Jinkela_wire_2345)
    );

    bfr new_Jinkela_buffer_1764 (
        .din(new_Jinkela_wire_2810),
        .dout(new_Jinkela_wire_2811)
    );

    and_bb _1445_ (
        .a(new_Jinkela_wire_831),
        .b(new_Jinkela_wire_2890),
        .c(_0610_)
    );

    or_bi _1446_ (
        .a(_0610_),
        .b(new_Jinkela_wire_1550),
        .c(_0611_)
    );

    spl2 new_Jinkela_splitter_354 (
        .a(_0189_),
        .b(new_Jinkela_wire_2381),
        .c(new_Jinkela_wire_2382)
    );

    bfr new_Jinkela_buffer_1787 (
        .din(new_Jinkela_wire_2837),
        .dout(new_Jinkela_wire_2838)
    );

    bfr new_Jinkela_buffer_1467 (
        .din(_0408_),
        .dout(new_Jinkela_wire_2379)
    );

    bfr new_Jinkela_buffer_1765 (
        .din(new_Jinkela_wire_2811),
        .dout(new_Jinkela_wire_2812)
    );

    and_bi _1447_ (
        .a(new_Jinkela_wire_2898),
        .b(new_Jinkela_wire_1735),
        .c(_0612_)
    );

    bfr new_Jinkela_buffer_1461 (
        .din(new_Jinkela_wire_2347),
        .dout(new_Jinkela_wire_2348)
    );

    and_ii _1448_ (
        .a(_0612_),
        .b(new_Jinkela_wire_2070),
        .c(_0613_)
    );

    spl4L new_Jinkela_splitter_349 (
        .a(new_Jinkela_wire_2355),
        .d(new_Jinkela_wire_2356),
        .e(new_Jinkela_wire_2357),
        .b(new_Jinkela_wire_2358),
        .c(new_Jinkela_wire_2359)
    );

    bfr new_Jinkela_buffer_1823 (
        .din(_0141_),
        .dout(new_Jinkela_wire_2874)
    );

    bfr new_Jinkela_buffer_1766 (
        .din(new_Jinkela_wire_2812),
        .dout(new_Jinkela_wire_2813)
    );

    or_bb _1449_ (
        .a(_0613_),
        .b(new_Jinkela_wire_2542),
        .c(_0614_)
    );

    spl4L new_Jinkela_splitter_348 (
        .a(new_Jinkela_wire_2350),
        .d(new_Jinkela_wire_2351),
        .e(new_Jinkela_wire_2352),
        .b(new_Jinkela_wire_2353),
        .c(new_Jinkela_wire_2354)
    );

    and_bi _1450_ (
        .a(new_Jinkela_wire_1199),
        .b(new_Jinkela_wire_2198),
        .c(_0615_)
    );

    bfr new_Jinkela_buffer_1788 (
        .din(new_Jinkela_wire_2838),
        .dout(new_Jinkela_wire_2839)
    );

    bfr new_Jinkela_buffer_1469 (
        .din(_0381_),
        .dout(new_Jinkela_wire_2383)
    );

    bfr new_Jinkela_buffer_1767 (
        .din(new_Jinkela_wire_2813),
        .dout(new_Jinkela_wire_2814)
    );

    or_bb _1451_ (
        .a(new_Jinkela_wire_1000),
        .b(new_Jinkela_wire_2003),
        .c(_0616_)
    );

    spl4L new_Jinkela_splitter_350 (
        .a(new_Jinkela_wire_2360),
        .d(new_Jinkela_wire_2361),
        .e(new_Jinkela_wire_2362),
        .b(new_Jinkela_wire_2363),
        .c(new_Jinkela_wire_2364)
    );

    and_bi _1452_ (
        .a(new_Jinkela_wire_1169),
        .b(new_Jinkela_wire_2968),
        .c(_0617_)
    );

    spl4L new_Jinkela_splitter_351 (
        .a(new_Jinkela_wire_2365),
        .d(new_Jinkela_wire_2366),
        .e(new_Jinkela_wire_2367),
        .b(new_Jinkela_wire_2368),
        .c(new_Jinkela_wire_2369)
    );

    bfr new_Jinkela_buffer_1794 (
        .din(new_Jinkela_wire_2844),
        .dout(new_Jinkela_wire_2845)
    );

    bfr new_Jinkela_buffer_1768 (
        .din(new_Jinkela_wire_2814),
        .dout(new_Jinkela_wire_2815)
    );

    inv _1453_ (
        .din(_0617_),
        .dout(_0618_)
    );

    and_bi _1454_ (
        .a(new_Jinkela_wire_2435),
        .b(new_Jinkela_wire_2303),
        .c(_0619_)
    );

    spl2 new_Jinkela_splitter_353 (
        .a(new_Jinkela_wire_2373),
        .b(new_Jinkela_wire_2374),
        .c(new_Jinkela_wire_2375)
    );

    bfr new_Jinkela_buffer_1789 (
        .din(new_Jinkela_wire_2839),
        .dout(new_Jinkela_wire_2840)
    );

    bfr new_Jinkela_buffer_1464 (
        .din(new_Jinkela_wire_2375),
        .dout(new_Jinkela_wire_2376)
    );

    bfr new_Jinkela_buffer_1769 (
        .din(new_Jinkela_wire_2815),
        .dout(new_Jinkela_wire_2816)
    );

    and_bi _1455_ (
        .a(new_Jinkela_wire_2304),
        .b(new_Jinkela_wire_2434),
        .c(_0621_)
    );

    bfr new_Jinkela_buffer_1468 (
        .din(new_Jinkela_wire_2379),
        .dout(new_Jinkela_wire_2380)
    );

    and_ii _1456_ (
        .a(_0621_),
        .b(_0619_),
        .c(_0622_)
    );

    bfr new_Jinkela_buffer_1819 (
        .din(new_Jinkela_wire_2869),
        .dout(new_Jinkela_wire_2870)
    );

    bfr new_Jinkela_buffer_1770 (
        .din(new_Jinkela_wire_2816),
        .dout(new_Jinkela_wire_2817)
    );

    bfr new_Jinkela_buffer_1011 (
        .din(new_Jinkela_wire_1682),
        .dout(new_Jinkela_wire_1683)
    );

    spl2 new_Jinkela_splitter_268 (
        .a(_0036_),
        .b(new_Jinkela_wire_1707),
        .c(new_Jinkela_wire_1708)
    );

    bfr new_Jinkela_buffer_1790 (
        .din(new_Jinkela_wire_2840),
        .dout(new_Jinkela_wire_2841)
    );

    bfr new_Jinkela_buffer_1771 (
        .din(new_Jinkela_wire_2817),
        .dout(new_Jinkela_wire_2818)
    );

    bfr new_Jinkela_buffer_1026 (
        .din(_0666_),
        .dout(new_Jinkela_wire_1706)
    );

    bfr new_Jinkela_buffer_1019 (
        .din(new_Jinkela_wire_1698),
        .dout(new_Jinkela_wire_1699)
    );

    bfr new_Jinkela_buffer_1012 (
        .din(new_Jinkela_wire_1685),
        .dout(new_Jinkela_wire_1686)
    );

    bfr new_Jinkela_buffer_1795 (
        .din(new_Jinkela_wire_2845),
        .dout(new_Jinkela_wire_2846)
    );

    bfr new_Jinkela_buffer_1772 (
        .din(new_Jinkela_wire_2818),
        .dout(new_Jinkela_wire_2819)
    );

    bfr new_Jinkela_buffer_1027 (
        .din(_0172_),
        .dout(new_Jinkela_wire_1709)
    );

    bfr new_Jinkela_buffer_1824 (
        .din(_0329_),
        .dout(new_Jinkela_wire_2875)
    );

    bfr new_Jinkela_buffer_1773 (
        .din(new_Jinkela_wire_2819),
        .dout(new_Jinkela_wire_2820)
    );

    spl2 new_Jinkela_splitter_266 (
        .a(new_Jinkela_wire_1688),
        .b(new_Jinkela_wire_1689),
        .c(new_Jinkela_wire_1690)
    );

    bfr new_Jinkela_buffer_1020 (
        .din(new_Jinkela_wire_1699),
        .dout(new_Jinkela_wire_1700)
    );

    spl2 new_Jinkela_splitter_265 (
        .a(new_Jinkela_wire_1686),
        .b(new_Jinkela_wire_1687),
        .c(new_Jinkela_wire_1688)
    );

    bfr new_Jinkela_buffer_1796 (
        .din(new_Jinkela_wire_2846),
        .dout(new_Jinkela_wire_2847)
    );

    bfr new_Jinkela_buffer_1013 (
        .din(new_Jinkela_wire_1690),
        .dout(new_Jinkela_wire_1691)
    );

    bfr new_Jinkela_buffer_1820 (
        .din(new_Jinkela_wire_2870),
        .dout(new_Jinkela_wire_2871)
    );

    bfr new_Jinkela_buffer_1797 (
        .din(new_Jinkela_wire_2847),
        .dout(new_Jinkela_wire_2848)
    );

    bfr new_Jinkela_buffer_1035 (
        .din(new_Jinkela_wire_1726),
        .dout(new_Jinkela_wire_1727)
    );

    bfr new_Jinkela_buffer_1021 (
        .din(new_Jinkela_wire_1700),
        .dout(new_Jinkela_wire_1701)
    );

    spl2 new_Jinkela_splitter_408 (
        .a(_0115_),
        .b(new_Jinkela_wire_2876),
        .c(new_Jinkela_wire_2877)
    );

    spl3L new_Jinkela_splitter_409 (
        .a(_0139_),
        .d(new_Jinkela_wire_2878),
        .b(new_Jinkela_wire_2879),
        .c(new_Jinkela_wire_2880)
    );

    bfr new_Jinkela_buffer_1014 (
        .din(new_Jinkela_wire_1691),
        .dout(new_Jinkela_wire_1692)
    );

    bfr new_Jinkela_buffer_1798 (
        .din(new_Jinkela_wire_2848),
        .dout(new_Jinkela_wire_2849)
    );

    bfr new_Jinkela_buffer_1821 (
        .din(new_Jinkela_wire_2871),
        .dout(new_Jinkela_wire_2872)
    );

    spl2 new_Jinkela_splitter_272 (
        .a(_0302_),
        .b(new_Jinkela_wire_1724),
        .c(new_Jinkela_wire_1725)
    );

    spl2 new_Jinkela_splitter_267 (
        .a(new_Jinkela_wire_1692),
        .b(new_Jinkela_wire_1693),
        .c(new_Jinkela_wire_1694)
    );

    bfr new_Jinkela_buffer_1799 (
        .din(new_Jinkela_wire_2849),
        .dout(new_Jinkela_wire_2850)
    );

    bfr new_Jinkela_buffer_1015 (
        .din(new_Jinkela_wire_1694),
        .dout(new_Jinkela_wire_1695)
    );

    spl3L new_Jinkela_splitter_413 (
        .a(new_net_2),
        .d(new_Jinkela_wire_2899),
        .b(new_Jinkela_wire_2900),
        .c(new_Jinkela_wire_2901)
    );

    bfr new_Jinkela_buffer_1826 (
        .din(new_Jinkela_wire_2883),
        .dout(new_Jinkela_wire_2884)
    );

    bfr new_Jinkela_buffer_1022 (
        .din(new_Jinkela_wire_1701),
        .dout(new_Jinkela_wire_1702)
    );

    bfr new_Jinkela_buffer_1800 (
        .din(new_Jinkela_wire_2850),
        .dout(new_Jinkela_wire_2851)
    );

    bfr new_Jinkela_buffer_1034 (
        .din(_0120_),
        .dout(new_Jinkela_wire_1726)
    );

    bfr new_Jinkela_buffer_1822 (
        .din(new_Jinkela_wire_2872),
        .dout(new_Jinkela_wire_2873)
    );

    bfr new_Jinkela_buffer_1016 (
        .din(new_Jinkela_wire_1695),
        .dout(new_Jinkela_wire_1696)
    );

    bfr new_Jinkela_buffer_1801 (
        .din(new_Jinkela_wire_2851),
        .dout(new_Jinkela_wire_2852)
    );

    bfr new_Jinkela_buffer_1023 (
        .din(new_Jinkela_wire_1702),
        .dout(new_Jinkela_wire_1703)
    );

    bfr new_Jinkela_buffer_1017 (
        .din(new_Jinkela_wire_1696),
        .dout(new_Jinkela_wire_1697)
    );

    bfr new_Jinkela_buffer_1802 (
        .din(new_Jinkela_wire_2852),
        .dout(new_Jinkela_wire_2853)
    );

    spl2 new_Jinkela_splitter_410 (
        .a(_0135_),
        .b(new_Jinkela_wire_2881),
        .c(new_Jinkela_wire_2882)
    );

    bfr new_Jinkela_buffer_1036 (
        .din(_0058_),
        .dout(new_Jinkela_wire_1728)
    );

    bfr new_Jinkela_buffer_1024 (
        .din(new_Jinkela_wire_1703),
        .dout(new_Jinkela_wire_1704)
    );

    bfr new_Jinkela_buffer_1803 (
        .din(new_Jinkela_wire_2853),
        .dout(new_Jinkela_wire_2854)
    );

    spl4L new_Jinkela_splitter_411 (
        .a(_0338_),
        .d(new_Jinkela_wire_2886),
        .e(new_Jinkela_wire_2887),
        .b(new_Jinkela_wire_2888),
        .c(new_Jinkela_wire_2889)
    );

    bfr new_Jinkela_buffer_1025 (
        .din(new_Jinkela_wire_1704),
        .dout(new_Jinkela_wire_1705)
    );

    bfr new_Jinkela_buffer_1804 (
        .din(new_Jinkela_wire_2854),
        .dout(new_Jinkela_wire_2855)
    );

    bfr new_Jinkela_buffer_1028 (
        .din(new_Jinkela_wire_1709),
        .dout(new_Jinkela_wire_1710)
    );

    bfr new_Jinkela_buffer_1825 (
        .din(_0702_),
        .dout(new_Jinkela_wire_2883)
    );

    bfr new_Jinkela_buffer_1029 (
        .din(new_Jinkela_wire_1710),
        .dout(new_Jinkela_wire_1711)
    );

    bfr new_Jinkela_buffer_1805 (
        .din(new_Jinkela_wire_2855),
        .dout(new_Jinkela_wire_2856)
    );

    bfr new_Jinkela_buffer_1037 (
        .din(_0654_),
        .dout(new_Jinkela_wire_1729)
    );

    spl4L new_Jinkela_splitter_269 (
        .a(new_Jinkela_wire_1711),
        .d(new_Jinkela_wire_1712),
        .e(new_Jinkela_wire_1713),
        .b(new_Jinkela_wire_1714),
        .c(new_Jinkela_wire_1715)
    );

    spl4L new_Jinkela_splitter_412 (
        .a(new_Jinkela_wire_2889),
        .d(new_Jinkela_wire_2890),
        .e(new_Jinkela_wire_2891),
        .b(new_Jinkela_wire_2892),
        .c(new_Jinkela_wire_2893)
    );

    bfr new_Jinkela_buffer_1844 (
        .din(_0090_),
        .dout(new_Jinkela_wire_2913)
    );

    bfr new_Jinkela_buffer_1806 (
        .din(new_Jinkela_wire_2856),
        .dout(new_Jinkela_wire_2857)
    );

    bfr new_Jinkela_buffer_1030 (
        .din(new_Jinkela_wire_1715),
        .dout(new_Jinkela_wire_1716)
    );

    bfr new_Jinkela_buffer_1827 (
        .din(new_Jinkela_wire_2884),
        .dout(new_Jinkela_wire_2885)
    );

    spl3L new_Jinkela_splitter_273 (
        .a(_0564_),
        .d(new_Jinkela_wire_1734),
        .b(new_Jinkela_wire_1735),
        .c(new_Jinkela_wire_1736)
    );

    bfr new_Jinkela_buffer_1807 (
        .din(new_Jinkela_wire_2857),
        .dout(new_Jinkela_wire_2858)
    );

    spl3L new_Jinkela_splitter_274 (
        .a(_0377_),
        .d(new_Jinkela_wire_1737),
        .b(new_Jinkela_wire_1742),
        .c(new_Jinkela_wire_1747)
    );

    bfr new_Jinkela_buffer_1038 (
        .din(new_Jinkela_wire_1729),
        .dout(new_Jinkela_wire_1730)
    );

    bfr new_Jinkela_buffer_1833 (
        .din(new_Jinkela_wire_2901),
        .dout(new_Jinkela_wire_2902)
    );

    spl2 new_Jinkela_splitter_270 (
        .a(new_Jinkela_wire_1716),
        .b(new_Jinkela_wire_1717),
        .c(new_Jinkela_wire_1718)
    );

    bfr new_Jinkela_buffer_1808 (
        .din(new_Jinkela_wire_2858),
        .dout(new_Jinkela_wire_2859)
    );

    spl2 new_Jinkela_splitter_271 (
        .a(new_Jinkela_wire_1718),
        .b(new_Jinkela_wire_1719),
        .c(new_Jinkela_wire_1720)
    );

    bfr new_Jinkela_buffer_1809 (
        .din(new_Jinkela_wire_2859),
        .dout(new_Jinkela_wire_2860)
    );

    bfr new_Jinkela_buffer_1031 (
        .din(new_Jinkela_wire_1720),
        .dout(new_Jinkela_wire_1721)
    );

    bfr new_Jinkela_buffer_1039 (
        .din(new_Jinkela_wire_1730),
        .dout(new_Jinkela_wire_1731)
    );

    bfr new_Jinkela_buffer_1810 (
        .din(new_Jinkela_wire_2860),
        .dout(new_Jinkela_wire_2861)
    );

    bfr new_Jinkela_buffer_1048 (
        .din(_0427_),
        .dout(new_Jinkela_wire_1761)
    );

    bfr new_Jinkela_buffer_1828 (
        .din(new_Jinkela_wire_2893),
        .dout(new_Jinkela_wire_2894)
    );

    bfr new_Jinkela_buffer_1032 (
        .din(new_Jinkela_wire_1721),
        .dout(new_Jinkela_wire_1722)
    );

    bfr new_Jinkela_buffer_1811 (
        .din(new_Jinkela_wire_2861),
        .dout(new_Jinkela_wire_2862)
    );

    bfr new_Jinkela_buffer_1040 (
        .din(new_Jinkela_wire_1731),
        .dout(new_Jinkela_wire_1732)
    );

    bfr new_Jinkela_buffer_1846 (
        .din(new_net_1479),
        .dout(new_Jinkela_wire_2915)
    );

    bfr new_Jinkela_buffer_1033 (
        .din(new_Jinkela_wire_1722),
        .dout(new_Jinkela_wire_1723)
    );

    bfr new_Jinkela_buffer_1812 (
        .din(new_Jinkela_wire_2862),
        .dout(new_Jinkela_wire_2863)
    );

    spl3L new_Jinkela_splitter_278 (
        .a(_0271_),
        .d(new_Jinkela_wire_1752),
        .b(new_Jinkela_wire_1753),
        .c(new_Jinkela_wire_1754)
    );

    bfr new_Jinkela_buffer_1829 (
        .din(new_Jinkela_wire_2894),
        .dout(new_Jinkela_wire_2895)
    );

    bfr new_Jinkela_buffer_1041 (
        .din(new_Jinkela_wire_1732),
        .dout(new_Jinkela_wire_1733)
    );

    bfr new_Jinkela_buffer_1813 (
        .din(new_Jinkela_wire_2863),
        .dout(new_Jinkela_wire_2864)
    );

    bfr new_Jinkela_buffer_688 (
        .din(new_Jinkela_wire_1217),
        .dout(new_Jinkela_wire_1218)
    );

    bfr new_Jinkela_buffer_706 (
        .din(_0378_),
        .dout(new_Jinkela_wire_1240)
    );

    bfr new_Jinkela_buffer_708 (
        .din(_0409_),
        .dout(new_Jinkela_wire_1244)
    );

    bfr new_Jinkela_buffer_689 (
        .din(new_Jinkela_wire_1218),
        .dout(new_Jinkela_wire_1219)
    );

    bfr new_Jinkela_buffer_705 (
        .din(new_Jinkela_wire_1238),
        .dout(new_Jinkela_wire_1239)
    );

    bfr new_Jinkela_buffer_690 (
        .din(new_Jinkela_wire_1219),
        .dout(new_Jinkela_wire_1220)
    );

    spl2 new_Jinkela_splitter_205 (
        .a(_0126_),
        .b(new_Jinkela_wire_1263),
        .c(new_Jinkela_wire_1264)
    );

    bfr new_Jinkela_buffer_691 (
        .din(new_Jinkela_wire_1220),
        .dout(new_Jinkela_wire_1221)
    );

    spl2 new_Jinkela_splitter_204 (
        .a(new_Jinkela_wire_1240),
        .b(new_Jinkela_wire_1241),
        .c(new_Jinkela_wire_1242)
    );

    bfr new_Jinkela_buffer_692 (
        .din(new_Jinkela_wire_1221),
        .dout(new_Jinkela_wire_1222)
    );

    bfr new_Jinkela_buffer_707 (
        .din(new_Jinkela_wire_1242),
        .dout(new_Jinkela_wire_1243)
    );

    bfr new_Jinkela_buffer_693 (
        .din(new_Jinkela_wire_1222),
        .dout(new_Jinkela_wire_1223)
    );

    bfr new_Jinkela_buffer_727 (
        .din(_0448_),
        .dout(new_Jinkela_wire_1267)
    );

    bfr new_Jinkela_buffer_694 (
        .din(new_Jinkela_wire_1223),
        .dout(new_Jinkela_wire_1224)
    );

    bfr new_Jinkela_buffer_709 (
        .din(new_Jinkela_wire_1244),
        .dout(new_Jinkela_wire_1245)
    );

    bfr new_Jinkela_buffer_695 (
        .din(new_Jinkela_wire_1224),
        .dout(new_Jinkela_wire_1225)
    );

    spl2 new_Jinkela_splitter_206 (
        .a(new_Jinkela_wire_1264),
        .b(new_Jinkela_wire_1265),
        .c(new_Jinkela_wire_1266)
    );

    bfr new_Jinkela_buffer_696 (
        .din(new_Jinkela_wire_1225),
        .dout(new_Jinkela_wire_1226)
    );

    bfr new_Jinkela_buffer_710 (
        .din(new_Jinkela_wire_1245),
        .dout(new_Jinkela_wire_1246)
    );

    bfr new_Jinkela_buffer_697 (
        .din(new_Jinkela_wire_1226),
        .dout(new_Jinkela_wire_1227)
    );

    spl2 new_Jinkela_splitter_207 (
        .a(_0020_),
        .b(new_Jinkela_wire_1269),
        .c(new_Jinkela_wire_1270)
    );

    bfr new_Jinkela_buffer_711 (
        .din(new_Jinkela_wire_1246),
        .dout(new_Jinkela_wire_1247)
    );

    spl2 new_Jinkela_splitter_208 (
        .a(_0784_),
        .b(new_Jinkela_wire_1271),
        .c(new_Jinkela_wire_1272)
    );

    bfr new_Jinkela_buffer_712 (
        .din(new_Jinkela_wire_1247),
        .dout(new_Jinkela_wire_1248)
    );

    spl2 new_Jinkela_splitter_209 (
        .a(_0663_),
        .b(new_Jinkela_wire_1276),
        .c(new_Jinkela_wire_1277)
    );

    bfr new_Jinkela_buffer_713 (
        .din(new_Jinkela_wire_1248),
        .dout(new_Jinkela_wire_1249)
    );

    bfr new_Jinkela_buffer_728 (
        .din(new_Jinkela_wire_1267),
        .dout(new_Jinkela_wire_1268)
    );

    bfr new_Jinkela_buffer_714 (
        .din(new_Jinkela_wire_1249),
        .dout(new_Jinkela_wire_1250)
    );

    bfr new_Jinkela_buffer_715 (
        .din(new_Jinkela_wire_1250),
        .dout(new_Jinkela_wire_1251)
    );

    bfr new_Jinkela_buffer_729 (
        .din(_0215_),
        .dout(new_Jinkela_wire_1273)
    );

    bfr new_Jinkela_buffer_716 (
        .din(new_Jinkela_wire_1251),
        .dout(new_Jinkela_wire_1252)
    );

    bfr new_Jinkela_buffer_730 (
        .din(_0668_),
        .dout(new_Jinkela_wire_1274)
    );

    spl2 new_Jinkela_splitter_210 (
        .a(_0199_),
        .b(new_Jinkela_wire_1278),
        .c(new_Jinkela_wire_1279)
    );

    bfr new_Jinkela_buffer_717 (
        .din(new_Jinkela_wire_1252),
        .dout(new_Jinkela_wire_1253)
    );

    bfr new_Jinkela_buffer_731 (
        .din(new_Jinkela_wire_1274),
        .dout(new_Jinkela_wire_1275)
    );

    bfr new_Jinkela_buffer_718 (
        .din(new_Jinkela_wire_1253),
        .dout(new_Jinkela_wire_1254)
    );

    bfr new_Jinkela_buffer_719 (
        .din(new_Jinkela_wire_1254),
        .dout(new_Jinkela_wire_1255)
    );

    spl4L new_Jinkela_splitter_211 (
        .a(_0057_),
        .d(new_Jinkela_wire_1280),
        .e(new_Jinkela_wire_1281),
        .b(new_Jinkela_wire_1282),
        .c(new_Jinkela_wire_1283)
    );

    bfr new_Jinkela_buffer_720 (
        .din(new_Jinkela_wire_1255),
        .dout(new_Jinkela_wire_1256)
    );

    spl2 new_Jinkela_splitter_212 (
        .a(_0069_),
        .b(new_Jinkela_wire_1284),
        .c(new_Jinkela_wire_1285)
    );

    bfr new_Jinkela_buffer_721 (
        .din(new_Jinkela_wire_1256),
        .dout(new_Jinkela_wire_1257)
    );

    bfr new_Jinkela_buffer_735 (
        .din(_0108_),
        .dout(new_Jinkela_wire_1289)
    );

    or_ii _1079_ (
        .a(new_Jinkela_wire_2655),
        .b(new_Jinkela_wire_2387),
        .c(_0251_)
    );

    spl2 new_Jinkela_splitter_17 (
        .a(G19),
        .b(new_Jinkela_wire_178),
        .c(new_Jinkela_wire_179)
    );

    bfr new_Jinkela_buffer_41 (
        .din(new_Jinkela_wire_56),
        .dout(new_Jinkela_wire_57)
    );

    inv _1080_ (
        .din(new_Jinkela_wire_276),
        .dout(_0252_)
    );

    and_bi _1081_ (
        .a(new_Jinkela_wire_2444),
        .b(new_Jinkela_wire_3194),
        .c(_0253_)
    );

    spl2 new_Jinkela_splitter_8 (
        .a(new_Jinkela_wire_101),
        .b(new_Jinkela_wire_102),
        .c(new_Jinkela_wire_103)
    );

    bfr new_Jinkela_buffer_42 (
        .din(new_Jinkela_wire_57),
        .dout(new_Jinkela_wire_58)
    );

    or_bb _1082_ (
        .a(_0253_),
        .b(new_Jinkela_wire_2401),
        .c(_0254_)
    );

    and_bi _1083_ (
        .a(new_Jinkela_wire_3300),
        .b(new_Jinkela_wire_289),
        .c(_0255_)
    );

    bfr new_Jinkela_buffer_82 (
        .din(new_Jinkela_wire_103),
        .dout(new_Jinkela_wire_104)
    );

    bfr new_Jinkela_buffer_43 (
        .din(new_Jinkela_wire_58),
        .dout(new_Jinkela_wire_59)
    );

    and_bb _1084_ (
        .a(new_Jinkela_wire_238),
        .b(new_Jinkela_wire_435),
        .c(_0256_)
    );

    and_bi _1085_ (
        .a(new_Jinkela_wire_2334),
        .b(new_Jinkela_wire_2407),
        .c(_0257_)
    );

    bfr new_Jinkela_buffer_44 (
        .din(new_Jinkela_wire_59),
        .dout(new_Jinkela_wire_60)
    );

    and_bi _1086_ (
        .a(new_Jinkela_wire_1033),
        .b(_0257_),
        .c(_0258_)
    );

    spl4L new_Jinkela_splitter_13 (
        .a(new_Jinkela_wire_159),
        .d(new_Jinkela_wire_160),
        .e(new_Jinkela_wire_161),
        .b(new_Jinkela_wire_162),
        .c(new_Jinkela_wire_163)
    );

    or_bb _1087_ (
        .a(_0258_),
        .b(_0255_),
        .c(_0259_)
    );

    bfr new_Jinkela_buffer_124 (
        .din(new_Jinkela_wire_153),
        .dout(new_Jinkela_wire_154)
    );

    bfr new_Jinkela_buffer_45 (
        .din(new_Jinkela_wire_60),
        .dout(new_Jinkela_wire_61)
    );

    and_bi _1088_ (
        .a(_0254_),
        .b(new_Jinkela_wire_2789),
        .c(_0260_)
    );

    or_ii _1089_ (
        .a(new_Jinkela_wire_2177),
        .b(new_Jinkela_wire_785),
        .c(_0261_)
    );

    bfr new_Jinkela_buffer_83 (
        .din(new_Jinkela_wire_104),
        .dout(new_Jinkela_wire_105)
    );

    bfr new_Jinkela_buffer_46 (
        .din(new_Jinkela_wire_61),
        .dout(new_Jinkela_wire_62)
    );

    and_bb _1090_ (
        .a(new_Jinkela_wire_430),
        .b(new_Jinkela_wire_515),
        .c(_0262_)
    );

    and_bi _1091_ (
        .a(new_Jinkela_wire_525),
        .b(new_Jinkela_wire_429),
        .c(_0263_)
    );

    spl4L new_Jinkela_splitter_12 (
        .a(new_Jinkela_wire_155),
        .d(new_Jinkela_wire_156),
        .e(new_Jinkela_wire_157),
        .b(new_Jinkela_wire_158),
        .c(new_Jinkela_wire_159)
    );

    bfr new_Jinkela_buffer_47 (
        .din(new_Jinkela_wire_62),
        .dout(new_Jinkela_wire_63)
    );

    or_bb _1092_ (
        .a(_0263_),
        .b(_0262_),
        .c(_0264_)
    );

    spl2 new_Jinkela_splitter_20 (
        .a(G9),
        .b(new_Jinkela_wire_191),
        .c(new_Jinkela_wire_193)
    );

    and_bi _1093_ (
        .a(new_Jinkela_wire_485),
        .b(new_Jinkela_wire_3033),
        .c(_0265_)
    );

    bfr new_Jinkela_buffer_84 (
        .din(new_Jinkela_wire_105),
        .dout(new_Jinkela_wire_106)
    );

    bfr new_Jinkela_buffer_48 (
        .din(new_Jinkela_wire_63),
        .dout(new_Jinkela_wire_64)
    );

    or_bb _1094_ (
        .a(_0265_),
        .b(new_Jinkela_wire_2431),
        .c(_0266_)
    );

    and_bi _1095_ (
        .a(new_Jinkela_wire_2575),
        .b(_0266_),
        .c(_0267_)
    );

    bfr new_Jinkela_buffer_49 (
        .din(new_Jinkela_wire_64),
        .dout(new_Jinkela_wire_65)
    );

    and_bi _1096_ (
        .a(new_Jinkela_wire_1044),
        .b(_0267_),
        .c(_0268_)
    );

    bfr new_Jinkela_buffer_129 (
        .din(new_Jinkela_wire_171),
        .dout(new_Jinkela_wire_172)
    );

    or_bb _1097_ (
        .a(new_Jinkela_wire_1355),
        .b(new_Jinkela_wire_964),
        .c(_0269_)
    );

    bfr new_Jinkela_buffer_85 (
        .din(new_Jinkela_wire_106),
        .dout(new_Jinkela_wire_107)
    );

    bfr new_Jinkela_buffer_50 (
        .din(new_Jinkela_wire_65),
        .dout(new_Jinkela_wire_66)
    );

    or_bb _1098_ (
        .a(new_Jinkela_wire_2274),
        .b(new_Jinkela_wire_3061),
        .c(_0270_)
    );

    or_bb _1099_ (
        .a(_0270_),
        .b(new_Jinkela_wire_1890),
        .c(_0271_)
    );

    bfr new_Jinkela_buffer_51 (
        .din(new_Jinkela_wire_66),
        .dout(new_Jinkela_wire_67)
    );

    or_bb _1100_ (
        .a(new_Jinkela_wire_1760),
        .b(new_Jinkela_wire_2938),
        .c(_0272_)
    );

    bfr new_Jinkela_buffer_125 (
        .din(new_Jinkela_wire_163),
        .dout(new_Jinkela_wire_164)
    );

    and_bi _1101_ (
        .a(new_Jinkela_wire_2386),
        .b(new_Jinkela_wire_1412),
        .c(_0273_)
    );

    bfr new_Jinkela_buffer_86 (
        .din(new_Jinkela_wire_107),
        .dout(new_Jinkela_wire_108)
    );

    bfr new_Jinkela_buffer_52 (
        .din(new_Jinkela_wire_67),
        .dout(new_Jinkela_wire_68)
    );

    and_bi _1102_ (
        .a(new_Jinkela_wire_1200),
        .b(new_Jinkela_wire_1278),
        .c(_0274_)
    );

    or_bb _1103_ (
        .a(_0274_),
        .b(new_Jinkela_wire_1501),
        .c(_0275_)
    );

    bfr new_Jinkela_buffer_53 (
        .din(new_Jinkela_wire_68),
        .dout(new_Jinkela_wire_69)
    );

    or_bb _1104_ (
        .a(new_Jinkela_wire_2338),
        .b(_0273_),
        .c(_0276_)
    );

    spl2 new_Jinkela_splitter_15 (
        .a(new_Jinkela_wire_172),
        .b(new_Jinkela_wire_173),
        .c(new_Jinkela_wire_174)
    );

    and_bi _1105_ (
        .a(_0272_),
        .b(new_Jinkela_wire_1627),
        .c(_0277_)
    );

    bfr new_Jinkela_buffer_87 (
        .din(new_Jinkela_wire_108),
        .dout(new_Jinkela_wire_109)
    );

    bfr new_Jinkela_buffer_54 (
        .din(new_Jinkela_wire_69),
        .dout(new_Jinkela_wire_70)
    );

    and_ii _1106_ (
        .a(new_Jinkela_wire_1646),
        .b(new_Jinkela_wire_2072),
        .c(_0278_)
    );

    and_bi _1107_ (
        .a(new_Jinkela_wire_2879),
        .b(new_Jinkela_wire_835),
        .c(_0279_)
    );

    spl4L new_Jinkela_splitter_21 (
        .a(new_Jinkela_wire_193),
        .d(new_Jinkela_wire_194),
        .e(new_Jinkela_wire_195),
        .b(new_Jinkela_wire_196),
        .c(new_Jinkela_wire_197)
    );

    bfr new_Jinkela_buffer_55 (
        .din(new_Jinkela_wire_70),
        .dout(new_Jinkela_wire_71)
    );

    and_ii _1108_ (
        .a(_0279_),
        .b(new_Jinkela_wire_3017),
        .c(_0280_)
    );

    and_bi _1109_ (
        .a(new_Jinkela_wire_2876),
        .b(new_Jinkela_wire_2385),
        .c(_0281_)
    );

    bfr new_Jinkela_buffer_88 (
        .din(new_Jinkela_wire_109),
        .dout(new_Jinkela_wire_110)
    );

    bfr new_Jinkela_buffer_56 (
        .din(new_Jinkela_wire_71),
        .dout(new_Jinkela_wire_72)
    );

    and_bb _1110_ (
        .a(new_Jinkela_wire_2284),
        .b(new_Jinkela_wire_1228),
        .c(_0282_)
    );

    or_bb _1111_ (
        .a(_0282_),
        .b(new_Jinkela_wire_2372),
        .c(_0283_)
    );

    spl2 new_Jinkela_splitter_18 (
        .a(new_Jinkela_wire_179),
        .b(new_Jinkela_wire_180),
        .c(new_Jinkela_wire_181)
    );

    bfr new_Jinkela_buffer_57 (
        .din(new_Jinkela_wire_72),
        .dout(new_Jinkela_wire_73)
    );

    or_bb _1112_ (
        .a(new_Jinkela_wire_1232),
        .b(_0281_),
        .c(_0284_)
    );

    bfr new_Jinkela_buffer_126 (
        .din(new_Jinkela_wire_164),
        .dout(new_Jinkela_wire_165)
    );

    or_bb _1113_ (
        .a(new_Jinkela_wire_2342),
        .b(_0278_),
        .c(new_net_1465)
    );

    bfr new_Jinkela_buffer_89 (
        .din(new_Jinkela_wire_110),
        .dout(new_Jinkela_wire_111)
    );

    bfr new_Jinkela_buffer_58 (
        .din(new_Jinkela_wire_73),
        .dout(new_Jinkela_wire_74)
    );

    or_ii _1114_ (
        .a(new_Jinkela_wire_95),
        .b(new_Jinkela_wire_343),
        .c(_0285_)
    );

    and_bi _1115_ (
        .a(new_Jinkela_wire_3231),
        .b(new_Jinkela_wire_2220),
        .c(_0286_)
    );

    bfr new_Jinkela_buffer_59 (
        .din(new_Jinkela_wire_74),
        .dout(new_Jinkela_wire_75)
    );

    inv _1116_ (
        .din(new_Jinkela_wire_2190),
        .dout(_0287_)
    );

    or_bb _1117_ (
        .a(new_Jinkela_wire_1354),
        .b(new_Jinkela_wire_2010),
        .c(_0288_)
    );

    bfr new_Jinkela_buffer_90 (
        .din(new_Jinkela_wire_111),
        .dout(new_Jinkela_wire_112)
    );

    bfr new_Jinkela_buffer_60 (
        .din(new_Jinkela_wire_75),
        .dout(new_Jinkela_wire_76)
    );

    or_bb _1118_ (
        .a(new_Jinkela_wire_1206),
        .b(new_Jinkela_wire_658),
        .c(_0289_)
    );

    or_bb _1119_ (
        .a(_0289_),
        .b(_0288_),
        .c(_0290_)
    );

    bfr new_Jinkela_buffer_61 (
        .din(new_Jinkela_wire_76),
        .dout(new_Jinkela_wire_77)
    );

    or_bb _1120_ (
        .a(_0290_),
        .b(new_Jinkela_wire_2586),
        .c(_0291_)
    );

    bfr new_Jinkela_buffer_1834 (
        .din(new_Jinkela_wire_2902),
        .dout(new_Jinkela_wire_2903)
    );

    bfr new_Jinkela_buffer_662 (
        .din(_0398_),
        .dout(new_Jinkela_wire_1183)
    );

    bfr new_Jinkela_buffer_1845 (
        .din(new_Jinkela_wire_2913),
        .dout(new_Jinkela_wire_2914)
    );

    bfr new_Jinkela_buffer_655 (
        .din(new_Jinkela_wire_1173),
        .dout(new_Jinkela_wire_1174)
    );

    bfr new_Jinkela_buffer_1814 (
        .din(new_Jinkela_wire_2864),
        .dout(new_Jinkela_wire_2865)
    );

    bfr new_Jinkela_buffer_668 (
        .din(_0096_),
        .dout(new_Jinkela_wire_1191)
    );

    bfr new_Jinkela_buffer_1830 (
        .din(new_Jinkela_wire_2895),
        .dout(new_Jinkela_wire_2896)
    );

    bfr new_Jinkela_buffer_669 (
        .din(new_Jinkela_wire_1191),
        .dout(new_Jinkela_wire_1192)
    );

    bfr new_Jinkela_buffer_656 (
        .din(new_Jinkela_wire_1174),
        .dout(new_Jinkela_wire_1175)
    );

    bfr new_Jinkela_buffer_1815 (
        .din(new_Jinkela_wire_2865),
        .dout(new_Jinkela_wire_2866)
    );

    bfr new_Jinkela_buffer_670 (
        .din(_0529_),
        .dout(new_Jinkela_wire_1193)
    );

    spl2 new_Jinkela_splitter_198 (
        .a(new_Jinkela_wire_1175),
        .b(new_Jinkela_wire_1176),
        .c(new_Jinkela_wire_1177)
    );

    bfr new_Jinkela_buffer_1816 (
        .din(new_Jinkela_wire_2866),
        .dout(new_Jinkela_wire_2867)
    );

    bfr new_Jinkela_buffer_657 (
        .din(new_Jinkela_wire_1177),
        .dout(new_Jinkela_wire_1178)
    );

    bfr new_Jinkela_buffer_1831 (
        .din(new_Jinkela_wire_2896),
        .dout(new_Jinkela_wire_2897)
    );

    bfr new_Jinkela_buffer_663 (
        .din(new_Jinkela_wire_1183),
        .dout(new_Jinkela_wire_1184)
    );

    bfr new_Jinkela_buffer_1817 (
        .din(new_Jinkela_wire_2867),
        .dout(new_Jinkela_wire_2868)
    );

    bfr new_Jinkela_buffer_664 (
        .din(new_Jinkela_wire_1184),
        .dout(new_Jinkela_wire_1185)
    );

    bfr new_Jinkela_buffer_1851 (
        .din(_0365_),
        .dout(new_Jinkela_wire_2920)
    );

    bfr new_Jinkela_buffer_1835 (
        .din(new_Jinkela_wire_2903),
        .dout(new_Jinkela_wire_2904)
    );

    bfr new_Jinkela_buffer_1832 (
        .din(new_Jinkela_wire_2897),
        .dout(new_Jinkela_wire_2898)
    );

    bfr new_Jinkela_buffer_672 (
        .din(_0694_),
        .dout(new_Jinkela_wire_1195)
    );

    bfr new_Jinkela_buffer_665 (
        .din(new_Jinkela_wire_1185),
        .dout(new_Jinkela_wire_1186)
    );

    spl2 new_Jinkela_splitter_415 (
        .a(_0414_),
        .b(new_Jinkela_wire_2927),
        .c(new_Jinkela_wire_2928)
    );

    bfr new_Jinkela_buffer_1847 (
        .din(new_Jinkela_wire_2915),
        .dout(new_Jinkela_wire_2916)
    );

    bfr new_Jinkela_buffer_1836 (
        .din(new_Jinkela_wire_2904),
        .dout(new_Jinkela_wire_2905)
    );

    bfr new_Jinkela_buffer_671 (
        .din(new_Jinkela_wire_1193),
        .dout(new_Jinkela_wire_1194)
    );

    bfr new_Jinkela_buffer_666 (
        .din(new_Jinkela_wire_1186),
        .dout(new_Jinkela_wire_1187)
    );

    bfr new_Jinkela_buffer_1837 (
        .din(new_Jinkela_wire_2905),
        .dout(new_Jinkela_wire_2906)
    );

    spl3L new_Jinkela_splitter_200 (
        .a(_0225_),
        .d(new_Jinkela_wire_1198),
        .b(new_Jinkela_wire_1199),
        .c(new_Jinkela_wire_1200)
    );

    spl2 new_Jinkela_splitter_417 (
        .a(_0251_),
        .b(new_Jinkela_wire_2937),
        .c(new_Jinkela_wire_2938)
    );

    spl2 new_Jinkela_splitter_199 (
        .a(new_Jinkela_wire_1187),
        .b(new_Jinkela_wire_1188),
        .c(new_Jinkela_wire_1189)
    );

    bfr new_Jinkela_buffer_1848 (
        .din(new_Jinkela_wire_2916),
        .dout(new_Jinkela_wire_2917)
    );

    bfr new_Jinkela_buffer_1838 (
        .din(new_Jinkela_wire_2906),
        .dout(new_Jinkela_wire_2907)
    );

    bfr new_Jinkela_buffer_667 (
        .din(new_Jinkela_wire_1189),
        .dout(new_Jinkela_wire_1190)
    );

    bfr new_Jinkela_buffer_675 (
        .din(_0705_),
        .dout(new_Jinkela_wire_1201)
    );

    bfr new_Jinkela_buffer_673 (
        .din(new_Jinkela_wire_1195),
        .dout(new_Jinkela_wire_1196)
    );

    bfr new_Jinkela_buffer_1839 (
        .din(new_Jinkela_wire_2907),
        .dout(new_Jinkela_wire_2908)
    );

    bfr new_Jinkela_buffer_1852 (
        .din(new_Jinkela_wire_2920),
        .dout(new_Jinkela_wire_2921)
    );

    spl4L new_Jinkela_splitter_201 (
        .a(_0195_),
        .d(new_Jinkela_wire_1203),
        .e(new_Jinkela_wire_1204),
        .b(new_Jinkela_wire_1205),
        .c(new_Jinkela_wire_1206)
    );

    bfr new_Jinkela_buffer_1849 (
        .din(new_Jinkela_wire_2917),
        .dout(new_Jinkela_wire_2918)
    );

    bfr new_Jinkela_buffer_674 (
        .din(new_Jinkela_wire_1196),
        .dout(new_Jinkela_wire_1197)
    );

    bfr new_Jinkela_buffer_1840 (
        .din(new_Jinkela_wire_2908),
        .dout(new_Jinkela_wire_2909)
    );

    bfr new_Jinkela_buffer_677 (
        .din(_0709_),
        .dout(new_Jinkela_wire_1207)
    );

    bfr new_Jinkela_buffer_676 (
        .din(new_Jinkela_wire_1201),
        .dout(new_Jinkela_wire_1202)
    );

    bfr new_Jinkela_buffer_1841 (
        .din(new_Jinkela_wire_2909),
        .dout(new_Jinkela_wire_2910)
    );

    bfr new_Jinkela_buffer_1850 (
        .din(new_Jinkela_wire_2918),
        .dout(new_Jinkela_wire_2919)
    );

    spl2 new_Jinkela_splitter_202 (
        .a(_0084_),
        .b(new_Jinkela_wire_1228),
        .c(new_Jinkela_wire_1229)
    );

    bfr new_Jinkela_buffer_1842 (
        .din(new_Jinkela_wire_2910),
        .dout(new_Jinkela_wire_2911)
    );

    bfr new_Jinkela_buffer_678 (
        .din(new_Jinkela_wire_1207),
        .dout(new_Jinkela_wire_1208)
    );

    bfr new_Jinkela_buffer_679 (
        .din(_0757_),
        .dout(new_Jinkela_wire_1209)
    );

    bfr new_Jinkela_buffer_698 (
        .din(_0283_),
        .dout(new_Jinkela_wire_1230)
    );

    bfr new_Jinkela_buffer_1843 (
        .din(new_Jinkela_wire_2911),
        .dout(new_Jinkela_wire_2912)
    );

    bfr new_Jinkela_buffer_680 (
        .din(new_Jinkela_wire_1209),
        .dout(new_Jinkela_wire_1210)
    );

    bfr new_Jinkela_buffer_1853 (
        .din(new_Jinkela_wire_2921),
        .dout(new_Jinkela_wire_2922)
    );

    bfr new_Jinkela_buffer_702 (
        .din(_0534_),
        .dout(new_Jinkela_wire_1236)
    );

    bfr new_Jinkela_buffer_699 (
        .din(new_Jinkela_wire_1230),
        .dout(new_Jinkela_wire_1231)
    );

    bfr new_Jinkela_buffer_1856 (
        .din(new_Jinkela_wire_2928),
        .dout(new_Jinkela_wire_2929)
    );

    bfr new_Jinkela_buffer_681 (
        .din(new_Jinkela_wire_1210),
        .dout(new_Jinkela_wire_1211)
    );

    bfr new_Jinkela_buffer_1854 (
        .din(new_Jinkela_wire_2922),
        .dout(new_Jinkela_wire_2923)
    );

    spl2 new_Jinkela_splitter_418 (
        .a(_0796_),
        .b(new_Jinkela_wire_2939),
        .c(new_Jinkela_wire_2940)
    );

    bfr new_Jinkela_buffer_682 (
        .din(new_Jinkela_wire_1211),
        .dout(new_Jinkela_wire_1212)
    );

    spl2 new_Jinkela_splitter_414 (
        .a(new_Jinkela_wire_2923),
        .b(new_Jinkela_wire_2924),
        .c(new_Jinkela_wire_2925)
    );

    bfr new_Jinkela_buffer_701 (
        .din(_0762_),
        .dout(new_Jinkela_wire_1233)
    );

    bfr new_Jinkela_buffer_1855 (
        .din(new_Jinkela_wire_2925),
        .dout(new_Jinkela_wire_2926)
    );

    bfr new_Jinkela_buffer_683 (
        .din(new_Jinkela_wire_1212),
        .dout(new_Jinkela_wire_1213)
    );

    spl4L new_Jinkela_splitter_419 (
        .a(_0791_),
        .d(new_Jinkela_wire_2944),
        .e(new_Jinkela_wire_2945),
        .b(new_Jinkela_wire_2946),
        .c(new_Jinkela_wire_2947)
    );

    bfr new_Jinkela_buffer_1857 (
        .din(new_Jinkela_wire_2929),
        .dout(new_Jinkela_wire_2930)
    );

    bfr new_Jinkela_buffer_703 (
        .din(_0166_),
        .dout(new_Jinkela_wire_1237)
    );

    bfr new_Jinkela_buffer_1862 (
        .din(new_Jinkela_wire_2940),
        .dout(new_Jinkela_wire_2941)
    );

    bfr new_Jinkela_buffer_684 (
        .din(new_Jinkela_wire_1213),
        .dout(new_Jinkela_wire_1214)
    );

    bfr new_Jinkela_buffer_1858 (
        .din(new_Jinkela_wire_2930),
        .dout(new_Jinkela_wire_2931)
    );

    bfr new_Jinkela_buffer_700 (
        .din(new_Jinkela_wire_1231),
        .dout(new_Jinkela_wire_1232)
    );

    bfr new_Jinkela_buffer_685 (
        .din(new_Jinkela_wire_1214),
        .dout(new_Jinkela_wire_1215)
    );

    bfr new_Jinkela_buffer_1868 (
        .din(_0560_),
        .dout(new_Jinkela_wire_2957)
    );

    bfr new_Jinkela_buffer_1859 (
        .din(new_Jinkela_wire_2931),
        .dout(new_Jinkela_wire_2932)
    );

    spl2 new_Jinkela_splitter_203 (
        .a(new_Jinkela_wire_1233),
        .b(new_Jinkela_wire_1234),
        .c(new_Jinkela_wire_1235)
    );

    bfr new_Jinkela_buffer_686 (
        .din(new_Jinkela_wire_1215),
        .dout(new_Jinkela_wire_1216)
    );

    bfr new_Jinkela_buffer_1869 (
        .din(_0697_),
        .dout(new_Jinkela_wire_2958)
    );

    bfr new_Jinkela_buffer_1863 (
        .din(new_Jinkela_wire_2941),
        .dout(new_Jinkela_wire_2942)
    );

    bfr new_Jinkela_buffer_1860 (
        .din(new_Jinkela_wire_2932),
        .dout(new_Jinkela_wire_2933)
    );

    bfr new_Jinkela_buffer_687 (
        .din(new_Jinkela_wire_1216),
        .dout(new_Jinkela_wire_1217)
    );

    bfr new_Jinkela_buffer_704 (
        .din(_0240_),
        .dout(new_Jinkela_wire_1238)
    );

    bfr new_Jinkela_buffer_1861 (
        .din(new_Jinkela_wire_2933),
        .dout(new_Jinkela_wire_2934)
    );

    or_bb _1457_ (
        .a(new_Jinkela_wire_1483),
        .b(new_Jinkela_wire_1894),
        .c(_0623_)
    );

    and_bb _1458_ (
        .a(new_Jinkela_wire_1482),
        .b(new_Jinkela_wire_1893),
        .c(_0624_)
    );

    bfr new_Jinkela_buffer_1043 (
        .din(new_Jinkela_wire_1755),
        .dout(new_Jinkela_wire_1756)
    );

    spl4L new_Jinkela_splitter_275 (
        .a(new_Jinkela_wire_1737),
        .d(new_Jinkela_wire_1738),
        .e(new_Jinkela_wire_1739),
        .b(new_Jinkela_wire_1740),
        .c(new_Jinkela_wire_1741)
    );

    and_bi _1459_ (
        .a(_0623_),
        .b(_0624_),
        .c(_0625_)
    );

    spl4L new_Jinkela_splitter_276 (
        .a(new_Jinkela_wire_1742),
        .d(new_Jinkela_wire_1743),
        .e(new_Jinkela_wire_1744),
        .b(new_Jinkela_wire_1745),
        .c(new_Jinkela_wire_1746)
    );

    or_ii _1460_ (
        .a(new_Jinkela_wire_1405),
        .b(new_Jinkela_wire_2574),
        .c(_0626_)
    );

    spl4L new_Jinkela_splitter_277 (
        .a(new_Jinkela_wire_1747),
        .d(new_Jinkela_wire_1748),
        .e(new_Jinkela_wire_1749),
        .b(new_Jinkela_wire_1750),
        .c(new_Jinkela_wire_1751)
    );

    or_bb _1461_ (
        .a(new_Jinkela_wire_1404),
        .b(new_Jinkela_wire_2573),
        .c(_0627_)
    );

    bfr new_Jinkela_buffer_1042 (
        .din(new_Jinkela_wire_1754),
        .dout(new_Jinkela_wire_1755)
    );

    bfr new_Jinkela_buffer_1050 (
        .din(_0181_),
        .dout(new_Jinkela_wire_1763)
    );

    and_bb _1462_ (
        .a(_0627_),
        .b(_0626_),
        .c(_0628_)
    );

    bfr new_Jinkela_buffer_1049 (
        .din(new_Jinkela_wire_1761),
        .dout(new_Jinkela_wire_1762)
    );

    and_bi _1463_ (
        .a(_0614_),
        .b(new_Jinkela_wire_3227),
        .c(_0629_)
    );

    or_bi _1464_ (
        .a(new_Jinkela_wire_1665),
        .b(new_Jinkela_wire_1473),
        .c(_0630_)
    );

    bfr new_Jinkela_buffer_1053 (
        .din(_0707_),
        .dout(new_Jinkela_wire_1766)
    );

    bfr new_Jinkela_buffer_1044 (
        .din(new_Jinkela_wire_1756),
        .dout(new_Jinkela_wire_1757)
    );

    and_ii _1465_ (
        .a(new_Jinkela_wire_1190),
        .b(new_Jinkela_wire_1139),
        .c(_0632_)
    );

    and_bi _1466_ (
        .a(new_Jinkela_wire_500),
        .b(new_Jinkela_wire_1871),
        .c(_0633_)
    );

    bfr new_Jinkela_buffer_1051 (
        .din(new_Jinkela_wire_1763),
        .dout(new_Jinkela_wire_1764)
    );

    bfr new_Jinkela_buffer_1045 (
        .din(new_Jinkela_wire_1757),
        .dout(new_Jinkela_wire_1758)
    );

    and_bi _1467_ (
        .a(new_Jinkela_wire_671),
        .b(new_Jinkela_wire_2359),
        .c(_0634_)
    );

    or_bb _1468_ (
        .a(_0634_),
        .b(new_Jinkela_wire_3228),
        .c(_0635_)
    );

    bfr new_Jinkela_buffer_1054 (
        .din(_0227_),
        .dout(new_Jinkela_wire_1767)
    );

    bfr new_Jinkela_buffer_1046 (
        .din(new_Jinkela_wire_1758),
        .dout(new_Jinkela_wire_1759)
    );

    or_bb _1469_ (
        .a(_0635_),
        .b(new_Jinkela_wire_1505),
        .c(_0636_)
    );

    or_bi _1470_ (
        .a(new_Jinkela_wire_394),
        .b(new_Jinkela_wire_737),
        .c(_0637_)
    );

    bfr new_Jinkela_buffer_1052 (
        .din(new_Jinkela_wire_1764),
        .dout(new_Jinkela_wire_1765)
    );

    bfr new_Jinkela_buffer_1047 (
        .din(new_Jinkela_wire_1759),
        .dout(new_Jinkela_wire_1760)
    );

    and_bi _1471_ (
        .a(new_Jinkela_wire_3297),
        .b(new_Jinkela_wire_2422),
        .c(_0638_)
    );

    or_bb _1472_ (
        .a(new_Jinkela_wire_951),
        .b(_0636_),
        .c(_0639_)
    );

    spl3L new_Jinkela_splitter_279 (
        .a(new_net_7),
        .d(new_Jinkela_wire_1768),
        .b(new_Jinkela_wire_1769),
        .c(new_Jinkela_wire_1770)
    );

    bfr new_Jinkela_buffer_1076 (
        .din(_0797_),
        .dout(new_Jinkela_wire_1792)
    );

    and_bi _1473_ (
        .a(new_Jinkela_wire_1068),
        .b(new_Jinkela_wire_3008),
        .c(_0640_)
    );

    bfr new_Jinkela_buffer_1077 (
        .din(new_net_1467),
        .dout(new_Jinkela_wire_1793)
    );

    or_bb _1474_ (
        .a(_0640_),
        .b(new_Jinkela_wire_3187),
        .c(_0641_)
    );

    bfr new_Jinkela_buffer_1055 (
        .din(new_Jinkela_wire_1770),
        .dout(new_Jinkela_wire_1771)
    );

    or_bb _1475_ (
        .a(_0641_),
        .b(new_Jinkela_wire_460),
        .c(_0642_)
    );

    or_bb _1476_ (
        .a(_0642_),
        .b(new_Jinkela_wire_2725),
        .c(_0643_)
    );

    bfr new_Jinkela_buffer_1126 (
        .din(_0449_),
        .dout(new_Jinkela_wire_1842)
    );

    bfr new_Jinkela_buffer_1056 (
        .din(new_Jinkela_wire_1771),
        .dout(new_Jinkela_wire_1772)
    );

    and_ii _1477_ (
        .a(new_Jinkela_wire_233),
        .b(new_Jinkela_wire_678),
        .c(_0644_)
    );

    or_bb _1478_ (
        .a(new_Jinkela_wire_2044),
        .b(new_Jinkela_wire_1121),
        .c(_0645_)
    );

    bfr new_Jinkela_buffer_1078 (
        .din(new_Jinkela_wire_1793),
        .dout(new_Jinkela_wire_1794)
    );

    bfr new_Jinkela_buffer_1057 (
        .din(new_Jinkela_wire_1772),
        .dout(new_Jinkela_wire_1773)
    );

    and_bi _1479_ (
        .a(new_Jinkela_wire_2924),
        .b(new_Jinkela_wire_2423),
        .c(_0646_)
    );

    and_bi _1480_ (
        .a(_0645_),
        .b(new_Jinkela_wire_2036),
        .c(_0647_)
    );

    bfr new_Jinkela_buffer_1145 (
        .din(_0483_),
        .dout(new_Jinkela_wire_1861)
    );

    bfr new_Jinkela_buffer_1058 (
        .din(new_Jinkela_wire_1773),
        .dout(new_Jinkela_wire_1774)
    );

    and_bi _1481_ (
        .a(new_Jinkela_wire_322),
        .b(new_Jinkela_wire_2354),
        .c(_0648_)
    );

    and_bi _1482_ (
        .a(new_Jinkela_wire_531),
        .b(new_Jinkela_wire_1873),
        .c(_0649_)
    );

    bfr new_Jinkela_buffer_1079 (
        .din(new_Jinkela_wire_1794),
        .dout(new_Jinkela_wire_1795)
    );

    bfr new_Jinkela_buffer_1059 (
        .din(new_Jinkela_wire_1774),
        .dout(new_Jinkela_wire_1775)
    );

    or_bb _1483_ (
        .a(new_Jinkela_wire_2721),
        .b(_0648_),
        .c(_0650_)
    );

    and_bi _1484_ (
        .a(new_Jinkela_wire_2404),
        .b(new_Jinkela_wire_3003),
        .c(_0651_)
    );

    bfr new_Jinkela_buffer_1127 (
        .din(new_Jinkela_wire_1842),
        .dout(new_Jinkela_wire_1843)
    );

    bfr new_Jinkela_buffer_1060 (
        .din(new_Jinkela_wire_1775),
        .dout(new_Jinkela_wire_1776)
    );

    and_bi _1485_ (
        .a(new_Jinkela_wire_923),
        .b(new_Jinkela_wire_1750),
        .c(_0653_)
    );

    or_bb _1486_ (
        .a(_0653_),
        .b(new_Jinkela_wire_3084),
        .c(_0654_)
    );

    bfr new_Jinkela_buffer_1080 (
        .din(new_Jinkela_wire_1795),
        .dout(new_Jinkela_wire_1796)
    );

    bfr new_Jinkela_buffer_1061 (
        .din(new_Jinkela_wire_1776),
        .dout(new_Jinkela_wire_1777)
    );

    or_bb _1487_ (
        .a(new_Jinkela_wire_1733),
        .b(_0651_),
        .c(_0655_)
    );

    or_bb _1488_ (
        .a(_0655_),
        .b(new_Jinkela_wire_2117),
        .c(_0656_)
    );

    bfr new_Jinkela_buffer_1146 (
        .din(_0770_),
        .dout(new_Jinkela_wire_1862)
    );

    bfr new_Jinkela_buffer_1062 (
        .din(new_Jinkela_wire_1777),
        .dout(new_Jinkela_wire_1778)
    );

    and_bi _1489_ (
        .a(new_Jinkela_wire_1095),
        .b(_0656_),
        .c(_0657_)
    );

    spl2 new_Jinkela_splitter_281 (
        .a(_0014_),
        .b(new_Jinkela_wire_1868),
        .c(new_Jinkela_wire_1869)
    );

    and_bi _1490_ (
        .a(_0643_),
        .b(_0657_),
        .c(_0658_)
    );

    bfr new_Jinkela_buffer_1081 (
        .din(new_Jinkela_wire_1796),
        .dout(new_Jinkela_wire_1797)
    );

    bfr new_Jinkela_buffer_1063 (
        .din(new_Jinkela_wire_1778),
        .dout(new_Jinkela_wire_1779)
    );

    and_bi _1491_ (
        .a(new_Jinkela_wire_1915),
        .b(_0658_),
        .c(_0659_)
    );

    or_bb _1492_ (
        .a(_0659_),
        .b(new_Jinkela_wire_1347),
        .c(_0660_)
    );

    bfr new_Jinkela_buffer_1128 (
        .din(new_Jinkela_wire_1843),
        .dout(new_Jinkela_wire_1844)
    );

    bfr new_Jinkela_buffer_1064 (
        .din(new_Jinkela_wire_1779),
        .dout(new_Jinkela_wire_1780)
    );

    and_bi _1493_ (
        .a(_0630_),
        .b(new_Jinkela_wire_913),
        .c(_0661_)
    );

    or_bb _1494_ (
        .a(new_Jinkela_wire_1113),
        .b(_0629_),
        .c(new_net_5)
    );

    bfr new_Jinkela_buffer_1082 (
        .din(new_Jinkela_wire_1797),
        .dout(new_Jinkela_wire_1798)
    );

    bfr new_Jinkela_buffer_1065 (
        .din(new_Jinkela_wire_1780),
        .dout(new_Jinkela_wire_1781)
    );

    or_bb _1495_ (
        .a(new_Jinkela_wire_2656),
        .b(new_Jinkela_wire_1418),
        .c(_0663_)
    );

    or_bi _1496_ (
        .a(new_Jinkela_wire_1666),
        .b(new_Jinkela_wire_2063),
        .c(_0664_)
    );

    bfr new_Jinkela_buffer_1066 (
        .din(new_Jinkela_wire_1781),
        .dout(new_Jinkela_wire_1782)
    );

    and_ii _1497_ (
        .a(new_Jinkela_wire_2042),
        .b(new_Jinkela_wire_2414),
        .c(_0665_)
    );

    and_bi _1498_ (
        .a(new_Jinkela_wire_523),
        .b(new_Jinkela_wire_158),
        .c(_0666_)
    );

    bfr new_Jinkela_buffer_1083 (
        .din(new_Jinkela_wire_1798),
        .dout(new_Jinkela_wire_1799)
    );

    bfr new_Jinkela_buffer_127 (
        .din(new_Jinkela_wire_165),
        .dout(new_Jinkela_wire_166)
    );

    bfr new_Jinkela_buffer_91 (
        .din(new_Jinkela_wire_112),
        .dout(new_Jinkela_wire_113)
    );

    bfr new_Jinkela_buffer_62 (
        .din(new_Jinkela_wire_77),
        .dout(new_Jinkela_wire_78)
    );

    bfr new_Jinkela_buffer_63 (
        .din(new_Jinkela_wire_78),
        .dout(new_Jinkela_wire_79)
    );

    bfr new_Jinkela_buffer_130 (
        .din(new_Jinkela_wire_174),
        .dout(new_Jinkela_wire_175)
    );

    bfr new_Jinkela_buffer_92 (
        .din(new_Jinkela_wire_113),
        .dout(new_Jinkela_wire_114)
    );

    bfr new_Jinkela_buffer_64 (
        .din(new_Jinkela_wire_79),
        .dout(new_Jinkela_wire_80)
    );

    bfr new_Jinkela_buffer_65 (
        .din(new_Jinkela_wire_80),
        .dout(new_Jinkela_wire_81)
    );

    bfr new_Jinkela_buffer_131 (
        .din(new_Jinkela_wire_181),
        .dout(new_Jinkela_wire_182)
    );

    bfr new_Jinkela_buffer_93 (
        .din(new_Jinkela_wire_114),
        .dout(new_Jinkela_wire_115)
    );

    bfr new_Jinkela_buffer_66 (
        .din(new_Jinkela_wire_81),
        .dout(new_Jinkela_wire_82)
    );

    bfr new_Jinkela_buffer_67 (
        .din(new_Jinkela_wire_82),
        .dout(new_Jinkela_wire_83)
    );

    bfr new_Jinkela_buffer_94 (
        .din(new_Jinkela_wire_115),
        .dout(new_Jinkela_wire_116)
    );

    bfr new_Jinkela_buffer_68 (
        .din(new_Jinkela_wire_83),
        .dout(new_Jinkela_wire_84)
    );

    bfr new_Jinkela_buffer_69 (
        .din(new_Jinkela_wire_84),
        .dout(new_Jinkela_wire_85)
    );

    spl2 new_Jinkela_splitter_16 (
        .a(new_Jinkela_wire_175),
        .b(new_Jinkela_wire_176),
        .c(new_Jinkela_wire_177)
    );

    bfr new_Jinkela_buffer_95 (
        .din(new_Jinkela_wire_116),
        .dout(new_Jinkela_wire_117)
    );

    bfr new_Jinkela_buffer_70 (
        .din(new_Jinkela_wire_85),
        .dout(new_Jinkela_wire_86)
    );

    bfr new_Jinkela_buffer_71 (
        .din(new_Jinkela_wire_86),
        .dout(new_Jinkela_wire_87)
    );

    bfr new_Jinkela_buffer_132 (
        .din(new_Jinkela_wire_182),
        .dout(new_Jinkela_wire_183)
    );

    bfr new_Jinkela_buffer_96 (
        .din(new_Jinkela_wire_117),
        .dout(new_Jinkela_wire_118)
    );

    bfr new_Jinkela_buffer_72 (
        .din(new_Jinkela_wire_87),
        .dout(new_Jinkela_wire_88)
    );

    bfr new_Jinkela_buffer_73 (
        .din(new_Jinkela_wire_88),
        .dout(new_Jinkela_wire_89)
    );

    spl4L new_Jinkela_splitter_24 (
        .a(new_Jinkela_wire_211),
        .d(new_Jinkela_wire_212),
        .e(new_Jinkela_wire_213),
        .b(new_Jinkela_wire_214),
        .c(new_Jinkela_wire_216)
    );

    bfr new_Jinkela_buffer_97 (
        .din(new_Jinkela_wire_118),
        .dout(new_Jinkela_wire_119)
    );

    bfr new_Jinkela_buffer_74 (
        .din(new_Jinkela_wire_89),
        .dout(new_Jinkela_wire_90)
    );

    bfr new_Jinkela_buffer_75 (
        .din(new_Jinkela_wire_90),
        .dout(new_Jinkela_wire_91)
    );

    bfr new_Jinkela_buffer_98 (
        .din(new_Jinkela_wire_119),
        .dout(new_Jinkela_wire_120)
    );

    bfr new_Jinkela_buffer_76 (
        .din(new_Jinkela_wire_91),
        .dout(new_Jinkela_wire_92)
    );

    bfr new_Jinkela_buffer_133 (
        .din(new_Jinkela_wire_183),
        .dout(new_Jinkela_wire_184)
    );

    spl2 new_Jinkela_splitter_6 (
        .a(new_Jinkela_wire_92),
        .b(new_Jinkela_wire_93),
        .c(new_Jinkela_wire_94)
    );

    bfr new_Jinkela_buffer_138 (
        .din(new_Jinkela_wire_191),
        .dout(new_Jinkela_wire_192)
    );

    bfr new_Jinkela_buffer_99 (
        .din(new_Jinkela_wire_120),
        .dout(new_Jinkela_wire_121)
    );

    bfr new_Jinkela_buffer_100 (
        .din(new_Jinkela_wire_121),
        .dout(new_Jinkela_wire_122)
    );

    spl3L new_Jinkela_splitter_22 (
        .a(new_Jinkela_wire_197),
        .d(new_Jinkela_wire_198),
        .b(new_Jinkela_wire_199),
        .c(new_Jinkela_wire_200)
    );

    bfr new_Jinkela_buffer_134 (
        .din(new_Jinkela_wire_184),
        .dout(new_Jinkela_wire_185)
    );

    bfr new_Jinkela_buffer_101 (
        .din(new_Jinkela_wire_122),
        .dout(new_Jinkela_wire_123)
    );

    bfr new_Jinkela_buffer_102 (
        .din(new_Jinkela_wire_123),
        .dout(new_Jinkela_wire_124)
    );

    bfr new_Jinkela_buffer_155 (
        .din(G39),
        .dout(new_Jinkela_wire_232)
    );

    bfr new_Jinkela_buffer_135 (
        .din(new_Jinkela_wire_185),
        .dout(new_Jinkela_wire_186)
    );

    bfr new_Jinkela_buffer_103 (
        .din(new_Jinkela_wire_124),
        .dout(new_Jinkela_wire_125)
    );

    bfr new_Jinkela_buffer_1871 (
        .din(_0426_),
        .dout(new_Jinkela_wire_2960)
    );

    bfr new_Jinkela_buffer_1864 (
        .din(new_Jinkela_wire_2942),
        .dout(new_Jinkela_wire_2943)
    );

    spl2 new_Jinkela_splitter_416 (
        .a(new_Jinkela_wire_2934),
        .b(new_Jinkela_wire_2935),
        .c(new_Jinkela_wire_2936)
    );

    spl2 new_Jinkela_splitter_421 (
        .a(new_Jinkela_wire_2949),
        .b(new_Jinkela_wire_2950),
        .c(new_Jinkela_wire_2951)
    );

    bfr new_Jinkela_buffer_1870 (
        .din(new_Jinkela_wire_2958),
        .dout(new_Jinkela_wire_2959)
    );

    spl2 new_Jinkela_splitter_420 (
        .a(new_Jinkela_wire_2947),
        .b(new_Jinkela_wire_2948),
        .c(new_Jinkela_wire_2949)
    );

    spl2 new_Jinkela_splitter_422 (
        .a(new_Jinkela_wire_2951),
        .b(new_Jinkela_wire_2952),
        .c(new_Jinkela_wire_2953)
    );

    bfr new_Jinkela_buffer_1874 (
        .din(_0287_),
        .dout(new_Jinkela_wire_2963)
    );

    bfr new_Jinkela_buffer_1885 (
        .din(_0196_),
        .dout(new_Jinkela_wire_2991)
    );

    bfr new_Jinkela_buffer_1865 (
        .din(new_Jinkela_wire_2953),
        .dout(new_Jinkela_wire_2954)
    );

    bfr new_Jinkela_buffer_1872 (
        .din(new_Jinkela_wire_2960),
        .dout(new_Jinkela_wire_2961)
    );

    bfr new_Jinkela_buffer_1886 (
        .din(new_Jinkela_wire_2991),
        .dout(new_Jinkela_wire_2992)
    );

    bfr new_Jinkela_buffer_1866 (
        .din(new_Jinkela_wire_2954),
        .dout(new_Jinkela_wire_2955)
    );

    bfr new_Jinkela_buffer_1873 (
        .din(new_Jinkela_wire_2961),
        .dout(new_Jinkela_wire_2962)
    );

    bfr new_Jinkela_buffer_1867 (
        .din(new_Jinkela_wire_2955),
        .dout(new_Jinkela_wire_2956)
    );

    spl3L new_Jinkela_splitter_429 (
        .a(_0369_),
        .d(new_Jinkela_wire_2997),
        .b(new_Jinkela_wire_3002),
        .c(new_Jinkela_wire_3007)
    );

    bfr new_Jinkela_buffer_1887 (
        .din(_0667_),
        .dout(new_Jinkela_wire_2993)
    );

    bfr new_Jinkela_buffer_1888 (
        .din(new_Jinkela_wire_2993),
        .dout(new_Jinkela_wire_2994)
    );

    bfr new_Jinkela_buffer_1875 (
        .din(new_Jinkela_wire_2963),
        .dout(new_Jinkela_wire_2964)
    );

    spl3L new_Jinkela_splitter_423 (
        .a(new_Jinkela_wire_2964),
        .d(new_Jinkela_wire_2965),
        .b(new_Jinkela_wire_2966),
        .c(new_Jinkela_wire_2969)
    );

    spl2 new_Jinkela_splitter_426 (
        .a(new_Jinkela_wire_2973),
        .b(new_Jinkela_wire_2974),
        .c(new_Jinkela_wire_2977)
    );

    spl2 new_Jinkela_splitter_424 (
        .a(new_Jinkela_wire_2966),
        .b(new_Jinkela_wire_2967),
        .c(new_Jinkela_wire_2968)
    );

    spl4L new_Jinkela_splitter_425 (
        .a(new_Jinkela_wire_2969),
        .d(new_Jinkela_wire_2970),
        .e(new_Jinkela_wire_2971),
        .b(new_Jinkela_wire_2972),
        .c(new_Jinkela_wire_2973)
    );

    spl2 new_Jinkela_splitter_433 (
        .a(_0766_),
        .b(new_Jinkela_wire_3012),
        .c(new_Jinkela_wire_3013)
    );

    bfr new_Jinkela_buffer_1889 (
        .din(new_Jinkela_wire_2994),
        .dout(new_Jinkela_wire_2995)
    );

    spl4L new_Jinkela_splitter_428 (
        .a(new_Jinkela_wire_2977),
        .d(new_Jinkela_wire_2978),
        .e(new_Jinkela_wire_2979),
        .b(new_Jinkela_wire_2980),
        .c(new_Jinkela_wire_2981)
    );

    spl2 new_Jinkela_splitter_427 (
        .a(new_Jinkela_wire_2974),
        .b(new_Jinkela_wire_2975),
        .c(new_Jinkela_wire_2976)
    );

    bfr new_Jinkela_buffer_1876 (
        .din(new_Jinkela_wire_2981),
        .dout(new_Jinkela_wire_2982)
    );

    spl4L new_Jinkela_splitter_431 (
        .a(new_Jinkela_wire_3002),
        .d(new_Jinkela_wire_3003),
        .e(new_Jinkela_wire_3004),
        .b(new_Jinkela_wire_3005),
        .c(new_Jinkela_wire_3006)
    );

    bfr new_Jinkela_buffer_1890 (
        .din(new_Jinkela_wire_2995),
        .dout(new_Jinkela_wire_2996)
    );

    bfr new_Jinkela_buffer_1877 (
        .din(new_Jinkela_wire_2982),
        .dout(new_Jinkela_wire_2983)
    );

    bfr new_Jinkela_buffer_1893 (
        .din(_0579_),
        .dout(new_Jinkela_wire_3019)
    );

    spl4L new_Jinkela_splitter_430 (
        .a(new_Jinkela_wire_2997),
        .d(new_Jinkela_wire_2998),
        .e(new_Jinkela_wire_2999),
        .b(new_Jinkela_wire_3000),
        .c(new_Jinkela_wire_3001)
    );

    bfr new_Jinkela_buffer_1878 (
        .din(new_Jinkela_wire_2983),
        .dout(new_Jinkela_wire_2984)
    );

    bfr new_Jinkela_buffer_1891 (
        .din(new_Jinkela_wire_3016),
        .dout(new_Jinkela_wire_3017)
    );

    bfr new_Jinkela_buffer_1879 (
        .din(new_Jinkela_wire_2984),
        .dout(new_Jinkela_wire_2985)
    );

    spl4L new_Jinkela_splitter_432 (
        .a(new_Jinkela_wire_3007),
        .d(new_Jinkela_wire_3008),
        .e(new_Jinkela_wire_3009),
        .b(new_Jinkela_wire_3010),
        .c(new_Jinkela_wire_3011)
    );

    bfr new_Jinkela_buffer_1880 (
        .din(new_Jinkela_wire_2985),
        .dout(new_Jinkela_wire_2986)
    );

    bfr new_Jinkela_buffer_1892 (
        .din(_0589_),
        .dout(new_Jinkela_wire_3018)
    );

    spl3L new_Jinkela_splitter_434 (
        .a(_0164_),
        .d(new_Jinkela_wire_3014),
        .b(new_Jinkela_wire_3015),
        .c(new_Jinkela_wire_3016)
    );

    bfr new_Jinkela_buffer_1881 (
        .din(new_Jinkela_wire_2986),
        .dout(new_Jinkela_wire_2987)
    );

    bfr new_Jinkela_buffer_1882 (
        .din(new_Jinkela_wire_2987),
        .dout(new_Jinkela_wire_2988)
    );

    bfr new_Jinkela_buffer_1067 (
        .din(new_Jinkela_wire_1782),
        .dout(new_Jinkela_wire_1783)
    );

    bfr new_Jinkela_buffer_1129 (
        .din(new_Jinkela_wire_1844),
        .dout(new_Jinkela_wire_1845)
    );

    bfr new_Jinkela_buffer_1068 (
        .din(new_Jinkela_wire_1783),
        .dout(new_Jinkela_wire_1784)
    );

    bfr new_Jinkela_buffer_1084 (
        .din(new_Jinkela_wire_1799),
        .dout(new_Jinkela_wire_1800)
    );

    bfr new_Jinkela_buffer_1069 (
        .din(new_Jinkela_wire_1784),
        .dout(new_Jinkela_wire_1785)
    );

    spl4L new_Jinkela_splitter_282 (
        .a(_0372_),
        .d(new_Jinkela_wire_1870),
        .e(new_Jinkela_wire_1875),
        .b(new_Jinkela_wire_1880),
        .c(new_Jinkela_wire_1885)
    );

    bfr new_Jinkela_buffer_1070 (
        .din(new_Jinkela_wire_1785),
        .dout(new_Jinkela_wire_1786)
    );

    spl2 new_Jinkela_splitter_280 (
        .a(new_Jinkela_wire_1862),
        .b(new_Jinkela_wire_1863),
        .c(new_Jinkela_wire_1864)
    );

    bfr new_Jinkela_buffer_1085 (
        .din(new_Jinkela_wire_1800),
        .dout(new_Jinkela_wire_1801)
    );

    bfr new_Jinkela_buffer_1071 (
        .din(new_Jinkela_wire_1786),
        .dout(new_Jinkela_wire_1787)
    );

    bfr new_Jinkela_buffer_1130 (
        .din(new_Jinkela_wire_1845),
        .dout(new_Jinkela_wire_1846)
    );

    bfr new_Jinkela_buffer_1072 (
        .din(new_Jinkela_wire_1787),
        .dout(new_Jinkela_wire_1788)
    );

    bfr new_Jinkela_buffer_1086 (
        .din(new_Jinkela_wire_1801),
        .dout(new_Jinkela_wire_1802)
    );

    bfr new_Jinkela_buffer_1073 (
        .din(new_Jinkela_wire_1788),
        .dout(new_Jinkela_wire_1789)
    );

    bfr new_Jinkela_buffer_1074 (
        .din(new_Jinkela_wire_1789),
        .dout(new_Jinkela_wire_1790)
    );

    bfr new_Jinkela_buffer_1147 (
        .din(new_Jinkela_wire_1864),
        .dout(new_Jinkela_wire_1865)
    );

    bfr new_Jinkela_buffer_1087 (
        .din(new_Jinkela_wire_1802),
        .dout(new_Jinkela_wire_1803)
    );

    bfr new_Jinkela_buffer_1075 (
        .din(new_Jinkela_wire_1790),
        .dout(new_Jinkela_wire_1791)
    );

    bfr new_Jinkela_buffer_1131 (
        .din(new_Jinkela_wire_1846),
        .dout(new_Jinkela_wire_1847)
    );

    bfr new_Jinkela_buffer_1088 (
        .din(new_Jinkela_wire_1803),
        .dout(new_Jinkela_wire_1804)
    );

    bfr new_Jinkela_buffer_1089 (
        .din(new_Jinkela_wire_1804),
        .dout(new_Jinkela_wire_1805)
    );

    bfr new_Jinkela_buffer_1132 (
        .din(new_Jinkela_wire_1847),
        .dout(new_Jinkela_wire_1848)
    );

    bfr new_Jinkela_buffer_1090 (
        .din(new_Jinkela_wire_1805),
        .dout(new_Jinkela_wire_1806)
    );

    spl2 new_Jinkela_splitter_288 (
        .a(_0616_),
        .b(new_Jinkela_wire_1893),
        .c(new_Jinkela_wire_1894)
    );

    bfr new_Jinkela_buffer_1091 (
        .din(new_Jinkela_wire_1806),
        .dout(new_Jinkela_wire_1807)
    );

    bfr new_Jinkela_buffer_1133 (
        .din(new_Jinkela_wire_1848),
        .dout(new_Jinkela_wire_1849)
    );

    bfr new_Jinkela_buffer_1092 (
        .din(new_Jinkela_wire_1807),
        .dout(new_Jinkela_wire_1808)
    );

    spl3L new_Jinkela_splitter_287 (
        .a(_0260_),
        .d(new_Jinkela_wire_1890),
        .b(new_Jinkela_wire_1891),
        .c(new_Jinkela_wire_1892)
    );

    bfr new_Jinkela_buffer_1148 (
        .din(new_Jinkela_wire_1865),
        .dout(new_Jinkela_wire_1866)
    );

    bfr new_Jinkela_buffer_1093 (
        .din(new_Jinkela_wire_1808),
        .dout(new_Jinkela_wire_1809)
    );

    bfr new_Jinkela_buffer_1134 (
        .din(new_Jinkela_wire_1849),
        .dout(new_Jinkela_wire_1850)
    );

    bfr new_Jinkela_buffer_1094 (
        .din(new_Jinkela_wire_1809),
        .dout(new_Jinkela_wire_1810)
    );

    bfr new_Jinkela_buffer_1095 (
        .din(new_Jinkela_wire_1810),
        .dout(new_Jinkela_wire_1811)
    );

    bfr new_Jinkela_buffer_1135 (
        .din(new_Jinkela_wire_1850),
        .dout(new_Jinkela_wire_1851)
    );

    bfr new_Jinkela_buffer_1096 (
        .din(new_Jinkela_wire_1811),
        .dout(new_Jinkela_wire_1812)
    );

    bfr new_Jinkela_buffer_1150 (
        .din(_0359_),
        .dout(new_Jinkela_wire_1895)
    );

    bfr new_Jinkela_buffer_1149 (
        .din(new_Jinkela_wire_1866),
        .dout(new_Jinkela_wire_1867)
    );

    bfr new_Jinkela_buffer_1097 (
        .din(new_Jinkela_wire_1812),
        .dout(new_Jinkela_wire_1813)
    );

    bfr new_Jinkela_buffer_1136 (
        .din(new_Jinkela_wire_1851),
        .dout(new_Jinkela_wire_1852)
    );

    bfr new_Jinkela_buffer_1098 (
        .din(new_Jinkela_wire_1813),
        .dout(new_Jinkela_wire_1814)
    );

    spl4L new_Jinkela_splitter_284 (
        .a(new_Jinkela_wire_1875),
        .d(new_Jinkela_wire_1876),
        .e(new_Jinkela_wire_1877),
        .b(new_Jinkela_wire_1878),
        .c(new_Jinkela_wire_1879)
    );

    bfr new_Jinkela_buffer_1099 (
        .din(new_Jinkela_wire_1814),
        .dout(new_Jinkela_wire_1815)
    );

    bfr new_Jinkela_buffer_1137 (
        .din(new_Jinkela_wire_1852),
        .dout(new_Jinkela_wire_1853)
    );

    and_bb _1121_ (
        .a(new_Jinkela_wire_2275),
        .b(new_Jinkela_wire_1038),
        .c(_0292_)
    );

    or_ii _1122_ (
        .a(new_Jinkela_wire_1205),
        .b(new_Jinkela_wire_659),
        .c(_0293_)
    );

    or_bi _1123_ (
        .a(new_Jinkela_wire_837),
        .b(new_Jinkela_wire_2587),
        .c(_0294_)
    );

    and_bi _1124_ (
        .a(_0292_),
        .b(_0294_),
        .c(_0295_)
    );

    and_bi _1125_ (
        .a(new_Jinkela_wire_2829),
        .b(_0295_),
        .c(_0296_)
    );

    and_bi _1126_ (
        .a(new_Jinkela_wire_2976),
        .b(_0296_),
        .c(_0297_)
    );

    and_bi _1127_ (
        .a(new_Jinkela_wire_2563),
        .b(new_Jinkela_wire_2276),
        .c(_0298_)
    );

    and_bi _1128_ (
        .a(new_Jinkela_wire_1892),
        .b(_0298_),
        .c(_0299_)
    );

    and_bi _1129_ (
        .a(new_Jinkela_wire_1753),
        .b(new_Jinkela_wire_917),
        .c(_0300_)
    );

    inv _1130_ (
        .din(new_Jinkela_wire_1144),
        .dout(_0301_)
    );

    or_bb _1131_ (
        .a(new_Jinkela_wire_1098),
        .b(new_Jinkela_wire_2937),
        .c(_0302_)
    );

    and_bi _1132_ (
        .a(new_Jinkela_wire_2207),
        .b(new_Jinkela_wire_1725),
        .c(_0303_)
    );

    or_bb _1133_ (
        .a(_0303_),
        .b(new_Jinkela_wire_2841),
        .c(_0304_)
    );

    and_bi _1134_ (
        .a(new_Jinkela_wire_33),
        .b(new_Jinkela_wire_2319),
        .c(_0305_)
    );

    or_bb _1135_ (
        .a(new_Jinkela_wire_2967),
        .b(new_Jinkela_wire_2448),
        .c(_0306_)
    );

    and_bi _1136_ (
        .a(new_Jinkela_wire_3099),
        .b(new_Jinkela_wire_1981),
        .c(_0307_)
    );

    and_bi _1137_ (
        .a(new_Jinkela_wire_1982),
        .b(new_Jinkela_wire_3098),
        .c(_0308_)
    );

    and_ii _1138_ (
        .a(_0308_),
        .b(_0307_),
        .c(_0309_)
    );

    and_bi _1139_ (
        .a(new_Jinkela_wire_1263),
        .b(new_Jinkela_wire_2965),
        .c(_0310_)
    );

    and_bi _1140_ (
        .a(new_Jinkela_wire_1630),
        .b(new_Jinkela_wire_3199),
        .c(_0311_)
    );

    and_bi _1141_ (
        .a(new_Jinkela_wire_3198),
        .b(new_Jinkela_wire_1629),
        .c(_0312_)
    );

    or_bb _1142_ (
        .a(_0312_),
        .b(_0311_),
        .c(_0313_)
    );

    or_bb _1143_ (
        .a(new_Jinkela_wire_3067),
        .b(new_Jinkela_wire_1074),
        .c(_0314_)
    );

    or_ii _1144_ (
        .a(new_Jinkela_wire_3232),
        .b(new_Jinkela_wire_102),
        .c(_0315_)
    );

    and_bi _1145_ (
        .a(new_Jinkela_wire_1290),
        .b(new_Jinkela_wire_2500),
        .c(_0316_)
    );

    or_bb _1146_ (
        .a(new_Jinkela_wire_1363),
        .b(new_Jinkela_wire_1366),
        .c(_0317_)
    );

    and_bb _1147_ (
        .a(new_Jinkela_wire_1362),
        .b(new_Jinkela_wire_1365),
        .c(_0318_)
    );

    and_bi _1148_ (
        .a(_0317_),
        .b(_0318_),
        .c(_0319_)
    );

    inv _1149_ (
        .din(new_Jinkela_wire_3209),
        .dout(_0320_)
    );

    and_ii _1150_ (
        .a(new_Jinkela_wire_3178),
        .b(new_Jinkela_wire_2323),
        .c(_0321_)
    );

    or_ii _1151_ (
        .a(new_Jinkela_wire_959),
        .b(new_Jinkela_wire_971),
        .c(_0322_)
    );

    or_bi _1152_ (
        .a(new_Jinkela_wire_2331),
        .b(new_Jinkela_wire_974),
        .c(_0323_)
    );

    and_bb _1153_ (
        .a(new_Jinkela_wire_2975),
        .b(new_Jinkela_wire_3015),
        .c(_0324_)
    );

    and_bb _1154_ (
        .a(new_Jinkela_wire_2980),
        .b(new_Jinkela_wire_2880),
        .c(_0325_)
    );

    and_ii _1155_ (
        .a(new_Jinkela_wire_3238),
        .b(new_Jinkela_wire_1075),
        .c(_0326_)
    );

    and_ii _1156_ (
        .a(_0326_),
        .b(new_Jinkela_wire_2440),
        .c(_0327_)
    );

    and_bi _1157_ (
        .a(new_Jinkela_wire_3214),
        .b(new_Jinkela_wire_941),
        .c(_0328_)
    );

    and_bi _1158_ (
        .a(new_Jinkela_wire_940),
        .b(new_Jinkela_wire_3213),
        .c(_0329_)
    );

    or_bb _1159_ (
        .a(new_Jinkela_wire_2875),
        .b(new_Jinkela_wire_961),
        .c(_0330_)
    );

    and_bi _1160_ (
        .a(new_Jinkela_wire_1489),
        .b(new_Jinkela_wire_1328),
        .c(_0331_)
    );

    and_bi _1161_ (
        .a(new_Jinkela_wire_2738),
        .b(_0331_),
        .c(_0332_)
    );

    or_bb _1162_ (
        .a(new_Jinkela_wire_1402),
        .b(new_Jinkela_wire_3258),
        .c(_0333_)
    );

    bfr new_Jinkela_buffer_1100 (
        .din(new_Jinkela_wire_1815),
        .dout(new_Jinkela_wire_1816)
    );

    bfr new_Jinkela_buffer_1899 (
        .din(_0739_),
        .dout(new_Jinkela_wire_3025)
    );

    spl2 new_Jinkela_splitter_293 (
        .a(_0367_),
        .b(new_Jinkela_wire_1924),
        .c(new_Jinkela_wire_1925)
    );

    bfr new_Jinkela_buffer_1883 (
        .din(new_Jinkela_wire_2988),
        .dout(new_Jinkela_wire_2989)
    );

    bfr new_Jinkela_buffer_1101 (
        .din(new_Jinkela_wire_1816),
        .dout(new_Jinkela_wire_1817)
    );

    bfr new_Jinkela_buffer_1894 (
        .din(new_Jinkela_wire_3019),
        .dout(new_Jinkela_wire_3020)
    );

    bfr new_Jinkela_buffer_1138 (
        .din(new_Jinkela_wire_1853),
        .dout(new_Jinkela_wire_1854)
    );

    bfr new_Jinkela_buffer_1884 (
        .din(new_Jinkela_wire_2989),
        .dout(new_Jinkela_wire_2990)
    );

    bfr new_Jinkela_buffer_1102 (
        .din(new_Jinkela_wire_1817),
        .dout(new_Jinkela_wire_1818)
    );

    spl2 new_Jinkela_splitter_435 (
        .a(_0074_),
        .b(new_Jinkela_wire_3026),
        .c(new_Jinkela_wire_3031)
    );

    bfr new_Jinkela_buffer_1895 (
        .din(new_Jinkela_wire_3020),
        .dout(new_Jinkela_wire_3021)
    );

    spl4L new_Jinkela_splitter_283 (
        .a(new_Jinkela_wire_1870),
        .d(new_Jinkela_wire_1871),
        .e(new_Jinkela_wire_1872),
        .b(new_Jinkela_wire_1873),
        .c(new_Jinkela_wire_1874)
    );

    bfr new_Jinkela_buffer_1103 (
        .din(new_Jinkela_wire_1818),
        .dout(new_Jinkela_wire_1819)
    );

    spl4L new_Jinkela_splitter_436 (
        .a(new_Jinkela_wire_3026),
        .d(new_Jinkela_wire_3027),
        .e(new_Jinkela_wire_3028),
        .b(new_Jinkela_wire_3029),
        .c(new_Jinkela_wire_3030)
    );

    bfr new_Jinkela_buffer_1139 (
        .din(new_Jinkela_wire_1854),
        .dout(new_Jinkela_wire_1855)
    );

    bfr new_Jinkela_buffer_1896 (
        .din(new_Jinkela_wire_3021),
        .dout(new_Jinkela_wire_3022)
    );

    bfr new_Jinkela_buffer_1104 (
        .din(new_Jinkela_wire_1819),
        .dout(new_Jinkela_wire_1820)
    );

    spl2 new_Jinkela_splitter_438 (
        .a(_0555_),
        .b(new_Jinkela_wire_3037),
        .c(new_Jinkela_wire_3038)
    );

    bfr new_Jinkela_buffer_1163 (
        .din(new_Jinkela_wire_1919),
        .dout(new_Jinkela_wire_1920)
    );

    bfr new_Jinkela_buffer_1897 (
        .din(new_Jinkela_wire_3022),
        .dout(new_Jinkela_wire_3023)
    );

    spl4L new_Jinkela_splitter_285 (
        .a(new_Jinkela_wire_1880),
        .d(new_Jinkela_wire_1881),
        .e(new_Jinkela_wire_1882),
        .b(new_Jinkela_wire_1883),
        .c(new_Jinkela_wire_1884)
    );

    bfr new_Jinkela_buffer_1105 (
        .din(new_Jinkela_wire_1820),
        .dout(new_Jinkela_wire_1821)
    );

    bfr new_Jinkela_buffer_1904 (
        .din(_0204_),
        .dout(new_Jinkela_wire_3042)
    );

    bfr new_Jinkela_buffer_1905 (
        .din(_0134_),
        .dout(new_Jinkela_wire_3043)
    );

    bfr new_Jinkela_buffer_1140 (
        .din(new_Jinkela_wire_1855),
        .dout(new_Jinkela_wire_1856)
    );

    bfr new_Jinkela_buffer_1898 (
        .din(new_Jinkela_wire_3023),
        .dout(new_Jinkela_wire_3024)
    );

    bfr new_Jinkela_buffer_1106 (
        .din(new_Jinkela_wire_1821),
        .dout(new_Jinkela_wire_1822)
    );

    spl4L new_Jinkela_splitter_437 (
        .a(new_Jinkela_wire_3031),
        .d(new_Jinkela_wire_3032),
        .e(new_Jinkela_wire_3033),
        .b(new_Jinkela_wire_3034),
        .c(new_Jinkela_wire_3035)
    );

    bfr new_Jinkela_buffer_1900 (
        .din(_0781_),
        .dout(new_Jinkela_wire_3036)
    );

    spl4L new_Jinkela_splitter_286 (
        .a(new_Jinkela_wire_1885),
        .d(new_Jinkela_wire_1886),
        .e(new_Jinkela_wire_1887),
        .b(new_Jinkela_wire_1888),
        .c(new_Jinkela_wire_1889)
    );

    bfr new_Jinkela_buffer_1107 (
        .din(new_Jinkela_wire_1822),
        .dout(new_Jinkela_wire_1823)
    );

    bfr new_Jinkela_buffer_1901 (
        .din(new_Jinkela_wire_3038),
        .dout(new_Jinkela_wire_3039)
    );

    bfr new_Jinkela_buffer_1141 (
        .din(new_Jinkela_wire_1856),
        .dout(new_Jinkela_wire_1857)
    );

    bfr new_Jinkela_buffer_1108 (
        .din(new_Jinkela_wire_1823),
        .dout(new_Jinkela_wire_1824)
    );

    bfr new_Jinkela_buffer_1906 (
        .din(_0101_),
        .dout(new_Jinkela_wire_3044)
    );

    bfr new_Jinkela_buffer_1902 (
        .din(new_Jinkela_wire_3039),
        .dout(new_Jinkela_wire_3040)
    );

    bfr new_Jinkela_buffer_1109 (
        .din(new_Jinkela_wire_1824),
        .dout(new_Jinkela_wire_1825)
    );

    bfr new_Jinkela_buffer_1907 (
        .din(_0387_),
        .dout(new_Jinkela_wire_3045)
    );

    bfr new_Jinkela_buffer_1903 (
        .din(new_Jinkela_wire_3040),
        .dout(new_Jinkela_wire_3041)
    );

    bfr new_Jinkela_buffer_1142 (
        .din(new_Jinkela_wire_1857),
        .dout(new_Jinkela_wire_1858)
    );

    bfr new_Jinkela_buffer_1110 (
        .din(new_Jinkela_wire_1825),
        .dout(new_Jinkela_wire_1826)
    );

    bfr new_Jinkela_buffer_1909 (
        .din(_0514_),
        .dout(new_Jinkela_wire_3047)
    );

    bfr new_Jinkela_buffer_1908 (
        .din(new_Jinkela_wire_3045),
        .dout(new_Jinkela_wire_3046)
    );

    spl2 new_Jinkela_splitter_292 (
        .a(_0384_),
        .b(new_Jinkela_wire_1918),
        .c(new_Jinkela_wire_1919)
    );

    bfr new_Jinkela_buffer_1111 (
        .din(new_Jinkela_wire_1826),
        .dout(new_Jinkela_wire_1827)
    );

    bfr new_Jinkela_buffer_1910 (
        .din(_0085_),
        .dout(new_Jinkela_wire_3048)
    );

    spl2 new_Jinkela_splitter_445 (
        .a(_0382_),
        .b(new_Jinkela_wire_3080),
        .c(new_Jinkela_wire_3081)
    );

    bfr new_Jinkela_buffer_1143 (
        .din(new_Jinkela_wire_1858),
        .dout(new_Jinkela_wire_1859)
    );

    bfr new_Jinkela_buffer_1112 (
        .din(new_Jinkela_wire_1827),
        .dout(new_Jinkela_wire_1828)
    );

    spl3L new_Jinkela_splitter_443 (
        .a(_0313_),
        .d(new_Jinkela_wire_3067),
        .b(new_Jinkela_wire_3068),
        .c(new_Jinkela_wire_3069)
    );

    bfr new_Jinkela_buffer_1162 (
        .din(_0421_),
        .dout(new_Jinkela_wire_1917)
    );

    bfr new_Jinkela_buffer_1926 (
        .din(new_Jinkela_wire_3081),
        .dout(new_Jinkela_wire_3082)
    );

    bfr new_Jinkela_buffer_1151 (
        .din(new_Jinkela_wire_1895),
        .dout(new_Jinkela_wire_1896)
    );

    bfr new_Jinkela_buffer_1113 (
        .din(new_Jinkela_wire_1828),
        .dout(new_Jinkela_wire_1829)
    );

    bfr new_Jinkela_buffer_1911 (
        .din(new_Jinkela_wire_3048),
        .dout(new_Jinkela_wire_3049)
    );

    bfr new_Jinkela_buffer_1144 (
        .din(new_Jinkela_wire_1859),
        .dout(new_Jinkela_wire_1860)
    );

    bfr new_Jinkela_buffer_1918 (
        .din(new_Jinkela_wire_3069),
        .dout(new_Jinkela_wire_3070)
    );

    bfr new_Jinkela_buffer_1114 (
        .din(new_Jinkela_wire_1829),
        .dout(new_Jinkela_wire_1830)
    );

    bfr new_Jinkela_buffer_1912 (
        .din(new_Jinkela_wire_3049),
        .dout(new_Jinkela_wire_3050)
    );

    bfr new_Jinkela_buffer_1913 (
        .din(new_Jinkela_wire_3050),
        .dout(new_Jinkela_wire_3051)
    );

    bfr new_Jinkela_buffer_1914 (
        .din(new_Jinkela_wire_3051),
        .dout(new_Jinkela_wire_3052)
    );

    bfr new_Jinkela_buffer_1115 (
        .din(new_Jinkela_wire_1830),
        .dout(new_Jinkela_wire_1831)
    );

    bfr new_Jinkela_buffer_1930 (
        .din(_0669_),
        .dout(new_Jinkela_wire_3094)
    );

    bfr new_Jinkela_buffer_1929 (
        .din(_0790_),
        .dout(new_Jinkela_wire_3093)
    );

    bfr new_Jinkela_buffer_1932 (
        .din(_0306_),
        .dout(new_Jinkela_wire_3096)
    );

    bfr new_Jinkela_buffer_1152 (
        .din(new_Jinkela_wire_1896),
        .dout(new_Jinkela_wire_1897)
    );

    bfr new_Jinkela_buffer_1116 (
        .din(new_Jinkela_wire_1831),
        .dout(new_Jinkela_wire_1832)
    );

    bfr new_Jinkela_buffer_1919 (
        .din(new_Jinkela_wire_3070),
        .dout(new_Jinkela_wire_3071)
    );

    bfr new_Jinkela_buffer_1117 (
        .din(new_Jinkela_wire_1832),
        .dout(new_Jinkela_wire_1833)
    );

    bfr new_Jinkela_buffer_1915 (
        .din(new_Jinkela_wire_3052),
        .dout(new_Jinkela_wire_3053)
    );

    bfr new_Jinkela_buffer_1154 (
        .din(new_Jinkela_wire_1898),
        .dout(new_Jinkela_wire_1899)
    );

    bfr new_Jinkela_buffer_1920 (
        .din(new_Jinkela_wire_3071),
        .dout(new_Jinkela_wire_3072)
    );

    bfr new_Jinkela_buffer_1118 (
        .din(new_Jinkela_wire_1833),
        .dout(new_Jinkela_wire_1834)
    );

    bfr new_Jinkela_buffer_1916 (
        .din(new_Jinkela_wire_3053),
        .dout(new_Jinkela_wire_3054)
    );

    bfr new_Jinkela_buffer_1167 (
        .din(_0745_),
        .dout(new_Jinkela_wire_1926)
    );

    bfr new_Jinkela_buffer_1168 (
        .din(_0042_),
        .dout(new_Jinkela_wire_1927)
    );

    bfr new_Jinkela_buffer_1934 (
        .din(new_net_1465),
        .dout(new_Jinkela_wire_3100)
    );

    bfr new_Jinkela_buffer_1119 (
        .din(new_Jinkela_wire_1834),
        .dout(new_Jinkela_wire_1835)
    );

    bfr new_Jinkela_buffer_1917 (
        .din(new_Jinkela_wire_3054),
        .dout(new_Jinkela_wire_3055)
    );

    bfr new_Jinkela_buffer_1921 (
        .din(new_Jinkela_wire_3072),
        .dout(new_Jinkela_wire_3073)
    );

    bfr new_Jinkela_buffer_1120 (
        .din(new_Jinkela_wire_1835),
        .dout(new_Jinkela_wire_1836)
    );

    spl2 new_Jinkela_splitter_439 (
        .a(new_Jinkela_wire_3055),
        .b(new_Jinkela_wire_3056),
        .c(new_Jinkela_wire_3057)
    );

    bfr new_Jinkela_buffer_1153 (
        .din(new_Jinkela_wire_1897),
        .dout(new_Jinkela_wire_1898)
    );

    spl2 new_Jinkela_splitter_440 (
        .a(new_Jinkela_wire_3057),
        .b(new_Jinkela_wire_3058),
        .c(new_Jinkela_wire_3062)
    );

    or_bb _1499_ (
        .a(new_Jinkela_wire_1706),
        .b(new_Jinkela_wire_3080),
        .c(_0667_)
    );

    bfr new_Jinkela_buffer_104 (
        .din(new_Jinkela_wire_125),
        .dout(new_Jinkela_wire_126)
    );

    or_bb _1500_ (
        .a(new_Jinkela_wire_2996),
        .b(_0665_),
        .c(_0668_)
    );

    bfr new_Jinkela_buffer_136 (
        .din(new_Jinkela_wire_186),
        .dout(new_Jinkela_wire_187)
    );

    and_bi _1501_ (
        .a(new_Jinkela_wire_722),
        .b(new_Jinkela_wire_1749),
        .c(_0669_)
    );

    bfr new_Jinkela_buffer_105 (
        .din(new_Jinkela_wire_126),
        .dout(new_Jinkela_wire_127)
    );

    and_bi _1502_ (
        .a(new_Jinkela_wire_698),
        .b(new_Jinkela_wire_1872),
        .c(_0670_)
    );

    bfr new_Jinkela_buffer_139 (
        .din(new_Jinkela_wire_200),
        .dout(new_Jinkela_wire_201)
    );

    or_bb _1503_ (
        .a(_0670_),
        .b(new_Jinkela_wire_3095),
        .c(_0671_)
    );

    bfr new_Jinkela_buffer_106 (
        .din(new_Jinkela_wire_127),
        .dout(new_Jinkela_wire_128)
    );

    and_ii _1504_ (
        .a(new_Jinkela_wire_520),
        .b(new_Jinkela_wire_787),
        .c(_0672_)
    );

    spl2 new_Jinkela_splitter_19 (
        .a(new_Jinkela_wire_187),
        .b(new_Jinkela_wire_188),
        .c(new_Jinkela_wire_189)
    );

    and_ii _1505_ (
        .a(new_Jinkela_wire_1301),
        .b(new_Jinkela_wire_2356),
        .c(_0674_)
    );

    bfr new_Jinkela_buffer_107 (
        .din(new_Jinkela_wire_128),
        .dout(new_Jinkela_wire_129)
    );

    or_bb _1506_ (
        .a(new_Jinkela_wire_274),
        .b(new_Jinkela_wire_311),
        .c(_0675_)
    );

    bfr new_Jinkela_buffer_137 (
        .din(new_Jinkela_wire_189),
        .dout(new_Jinkela_wire_190)
    );

    and_bi _1507_ (
        .a(new_Jinkela_wire_984),
        .b(new_Jinkela_wire_1126),
        .c(_0676_)
    );

    bfr new_Jinkela_buffer_108 (
        .din(new_Jinkela_wire_129),
        .dout(new_Jinkela_wire_130)
    );

    or_bb _1508_ (
        .a(_0676_),
        .b(_0674_),
        .c(_0677_)
    );

    bfr new_Jinkela_buffer_147 (
        .din(new_Jinkela_wire_209),
        .dout(new_Jinkela_wire_210)
    );

    or_bb _1509_ (
        .a(_0677_),
        .b(new_Jinkela_wire_2408),
        .c(_0678_)
    );

    bfr new_Jinkela_buffer_109 (
        .din(new_Jinkela_wire_130),
        .dout(new_Jinkela_wire_131)
    );

    or_bb _1510_ (
        .a(_0678_),
        .b(new_Jinkela_wire_1275),
        .c(_0679_)
    );

    bfr new_Jinkela_buffer_140 (
        .din(new_Jinkela_wire_201),
        .dout(new_Jinkela_wire_202)
    );

    and_ii _1511_ (
        .a(new_Jinkela_wire_1923),
        .b(new_Jinkela_wire_1569),
        .c(_0680_)
    );

    bfr new_Jinkela_buffer_110 (
        .din(new_Jinkela_wire_131),
        .dout(new_Jinkela_wire_132)
    );

    and_bi _1512_ (
        .a(new_Jinkela_wire_1693),
        .b(new_Jinkela_wire_2358),
        .c(_0681_)
    );

    spl4L new_Jinkela_splitter_25 (
        .a(new_Jinkela_wire_216),
        .d(new_Jinkela_wire_217),
        .e(new_Jinkela_wire_218),
        .b(new_Jinkela_wire_219),
        .c(new_Jinkela_wire_220)
    );

    or_bb _1513_ (
        .a(_0681_),
        .b(new_Jinkela_wire_2578),
        .c(_0682_)
    );

    bfr new_Jinkela_buffer_111 (
        .din(new_Jinkela_wire_132),
        .dout(new_Jinkela_wire_133)
    );

    and_bi _1514_ (
        .a(new_Jinkela_wire_2765),
        .b(new_Jinkela_wire_1117),
        .c(_0683_)
    );

    spl4L new_Jinkela_splitter_37 (
        .a(new_Jinkela_wire_265),
        .d(new_Jinkela_wire_266),
        .e(new_Jinkela_wire_267),
        .b(new_Jinkela_wire_268),
        .c(new_Jinkela_wire_269)
    );

    bfr new_Jinkela_buffer_141 (
        .din(new_Jinkela_wire_202),
        .dout(new_Jinkela_wire_203)
    );

    and_bi _1515_ (
        .a(new_Jinkela_wire_1060),
        .b(new_Jinkela_wire_1879),
        .c(_0685_)
    );

    bfr new_Jinkela_buffer_112 (
        .din(new_Jinkela_wire_133),
        .dout(new_Jinkela_wire_134)
    );

    or_bb _1516_ (
        .a(new_Jinkela_wire_833),
        .b(_0683_),
        .c(_0686_)
    );

    or_bb _1517_ (
        .a(_0686_),
        .b(_0682_),
        .c(_0687_)
    );

    bfr new_Jinkela_buffer_113 (
        .din(new_Jinkela_wire_134),
        .dout(new_Jinkela_wire_135)
    );

    or_bb _1518_ (
        .a(new_Jinkela_wire_2378),
        .b(new_Jinkela_wire_1643),
        .c(_0688_)
    );

    spl2 new_Jinkela_splitter_33 (
        .a(G34),
        .b(new_Jinkela_wire_252),
        .c(new_Jinkela_wire_254)
    );

    bfr new_Jinkela_buffer_142 (
        .din(new_Jinkela_wire_203),
        .dout(new_Jinkela_wire_204)
    );

    or_bb _1519_ (
        .a(_0688_),
        .b(new_Jinkela_wire_2432),
        .c(_0689_)
    );

    bfr new_Jinkela_buffer_114 (
        .din(new_Jinkela_wire_135),
        .dout(new_Jinkela_wire_136)
    );

    and_bi _1520_ (
        .a(_0680_),
        .b(new_Jinkela_wire_1647),
        .c(_0690_)
    );

    bfr new_Jinkela_buffer_148 (
        .din(new_Jinkela_wire_214),
        .dout(new_Jinkela_wire_215)
    );

    and_bi _1521_ (
        .a(new_Jinkela_wire_1151),
        .b(_0690_),
        .c(_0691_)
    );

    bfr new_Jinkela_buffer_115 (
        .din(new_Jinkela_wire_136),
        .dout(new_Jinkela_wire_137)
    );

    and_bi _1522_ (
        .a(new_Jinkela_wire_1916),
        .b(_0691_),
        .c(_0692_)
    );

    spl3L new_Jinkela_splitter_26 (
        .a(new_Jinkela_wire_220),
        .d(new_Jinkela_wire_221),
        .b(new_Jinkela_wire_222),
        .c(new_Jinkela_wire_223)
    );

    bfr new_Jinkela_buffer_143 (
        .din(new_Jinkela_wire_204),
        .dout(new_Jinkela_wire_205)
    );

    or_bb _1523_ (
        .a(_0692_),
        .b(new_Jinkela_wire_1348),
        .c(_0693_)
    );

    bfr new_Jinkela_buffer_116 (
        .din(new_Jinkela_wire_137),
        .dout(new_Jinkela_wire_138)
    );

    and_bi _1524_ (
        .a(_0664_),
        .b(new_Jinkela_wire_1567),
        .c(_0694_)
    );

    spl3L new_Jinkela_splitter_28 (
        .a(new_Jinkela_wire_232),
        .d(new_Jinkela_wire_233),
        .b(new_Jinkela_wire_234),
        .c(new_Jinkela_wire_235)
    );

    and_bi _1525_ (
        .a(new_Jinkela_wire_2064),
        .b(new_Jinkela_wire_24),
        .c(_0696_)
    );

    bfr new_Jinkela_buffer_117 (
        .din(new_Jinkela_wire_138),
        .dout(new_Jinkela_wire_139)
    );

    or_bb _1526_ (
        .a(_0696_),
        .b(new_Jinkela_wire_1451),
        .c(_0697_)
    );

    bfr new_Jinkela_buffer_144 (
        .din(new_Jinkela_wire_205),
        .dout(new_Jinkela_wire_206)
    );

    and_bi _1527_ (
        .a(new_Jinkela_wire_2782),
        .b(new_Jinkela_wire_2959),
        .c(_0698_)
    );

    bfr new_Jinkela_buffer_118 (
        .din(new_Jinkela_wire_139),
        .dout(new_Jinkela_wire_140)
    );

    or_bb _1528_ (
        .a(_0698_),
        .b(new_Jinkela_wire_1197),
        .c(new_net_8)
    );

    and_bi _1529_ (
        .a(new_Jinkela_wire_1487),
        .b(new_Jinkela_wire_2066),
        .c(_0699_)
    );

    bfr new_Jinkela_buffer_119 (
        .din(new_Jinkela_wire_140),
        .dout(new_Jinkela_wire_141)
    );

    and_bi _1530_ (
        .a(new_Jinkela_wire_2533),
        .b(new_Jinkela_wire_832),
        .c(_0700_)
    );

    bfr new_Jinkela_buffer_145 (
        .din(new_Jinkela_wire_206),
        .dout(new_Jinkela_wire_207)
    );

    or_bb _1531_ (
        .a(new_Jinkela_wire_1664),
        .b(new_Jinkela_wire_3200),
        .c(_0701_)
    );

    bfr new_Jinkela_buffer_120 (
        .din(new_Jinkela_wire_141),
        .dout(new_Jinkela_wire_142)
    );

    and_bi _1532_ (
        .a(new_Jinkela_wire_242),
        .b(new_Jinkela_wire_1745),
        .c(_0702_)
    );

    and_bi _1533_ (
        .a(new_Jinkela_wire_700),
        .b(new_Jinkela_wire_2351),
        .c(_0703_)
    );

    bfr new_Jinkela_buffer_121 (
        .din(new_Jinkela_wire_142),
        .dout(new_Jinkela_wire_143)
    );

    or_bb _1534_ (
        .a(_0703_),
        .b(new_Jinkela_wire_2885),
        .c(_0704_)
    );

    bfr new_Jinkela_buffer_146 (
        .din(new_Jinkela_wire_207),
        .dout(new_Jinkela_wire_208)
    );

    and_ii _1535_ (
        .a(new_Jinkela_wire_1300),
        .b(new_Jinkela_wire_1128),
        .c(_0706_)
    );

    bfr new_Jinkela_buffer_122 (
        .din(new_Jinkela_wire_143),
        .dout(new_Jinkela_wire_144)
    );

    and_bi _1536_ (
        .a(new_Jinkela_wire_686),
        .b(new_Jinkela_wire_1888),
        .c(_0707_)
    );

    bfr new_Jinkela_buffer_156 (
        .din(new_Jinkela_wire_235),
        .dout(new_Jinkela_wire_236)
    );

    or_bb _1537_ (
        .a(new_Jinkela_wire_1766),
        .b(_0706_),
        .c(_0708_)
    );

    bfr new_Jinkela_buffer_123 (
        .din(new_Jinkela_wire_144),
        .dout(new_Jinkela_wire_145)
    );

    or_bb _1538_ (
        .a(_0708_),
        .b(_0704_),
        .c(_0709_)
    );

    bfr new_Jinkela_buffer_149 (
        .din(new_Jinkela_wire_223),
        .dout(new_Jinkela_wire_224)
    );

    spl2 new_Jinkela_splitter_36 (
        .a(G8),
        .b(new_Jinkela_wire_264),
        .c(new_Jinkela_wire_265)
    );

    and_bi _1539_ (
        .a(new_Jinkela_wire_731),
        .b(new_Jinkela_wire_3009),
        .c(_0710_)
    );

    spl4L new_Jinkela_splitter_34 (
        .a(new_Jinkela_wire_254),
        .d(new_Jinkela_wire_255),
        .e(new_Jinkela_wire_256),
        .b(new_Jinkela_wire_257),
        .c(new_Jinkela_wire_258)
    );

    and_ii _1540_ (
        .a(new_Jinkela_wire_2746),
        .b(new_Jinkela_wire_2418),
        .c(_0711_)
    );

    bfr new_Jinkela_buffer_163 (
        .din(new_Jinkela_wire_252),
        .dout(new_Jinkela_wire_253)
    );

    spl4L new_Jinkela_splitter_187 (
        .a(new_Jinkela_wire_1119),
        .d(new_Jinkela_wire_1120),
        .e(new_Jinkela_wire_1125),
        .b(new_Jinkela_wire_1130),
        .c(new_Jinkela_wire_1135)
    );

    bfr new_Jinkela_buffer_626 (
        .din(new_Jinkela_wire_1104),
        .dout(new_Jinkela_wire_1105)
    );

    bfr new_Jinkela_buffer_635 (
        .din(new_Jinkela_wire_1114),
        .dout(new_Jinkela_wire_1115)
    );

    bfr new_Jinkela_buffer_627 (
        .din(new_Jinkela_wire_1105),
        .dout(new_Jinkela_wire_1106)
    );

    bfr new_Jinkela_buffer_628 (
        .din(new_Jinkela_wire_1106),
        .dout(new_Jinkela_wire_1107)
    );

    spl3L new_Jinkela_splitter_186 (
        .a(new_Jinkela_wire_1115),
        .d(new_Jinkela_wire_1116),
        .b(new_Jinkela_wire_1117),
        .c(new_Jinkela_wire_1118)
    );

    bfr new_Jinkela_buffer_629 (
        .din(new_Jinkela_wire_1107),
        .dout(new_Jinkela_wire_1108)
    );

    spl4L new_Jinkela_splitter_189 (
        .a(new_Jinkela_wire_1125),
        .d(new_Jinkela_wire_1126),
        .e(new_Jinkela_wire_1127),
        .b(new_Jinkela_wire_1128),
        .c(new_Jinkela_wire_1129)
    );

    bfr new_Jinkela_buffer_630 (
        .din(new_Jinkela_wire_1108),
        .dout(new_Jinkela_wire_1109)
    );

    spl4L new_Jinkela_splitter_188 (
        .a(new_Jinkela_wire_1120),
        .d(new_Jinkela_wire_1121),
        .e(new_Jinkela_wire_1122),
        .b(new_Jinkela_wire_1123),
        .c(new_Jinkela_wire_1124)
    );

    bfr new_Jinkela_buffer_631 (
        .din(new_Jinkela_wire_1109),
        .dout(new_Jinkela_wire_1110)
    );

    bfr new_Jinkela_buffer_632 (
        .din(new_Jinkela_wire_1110),
        .dout(new_Jinkela_wire_1111)
    );

    spl3L new_Jinkela_splitter_196 (
        .a(_0236_),
        .d(new_Jinkela_wire_1154),
        .b(new_Jinkela_wire_1155),
        .c(new_Jinkela_wire_1156)
    );

    spl4L new_Jinkela_splitter_190 (
        .a(new_Jinkela_wire_1130),
        .d(new_Jinkela_wire_1131),
        .e(new_Jinkela_wire_1132),
        .b(new_Jinkela_wire_1133),
        .c(new_Jinkela_wire_1134)
    );

    bfr new_Jinkela_buffer_633 (
        .din(new_Jinkela_wire_1111),
        .dout(new_Jinkela_wire_1112)
    );

    spl4L new_Jinkela_splitter_191 (
        .a(new_Jinkela_wire_1135),
        .d(new_Jinkela_wire_1136),
        .e(new_Jinkela_wire_1137),
        .b(new_Jinkela_wire_1138),
        .c(new_Jinkela_wire_1139)
    );

    bfr new_Jinkela_buffer_634 (
        .din(new_Jinkela_wire_1112),
        .dout(new_Jinkela_wire_1113)
    );

    bfr new_Jinkela_buffer_637 (
        .din(new_Jinkela_wire_1149),
        .dout(new_Jinkela_wire_1150)
    );

    bfr new_Jinkela_buffer_639 (
        .din(_0466_),
        .dout(new_Jinkela_wire_1152)
    );

    bfr new_Jinkela_buffer_636 (
        .din(_0679_),
        .dout(new_Jinkela_wire_1149)
    );

    bfr new_Jinkela_buffer_641 (
        .din(_0537_),
        .dout(new_Jinkela_wire_1157)
    );

    bfr new_Jinkela_buffer_638 (
        .din(new_Jinkela_wire_1150),
        .dout(new_Jinkela_wire_1151)
    );

    bfr new_Jinkela_buffer_640 (
        .din(new_Jinkela_wire_1152),
        .dout(new_Jinkela_wire_1153)
    );

    bfr new_Jinkela_buffer_644 (
        .din(_0496_),
        .dout(new_Jinkela_wire_1160)
    );

    bfr new_Jinkela_buffer_642 (
        .din(new_Jinkela_wire_1157),
        .dout(new_Jinkela_wire_1158)
    );

    bfr new_Jinkela_buffer_647 (
        .din(_0159_),
        .dout(new_Jinkela_wire_1163)
    );

    bfr new_Jinkela_buffer_643 (
        .din(new_Jinkela_wire_1158),
        .dout(new_Jinkela_wire_1159)
    );

    bfr new_Jinkela_buffer_645 (
        .din(new_Jinkela_wire_1160),
        .dout(new_Jinkela_wire_1161)
    );

    bfr new_Jinkela_buffer_648 (
        .din(_0391_),
        .dout(new_Jinkela_wire_1164)
    );

    bfr new_Jinkela_buffer_646 (
        .din(new_Jinkela_wire_1161),
        .dout(new_Jinkela_wire_1162)
    );

    spl3L new_Jinkela_splitter_197 (
        .a(_0183_),
        .d(new_Jinkela_wire_1167),
        .b(new_Jinkela_wire_1168),
        .c(new_Jinkela_wire_1169)
    );

    bfr new_Jinkela_buffer_651 (
        .din(_0416_),
        .dout(new_Jinkela_wire_1170)
    );

    bfr new_Jinkela_buffer_649 (
        .din(new_Jinkela_wire_1164),
        .dout(new_Jinkela_wire_1165)
    );

    bfr new_Jinkela_buffer_658 (
        .din(_0131_),
        .dout(new_Jinkela_wire_1179)
    );

    bfr new_Jinkela_buffer_650 (
        .din(new_Jinkela_wire_1165),
        .dout(new_Jinkela_wire_1166)
    );

    bfr new_Jinkela_buffer_652 (
        .din(new_Jinkela_wire_1170),
        .dout(new_Jinkela_wire_1171)
    );

    bfr new_Jinkela_buffer_659 (
        .din(_0003_),
        .dout(new_Jinkela_wire_1180)
    );

    bfr new_Jinkela_buffer_661 (
        .din(_0607_),
        .dout(new_Jinkela_wire_1182)
    );

    bfr new_Jinkela_buffer_653 (
        .din(new_Jinkela_wire_1171),
        .dout(new_Jinkela_wire_1172)
    );

    bfr new_Jinkela_buffer_660 (
        .din(new_Jinkela_wire_1180),
        .dout(new_Jinkela_wire_1181)
    );

    bfr new_Jinkela_buffer_654 (
        .din(new_Jinkela_wire_1172),
        .dout(new_Jinkela_wire_1173)
    );

    bfr new_Jinkela_buffer_1121 (
        .din(new_Jinkela_wire_1836),
        .dout(new_Jinkela_wire_1837)
    );

    bfr new_Jinkela_buffer_1155 (
        .din(new_Jinkela_wire_1899),
        .dout(new_Jinkela_wire_1900)
    );

    bfr new_Jinkela_buffer_1170 (
        .din(_0546_),
        .dout(new_Jinkela_wire_1931)
    );

    bfr new_Jinkela_buffer_1122 (
        .din(new_Jinkela_wire_1837),
        .dout(new_Jinkela_wire_1838)
    );

    bfr new_Jinkela_buffer_1164 (
        .din(new_Jinkela_wire_1920),
        .dout(new_Jinkela_wire_1921)
    );

    bfr new_Jinkela_buffer_1123 (
        .din(new_Jinkela_wire_1838),
        .dout(new_Jinkela_wire_1839)
    );

    bfr new_Jinkela_buffer_1169 (
        .din(new_Jinkela_wire_1927),
        .dout(new_Jinkela_wire_1928)
    );

    bfr new_Jinkela_buffer_1156 (
        .din(new_Jinkela_wire_1900),
        .dout(new_Jinkela_wire_1901)
    );

    bfr new_Jinkela_buffer_1124 (
        .din(new_Jinkela_wire_1839),
        .dout(new_Jinkela_wire_1840)
    );

    bfr new_Jinkela_buffer_1165 (
        .din(new_Jinkela_wire_1921),
        .dout(new_Jinkela_wire_1922)
    );

    bfr new_Jinkela_buffer_1125 (
        .din(new_Jinkela_wire_1840),
        .dout(new_Jinkela_wire_1841)
    );

    bfr new_Jinkela_buffer_1157 (
        .din(new_Jinkela_wire_1901),
        .dout(new_Jinkela_wire_1902)
    );

    bfr new_Jinkela_buffer_1172 (
        .din(_0093_),
        .dout(new_Jinkela_wire_1935)
    );

    bfr new_Jinkela_buffer_1158 (
        .din(new_Jinkela_wire_1902),
        .dout(new_Jinkela_wire_1903)
    );

    bfr new_Jinkela_buffer_1166 (
        .din(new_Jinkela_wire_1922),
        .dout(new_Jinkela_wire_1923)
    );

    bfr new_Jinkela_buffer_1159 (
        .din(new_Jinkela_wire_1903),
        .dout(new_Jinkela_wire_1904)
    );

    spl2 new_Jinkela_splitter_289 (
        .a(new_Jinkela_wire_1904),
        .b(new_Jinkela_wire_1905),
        .c(new_Jinkela_wire_1907)
    );

    spl4L new_Jinkela_splitter_290 (
        .a(new_Jinkela_wire_1907),
        .d(new_Jinkela_wire_1908),
        .e(new_Jinkela_wire_1909),
        .b(new_Jinkela_wire_1910),
        .c(new_Jinkela_wire_1912)
    );

    bfr new_Jinkela_buffer_1160 (
        .din(new_Jinkela_wire_1905),
        .dout(new_Jinkela_wire_1906)
    );

    spl3L new_Jinkela_splitter_300 (
        .a(_0165_),
        .d(new_Jinkela_wire_1980),
        .b(new_Jinkela_wire_1981),
        .c(new_Jinkela_wire_1982)
    );

    spl4L new_Jinkela_splitter_291 (
        .a(new_Jinkela_wire_1912),
        .d(new_Jinkela_wire_1913),
        .e(new_Jinkela_wire_1914),
        .b(new_Jinkela_wire_1915),
        .c(new_Jinkela_wire_1916)
    );

    bfr new_Jinkela_buffer_1161 (
        .din(new_Jinkela_wire_1910),
        .dout(new_Jinkela_wire_1911)
    );

    spl2 new_Jinkela_splitter_294 (
        .a(new_Jinkela_wire_1928),
        .b(new_Jinkela_wire_1929),
        .c(new_Jinkela_wire_1930)
    );

    bfr new_Jinkela_buffer_1171 (
        .din(new_Jinkela_wire_1931),
        .dout(new_Jinkela_wire_1932)
    );

    bfr new_Jinkela_buffer_1179 (
        .din(new_Jinkela_wire_1951),
        .dout(new_Jinkela_wire_1952)
    );

    spl2 new_Jinkela_splitter_295 (
        .a(new_Jinkela_wire_1932),
        .b(new_Jinkela_wire_1933),
        .c(new_Jinkela_wire_1934)
    );

    bfr new_Jinkela_buffer_1207 (
        .din(_0580_),
        .dout(new_Jinkela_wire_1983)
    );

    bfr new_Jinkela_buffer_1208 (
        .din(new_net_1485),
        .dout(new_Jinkela_wire_1984)
    );

    bfr new_Jinkela_buffer_1178 (
        .din(_0771_),
        .dout(new_Jinkela_wire_1951)
    );

    spl3L new_Jinkela_splitter_297 (
        .a(new_Jinkela_wire_1938),
        .d(new_Jinkela_wire_1939),
        .b(new_Jinkela_wire_1940),
        .c(new_Jinkela_wire_1941)
    );

    bfr new_Jinkela_buffer_1180 (
        .din(new_Jinkela_wire_1952),
        .dout(new_Jinkela_wire_1953)
    );

    bfr new_Jinkela_buffer_1173 (
        .din(new_Jinkela_wire_1935),
        .dout(new_Jinkela_wire_1936)
    );

    spl2 new_Jinkela_splitter_296 (
        .a(new_Jinkela_wire_1936),
        .b(new_Jinkela_wire_1937),
        .c(new_Jinkela_wire_1938)
    );

    bfr new_Jinkela_buffer_1174 (
        .din(new_Jinkela_wire_1941),
        .dout(new_Jinkela_wire_1942)
    );

    bfr new_Jinkela_buffer_1181 (
        .din(new_Jinkela_wire_1953),
        .dout(new_Jinkela_wire_1954)
    );

    spl3L new_Jinkela_splitter_298 (
        .a(new_Jinkela_wire_1942),
        .d(new_Jinkela_wire_1943),
        .b(new_Jinkela_wire_1944),
        .c(new_Jinkela_wire_1945)
    );

    bfr new_Jinkela_buffer_1226 (
        .din(_0149_),
        .dout(new_Jinkela_wire_2002)
    );

    spl2 new_Jinkela_splitter_299 (
        .a(new_Jinkela_wire_1945),
        .b(new_Jinkela_wire_1946),
        .c(new_Jinkela_wire_1947)
    );

    bfr new_Jinkela_buffer_1175 (
        .din(new_Jinkela_wire_1947),
        .dout(new_Jinkela_wire_1948)
    );

    bfr new_Jinkela_buffer_1182 (
        .din(new_Jinkela_wire_1954),
        .dout(new_Jinkela_wire_1955)
    );

    bfr new_Jinkela_buffer_1209 (
        .din(new_Jinkela_wire_1984),
        .dout(new_Jinkela_wire_1985)
    );

    bfr new_Jinkela_buffer_1176 (
        .din(new_Jinkela_wire_1948),
        .dout(new_Jinkela_wire_1949)
    );

    bfr new_Jinkela_buffer_1465 (
        .din(new_Jinkela_wire_2376),
        .dout(new_Jinkela_wire_2377)
    );

    and_bi _1163_ (
        .a(new_Jinkela_wire_2512),
        .b(_0333_),
        .c(_0334_)
    );

    inv _1164_ (
        .din(new_Jinkela_wire_534),
        .dout(_0335_)
    );

    spl2 new_Jinkela_splitter_355 (
        .a(_0229_),
        .b(new_Jinkela_wire_2386),
        .c(new_Jinkela_wire_2387)
    );

    bfr new_Jinkela_buffer_1466 (
        .din(new_Jinkela_wire_2377),
        .dout(new_Jinkela_wire_2378)
    );

    and_bi _1165_ (
        .a(new_Jinkela_wire_3230),
        .b(new_Jinkela_wire_2873),
        .c(_0336_)
    );

    inv _1166_ (
        .din(new_Jinkela_wire_2646),
        .dout(_0337_)
    );

    bfr new_Jinkela_buffer_1470 (
        .din(_0280_),
        .dout(new_Jinkela_wire_2384)
    );

    bfr new_Jinkela_buffer_1472 (
        .din(_0029_),
        .dout(new_Jinkela_wire_2388)
    );

    and_bi _1167_ (
        .a(new_Jinkela_wire_2990),
        .b(new_Jinkela_wire_1645),
        .c(_0338_)
    );

    bfr new_Jinkela_buffer_1471 (
        .din(new_Jinkela_wire_2384),
        .dout(new_Jinkela_wire_2385)
    );

    and_ii _1168_ (
        .a(new_Jinkela_wire_2887),
        .b(new_Jinkela_wire_3075),
        .c(_0339_)
    );

    bfr new_Jinkela_buffer_1480 (
        .din(new_Jinkela_wire_2405),
        .dout(new_Jinkela_wire_2406)
    );

    or_bb _1169_ (
        .a(new_Jinkela_wire_899),
        .b(new_Jinkela_wire_3247),
        .c(_0340_)
    );

    and_bi _1170_ (
        .a(new_Jinkela_wire_975),
        .b(new_Jinkela_wire_3079),
        .c(_0341_)
    );

    bfr new_Jinkela_buffer_1473 (
        .din(_0252_),
        .dout(new_Jinkela_wire_2389)
    );

    and_bi _1171_ (
        .a(new_Jinkela_wire_1087),
        .b(_0341_),
        .c(_0342_)
    );

    bfr new_Jinkela_buffer_1479 (
        .din(_0582_),
        .dout(new_Jinkela_wire_2405)
    );

    bfr new_Jinkela_buffer_1481 (
        .din(_0256_),
        .dout(new_Jinkela_wire_2407)
    );

    or_bi _1172_ (
        .a(_0342_),
        .b(new_Jinkela_wire_1488),
        .c(_0343_)
    );

    or_bi _1173_ (
        .a(new_Jinkela_wire_2456),
        .b(new_Jinkela_wire_2451),
        .c(_0344_)
    );

    bfr new_Jinkela_buffer_1482 (
        .din(_0671_),
        .dout(new_Jinkela_wire_2408)
    );

    spl4L new_Jinkela_splitter_361 (
        .a(_0374_),
        .d(new_Jinkela_wire_2411),
        .e(new_Jinkela_wire_2416),
        .b(new_Jinkela_wire_2421),
        .c(new_Jinkela_wire_2426)
    );

    and_bi _1174_ (
        .a(new_Jinkela_wire_2455),
        .b(new_Jinkela_wire_2450),
        .c(_0345_)
    );

    bfr new_Jinkela_buffer_1474 (
        .din(new_Jinkela_wire_2389),
        .dout(new_Jinkela_wire_2390)
    );

    and_bi _1175_ (
        .a(_0344_),
        .b(_0345_),
        .c(_0346_)
    );

    bfr new_Jinkela_buffer_1475 (
        .din(new_Jinkela_wire_2390),
        .dout(new_Jinkela_wire_2391)
    );

    and_bi _1176_ (
        .a(new_Jinkela_wire_2076),
        .b(new_Jinkela_wire_2888),
        .c(_0347_)
    );

    bfr new_Jinkela_buffer_1483 (
        .din(_0522_),
        .dout(new_Jinkela_wire_2409)
    );

    spl2 new_Jinkela_splitter_356 (
        .a(new_Jinkela_wire_2391),
        .b(new_Jinkela_wire_2392),
        .c(new_Jinkela_wire_2393)
    );

    and_ii _1177_ (
        .a(_0347_),
        .b(new_Jinkela_wire_2345),
        .c(_0348_)
    );

    or_bi _1178_ (
        .a(new_Jinkela_wire_2709),
        .b(new_Jinkela_wire_976),
        .c(_0349_)
    );

    spl2 new_Jinkela_splitter_357 (
        .a(new_Jinkela_wire_2393),
        .b(new_Jinkela_wire_2394),
        .c(new_Jinkela_wire_2395)
    );

    and_bi _1179_ (
        .a(new_Jinkela_wire_2025),
        .b(new_Jinkela_wire_1502),
        .c(_0350_)
    );

    and_bb _1180_ (
        .a(new_Jinkela_wire_1143),
        .b(new_Jinkela_wire_1564),
        .c(_0351_)
    );

    bfr new_Jinkela_buffer_1484 (
        .din(new_Jinkela_wire_2409),
        .dout(new_Jinkela_wire_2410)
    );

    bfr new_Jinkela_buffer_1476 (
        .din(new_Jinkela_wire_2395),
        .dout(new_Jinkela_wire_2396)
    );

    and_ii _1181_ (
        .a(_0351_),
        .b(new_Jinkela_wire_2550),
        .c(_0352_)
    );

    and_ii _1182_ (
        .a(_0352_),
        .b(new_Jinkela_wire_2085),
        .c(_0353_)
    );

    bfr new_Jinkela_buffer_1485 (
        .din(_0264_),
        .dout(new_Jinkela_wire_2431)
    );

    spl4L new_Jinkela_splitter_362 (
        .a(new_Jinkela_wire_2411),
        .d(new_Jinkela_wire_2412),
        .e(new_Jinkela_wire_2413),
        .b(new_Jinkela_wire_2414),
        .c(new_Jinkela_wire_2415)
    );

    and_bi _1183_ (
        .a(new_Jinkela_wire_1565),
        .b(new_Jinkela_wire_1142),
        .c(_0354_)
    );

    spl4L new_Jinkela_splitter_363 (
        .a(new_Jinkela_wire_2416),
        .d(new_Jinkela_wire_2417),
        .e(new_Jinkela_wire_2418),
        .b(new_Jinkela_wire_2419),
        .c(new_Jinkela_wire_2420)
    );

    spl2 new_Jinkela_splitter_358 (
        .a(new_Jinkela_wire_2396),
        .b(new_Jinkela_wire_2397),
        .c(new_Jinkela_wire_2398)
    );

    and_bb _1184_ (
        .a(new_Jinkela_wire_919),
        .b(new_Jinkela_wire_2084),
        .c(_0355_)
    );

    spl2 new_Jinkela_splitter_359 (
        .a(new_Jinkela_wire_2398),
        .b(new_Jinkela_wire_2399),
        .c(new_Jinkela_wire_2400)
    );

    or_bi _1185_ (
        .a(new_Jinkela_wire_797),
        .b(new_Jinkela_wire_413),
        .c(_0356_)
    );

    or_bi _1186_ (
        .a(new_Jinkela_wire_2106),
        .b(new_Jinkela_wire_3208),
        .c(_0357_)
    );

    bfr new_Jinkela_buffer_1487 (
        .din(_0618_),
        .dout(new_Jinkela_wire_2433)
    );

    spl2 new_Jinkela_splitter_360 (
        .a(new_Jinkela_wire_2400),
        .b(new_Jinkela_wire_2401),
        .c(new_Jinkela_wire_2402)
    );

    and_bi _1187_ (
        .a(new_Jinkela_wire_147),
        .b(new_Jinkela_wire_488),
        .c(_0358_)
    );

    or_bb _1188_ (
        .a(new_Jinkela_wire_3262),
        .b(new_Jinkela_wire_2508),
        .c(_0359_)
    );

    bfr new_Jinkela_buffer_1486 (
        .din(_0687_),
        .dout(new_Jinkela_wire_2432)
    );

    bfr new_Jinkela_buffer_1477 (
        .din(new_Jinkela_wire_2402),
        .dout(new_Jinkela_wire_2403)
    );

    or_ii _1189_ (
        .a(new_Jinkela_wire_151),
        .b(new_Jinkela_wire_2),
        .c(_0360_)
    );

    and_bb _1190_ (
        .a(new_Jinkela_wire_647),
        .b(new_Jinkela_wire_148),
        .c(_0361_)
    );

    or_bb _1191_ (
        .a(new_Jinkela_wire_2333),
        .b(new_Jinkela_wire_566),
        .c(_0362_)
    );

    bfr new_Jinkela_buffer_1478 (
        .din(new_Jinkela_wire_2403),
        .dout(new_Jinkela_wire_2404)
    );

    and_ii _1192_ (
        .a(new_Jinkela_wire_1358),
        .b(new_Jinkela_wire_2028),
        .c(_0363_)
    );

    spl4L new_Jinkela_splitter_364 (
        .a(new_Jinkela_wire_2421),
        .d(new_Jinkela_wire_2422),
        .e(new_Jinkela_wire_2423),
        .b(new_Jinkela_wire_2424),
        .c(new_Jinkela_wire_2425)
    );

    and_bi _1193_ (
        .a(new_Jinkela_wire_705),
        .b(new_Jinkela_wire_715),
        .c(_0364_)
    );

    spl4L new_Jinkela_splitter_365 (
        .a(new_Jinkela_wire_2426),
        .d(new_Jinkela_wire_2427),
        .e(new_Jinkela_wire_2428),
        .b(new_Jinkela_wire_2429),
        .c(new_Jinkela_wire_2430)
    );

    inv _1194_ (
        .din(_0364_),
        .dout(_0365_)
    );

    bfr new_Jinkela_buffer_1488 (
        .din(_0324_),
        .dout(new_Jinkela_wire_2436)
    );

    and_bi _1195_ (
        .a(new_Jinkela_wire_2926),
        .b(new_Jinkela_wire_1123),
        .c(_0366_)
    );

    spl4L new_Jinkela_splitter_367 (
        .a(_0179_),
        .d(new_Jinkela_wire_2441),
        .e(new_Jinkela_wire_2442),
        .b(new_Jinkela_wire_2443),
        .c(new_Jinkela_wire_2444)
    );

    or_bi _1196_ (
        .a(new_Jinkela_wire_2332),
        .b(new_Jinkela_wire_565),
        .c(_0367_)
    );

    spl2 new_Jinkela_splitter_366 (
        .a(new_Jinkela_wire_2433),
        .b(new_Jinkela_wire_2434),
        .c(new_Jinkela_wire_2435)
    );

    and_bi _1197_ (
        .a(new_Jinkela_wire_2031),
        .b(new_Jinkela_wire_1925),
        .c(_0368_)
    );

    spl2 new_Jinkela_splitter_369 (
        .a(_0343_),
        .b(new_Jinkela_wire_2450),
        .c(new_Jinkela_wire_2451)
    );

    bfr new_Jinkela_buffer_1493 (
        .din(_0373_),
        .dout(new_Jinkela_wire_2445)
    );

    and_bi _1198_ (
        .a(new_Jinkela_wire_2366),
        .b(new_Jinkela_wire_2956),
        .c(_0369_)
    );

    bfr new_Jinkela_buffer_1489 (
        .din(new_Jinkela_wire_2436),
        .dout(new_Jinkela_wire_2437)
    );

    and_bi _1199_ (
        .a(new_Jinkela_wire_2060),
        .b(new_Jinkela_wire_3005),
        .c(_0370_)
    );

    bfr new_Jinkela_buffer_1490 (
        .din(new_Jinkela_wire_2437),
        .dout(new_Jinkela_wire_2438)
    );

    or_bb _1200_ (
        .a(new_Jinkela_wire_1570),
        .b(new_Jinkela_wire_2643),
        .c(_0371_)
    );

    bfr new_Jinkela_buffer_1494 (
        .din(new_Jinkela_wire_2445),
        .dout(new_Jinkela_wire_2446)
    );

    and_bi _1201_ (
        .a(new_Jinkela_wire_2029),
        .b(new_Jinkela_wire_1357),
        .c(_0372_)
    );

    bfr new_Jinkela_buffer_1491 (
        .din(new_Jinkela_wire_2438),
        .dout(new_Jinkela_wire_2439)
    );

    and_bi _1202_ (
        .a(new_Jinkela_wire_2397),
        .b(new_Jinkela_wire_1884),
        .c(_0373_)
    );

    spl3L new_Jinkela_splitter_368 (
        .a(_0150_),
        .d(new_Jinkela_wire_2447),
        .b(new_Jinkela_wire_2448),
        .c(new_Jinkela_wire_2449)
    );

    and_ii _1203_ (
        .a(new_Jinkela_wire_1924),
        .b(new_Jinkela_wire_2030),
        .c(_0374_)
    );

    bfr new_Jinkela_buffer_1492 (
        .din(new_Jinkela_wire_2439),
        .dout(new_Jinkela_wire_2440)
    );

    and_bi _1204_ (
        .a(new_Jinkela_wire_1943),
        .b(new_Jinkela_wire_2424),
        .c(_0375_)
    );

    bfr new_Jinkela_buffer_591 (
        .din(new_Jinkela_wire_1051),
        .dout(new_Jinkela_wire_1052)
    );

    spl2 new_Jinkela_splitter_446 (
        .a(new_Jinkela_wire_3083),
        .b(new_Jinkela_wire_3084),
        .c(new_Jinkela_wire_3085)
    );

    spl4L new_Jinkela_splitter_182 (
        .a(_0309_),
        .d(new_Jinkela_wire_1074),
        .e(new_Jinkela_wire_1075),
        .b(new_Jinkela_wire_1076),
        .c(new_Jinkela_wire_1077)
    );

    spl4L new_Jinkela_splitter_442 (
        .a(new_Jinkela_wire_3062),
        .d(new_Jinkela_wire_3063),
        .e(new_Jinkela_wire_3064),
        .b(new_Jinkela_wire_3065),
        .c(new_Jinkela_wire_3066)
    );

    bfr new_Jinkela_buffer_592 (
        .din(new_Jinkela_wire_1052),
        .dout(new_Jinkela_wire_1053)
    );

    spl3L new_Jinkela_splitter_441 (
        .a(new_Jinkela_wire_3058),
        .d(new_Jinkela_wire_3059),
        .b(new_Jinkela_wire_3060),
        .c(new_Jinkela_wire_3061)
    );

    spl2 new_Jinkela_splitter_183 (
        .a(_0442_),
        .b(new_Jinkela_wire_1088),
        .c(new_Jinkela_wire_1089)
    );

    bfr new_Jinkela_buffer_601 (
        .din(new_Jinkela_wire_1071),
        .dout(new_Jinkela_wire_1072)
    );

    bfr new_Jinkela_buffer_1922 (
        .din(new_Jinkela_wire_3073),
        .dout(new_Jinkela_wire_3074)
    );

    bfr new_Jinkela_buffer_593 (
        .din(new_Jinkela_wire_1053),
        .dout(new_Jinkela_wire_1054)
    );

    spl2 new_Jinkela_splitter_444 (
        .a(new_Jinkela_wire_3074),
        .b(new_Jinkela_wire_3075),
        .c(new_Jinkela_wire_3076)
    );

    bfr new_Jinkela_buffer_603 (
        .din(new_Jinkela_wire_1077),
        .dout(new_Jinkela_wire_1078)
    );

    bfr new_Jinkela_buffer_1931 (
        .din(new_Jinkela_wire_3094),
        .dout(new_Jinkela_wire_3095)
    );

    spl4L new_Jinkela_splitter_179 (
        .a(new_Jinkela_wire_1054),
        .d(new_Jinkela_wire_1055),
        .e(new_Jinkela_wire_1056),
        .b(new_Jinkela_wire_1057),
        .c(new_Jinkela_wire_1058)
    );

    bfr new_Jinkela_buffer_1927 (
        .din(new_Jinkela_wire_3082),
        .dout(new_Jinkela_wire_3083)
    );

    bfr new_Jinkela_buffer_1923 (
        .din(new_Jinkela_wire_3076),
        .dout(new_Jinkela_wire_3077)
    );

    bfr new_Jinkela_buffer_594 (
        .din(new_Jinkela_wire_1058),
        .dout(new_Jinkela_wire_1059)
    );

    bfr new_Jinkela_buffer_1962 (
        .din(_0218_),
        .dout(new_Jinkela_wire_3128)
    );

    bfr new_Jinkela_buffer_602 (
        .din(new_Jinkela_wire_1072),
        .dout(new_Jinkela_wire_1073)
    );

    bfr new_Jinkela_buffer_1924 (
        .din(new_Jinkela_wire_3077),
        .dout(new_Jinkela_wire_3078)
    );

    spl4L new_Jinkela_splitter_180 (
        .a(new_Jinkela_wire_1059),
        .d(new_Jinkela_wire_1060),
        .e(new_Jinkela_wire_1061),
        .b(new_Jinkela_wire_1062),
        .c(new_Jinkela_wire_1063)
    );

    spl2 new_Jinkela_splitter_181 (
        .a(new_Jinkela_wire_1063),
        .b(new_Jinkela_wire_1064),
        .c(new_Jinkela_wire_1065)
    );

    bfr new_Jinkela_buffer_1925 (
        .din(new_Jinkela_wire_3078),
        .dout(new_Jinkela_wire_3079)
    );

    bfr new_Jinkela_buffer_595 (
        .din(new_Jinkela_wire_1065),
        .dout(new_Jinkela_wire_1066)
    );

    bfr new_Jinkela_buffer_1933 (
        .din(new_Jinkela_wire_3096),
        .dout(new_Jinkela_wire_3097)
    );

    bfr new_Jinkela_buffer_1928 (
        .din(new_Jinkela_wire_3085),
        .dout(new_Jinkela_wire_3086)
    );

    bfr new_Jinkela_buffer_613 (
        .din(_0647_),
        .dout(new_Jinkela_wire_1092)
    );

    spl3L new_Jinkela_splitter_447 (
        .a(new_Jinkela_wire_3086),
        .d(new_Jinkela_wire_3087),
        .b(new_Jinkela_wire_3088),
        .c(new_Jinkela_wire_3089)
    );

    bfr new_Jinkela_buffer_604 (
        .din(new_Jinkela_wire_1078),
        .dout(new_Jinkela_wire_1079)
    );

    bfr new_Jinkela_buffer_1935 (
        .din(new_Jinkela_wire_3100),
        .dout(new_Jinkela_wire_3101)
    );

    bfr new_Jinkela_buffer_596 (
        .din(new_Jinkela_wire_1066),
        .dout(new_Jinkela_wire_1067)
    );

    spl2 new_Jinkela_splitter_449 (
        .a(new_Jinkela_wire_3097),
        .b(new_Jinkela_wire_3098),
        .c(new_Jinkela_wire_3099)
    );

    spl3L new_Jinkela_splitter_448 (
        .a(new_Jinkela_wire_3089),
        .d(new_Jinkela_wire_3090),
        .b(new_Jinkela_wire_3091),
        .c(new_Jinkela_wire_3092)
    );

    spl2 new_Jinkela_splitter_184 (
        .a(new_Jinkela_wire_1089),
        .b(new_Jinkela_wire_1090),
        .c(new_Jinkela_wire_1091)
    );

    bfr new_Jinkela_buffer_597 (
        .din(new_Jinkela_wire_1067),
        .dout(new_Jinkela_wire_1068)
    );

    bfr new_Jinkela_buffer_1936 (
        .din(new_Jinkela_wire_3101),
        .dout(new_Jinkela_wire_3102)
    );

    bfr new_Jinkela_buffer_605 (
        .din(new_Jinkela_wire_1079),
        .dout(new_Jinkela_wire_1080)
    );

    bfr new_Jinkela_buffer_1963 (
        .din(_0467_),
        .dout(new_Jinkela_wire_3129)
    );

    bfr new_Jinkela_buffer_620 (
        .din(_0111_),
        .dout(new_Jinkela_wire_1099)
    );

    bfr new_Jinkela_buffer_617 (
        .din(_0301_),
        .dout(new_Jinkela_wire_1096)
    );

    bfr new_Jinkela_buffer_1966 (
        .din(_0144_),
        .dout(new_Jinkela_wire_3132)
    );

    bfr new_Jinkela_buffer_606 (
        .din(new_Jinkela_wire_1080),
        .dout(new_Jinkela_wire_1081)
    );

    bfr new_Jinkela_buffer_1937 (
        .din(new_Jinkela_wire_3102),
        .dout(new_Jinkela_wire_3103)
    );

    bfr new_Jinkela_buffer_614 (
        .din(new_Jinkela_wire_1092),
        .dout(new_Jinkela_wire_1093)
    );

    bfr new_Jinkela_buffer_1964 (
        .din(new_Jinkela_wire_3129),
        .dout(new_Jinkela_wire_3130)
    );

    bfr new_Jinkela_buffer_607 (
        .din(new_Jinkela_wire_1081),
        .dout(new_Jinkela_wire_1082)
    );

    bfr new_Jinkela_buffer_1938 (
        .din(new_Jinkela_wire_3103),
        .dout(new_Jinkela_wire_3104)
    );

    bfr new_Jinkela_buffer_615 (
        .din(new_Jinkela_wire_1093),
        .dout(new_Jinkela_wire_1094)
    );

    bfr new_Jinkela_buffer_1967 (
        .din(_0485_),
        .dout(new_Jinkela_wire_3133)
    );

    bfr new_Jinkela_buffer_608 (
        .din(new_Jinkela_wire_1082),
        .dout(new_Jinkela_wire_1083)
    );

    bfr new_Jinkela_buffer_1939 (
        .din(new_Jinkela_wire_3104),
        .dout(new_Jinkela_wire_3105)
    );

    bfr new_Jinkela_buffer_618 (
        .din(new_Jinkela_wire_1096),
        .dout(new_Jinkela_wire_1097)
    );

    bfr new_Jinkela_buffer_1965 (
        .din(new_Jinkela_wire_3130),
        .dout(new_Jinkela_wire_3131)
    );

    bfr new_Jinkela_buffer_609 (
        .din(new_Jinkela_wire_1083),
        .dout(new_Jinkela_wire_1084)
    );

    bfr new_Jinkela_buffer_1940 (
        .din(new_Jinkela_wire_3105),
        .dout(new_Jinkela_wire_3106)
    );

    bfr new_Jinkela_buffer_616 (
        .din(new_Jinkela_wire_1094),
        .dout(new_Jinkela_wire_1095)
    );

    spl3L new_Jinkela_splitter_450 (
        .a(_0028_),
        .d(new_Jinkela_wire_3134),
        .b(new_Jinkela_wire_3135),
        .c(new_Jinkela_wire_3136)
    );

    bfr new_Jinkela_buffer_610 (
        .din(new_Jinkela_wire_1084),
        .dout(new_Jinkela_wire_1085)
    );

    bfr new_Jinkela_buffer_1969 (
        .din(_0498_),
        .dout(new_Jinkela_wire_3138)
    );

    bfr new_Jinkela_buffer_1941 (
        .din(new_Jinkela_wire_3106),
        .dout(new_Jinkela_wire_3107)
    );

    bfr new_Jinkela_buffer_621 (
        .din(_0661_),
        .dout(new_Jinkela_wire_1100)
    );

    bfr new_Jinkela_buffer_611 (
        .din(new_Jinkela_wire_1085),
        .dout(new_Jinkela_wire_1086)
    );

    spl3L new_Jinkela_splitter_451 (
        .a(new_net_1),
        .d(new_Jinkela_wire_3163),
        .b(new_Jinkela_wire_3164),
        .c(new_Jinkela_wire_3165)
    );

    bfr new_Jinkela_buffer_1942 (
        .din(new_Jinkela_wire_3107),
        .dout(new_Jinkela_wire_3108)
    );

    bfr new_Jinkela_buffer_619 (
        .din(new_Jinkela_wire_1097),
        .dout(new_Jinkela_wire_1098)
    );

    bfr new_Jinkela_buffer_1968 (
        .din(new_Jinkela_wire_3136),
        .dout(new_Jinkela_wire_3137)
    );

    bfr new_Jinkela_buffer_612 (
        .din(new_Jinkela_wire_1086),
        .dout(new_Jinkela_wire_1087)
    );

    spl2 new_Jinkela_splitter_452 (
        .a(_0103_),
        .b(new_Jinkela_wire_3176),
        .c(new_Jinkela_wire_3177)
    );

    bfr new_Jinkela_buffer_1943 (
        .din(new_Jinkela_wire_3108),
        .dout(new_Jinkela_wire_3109)
    );

    spl2 new_Jinkela_splitter_185 (
        .a(_0363_),
        .b(new_Jinkela_wire_1114),
        .c(new_Jinkela_wire_1119)
    );

    spl2 new_Jinkela_splitter_193 (
        .a(_0350_),
        .b(new_Jinkela_wire_1142),
        .c(new_Jinkela_wire_1143)
    );

    bfr new_Jinkela_buffer_622 (
        .din(new_Jinkela_wire_1100),
        .dout(new_Jinkela_wire_1101)
    );

    bfr new_Jinkela_buffer_1944 (
        .din(new_Jinkela_wire_3109),
        .dout(new_Jinkela_wire_3110)
    );

    spl2 new_Jinkela_splitter_192 (
        .a(_0001_),
        .b(new_Jinkela_wire_1140),
        .c(new_Jinkela_wire_1141)
    );

    bfr new_Jinkela_buffer_1970 (
        .din(new_Jinkela_wire_3138),
        .dout(new_Jinkela_wire_3139)
    );

    bfr new_Jinkela_buffer_623 (
        .din(new_Jinkela_wire_1101),
        .dout(new_Jinkela_wire_1102)
    );

    bfr new_Jinkela_buffer_1945 (
        .din(new_Jinkela_wire_3110),
        .dout(new_Jinkela_wire_3111)
    );

    bfr new_Jinkela_buffer_2004 (
        .din(_0320_),
        .dout(new_Jinkela_wire_3178)
    );

    bfr new_Jinkela_buffer_624 (
        .din(new_Jinkela_wire_1102),
        .dout(new_Jinkela_wire_1103)
    );

    bfr new_Jinkela_buffer_1946 (
        .din(new_Jinkela_wire_3111),
        .dout(new_Jinkela_wire_3112)
    );

    spl2 new_Jinkela_splitter_195 (
        .a(_0017_),
        .b(new_Jinkela_wire_1147),
        .c(new_Jinkela_wire_1148)
    );

    bfr new_Jinkela_buffer_1971 (
        .din(new_Jinkela_wire_3139),
        .dout(new_Jinkela_wire_3140)
    );

    spl3L new_Jinkela_splitter_194 (
        .a(_0300_),
        .d(new_Jinkela_wire_1144),
        .b(new_Jinkela_wire_1145),
        .c(new_Jinkela_wire_1146)
    );

    bfr new_Jinkela_buffer_625 (
        .din(new_Jinkela_wire_1103),
        .dout(new_Jinkela_wire_1104)
    );

    bfr new_Jinkela_buffer_1947 (
        .din(new_Jinkela_wire_3112),
        .dout(new_Jinkela_wire_3113)
    );

    spl2 new_Jinkela_splitter_371 (
        .a(_0450_),
        .b(new_Jinkela_wire_2458),
        .c(new_Jinkela_wire_2459)
    );

    bfr new_Jinkela_buffer_1495 (
        .din(_0340_),
        .dout(new_Jinkela_wire_2452)
    );

    bfr new_Jinkela_buffer_1501 (
        .din(new_net_4),
        .dout(new_Jinkela_wire_2462)
    );

    bfr new_Jinkela_buffer_1498 (
        .din(_0081_),
        .dout(new_Jinkela_wire_2457)
    );

    bfr new_Jinkela_buffer_1496 (
        .din(new_Jinkela_wire_2452),
        .dout(new_Jinkela_wire_2453)
    );

    bfr new_Jinkela_buffer_1499 (
        .din(new_Jinkela_wire_2459),
        .dout(new_Jinkela_wire_2460)
    );

    bfr new_Jinkela_buffer_1497 (
        .din(new_Jinkela_wire_2453),
        .dout(new_Jinkela_wire_2454)
    );

    spl2 new_Jinkela_splitter_370 (
        .a(new_Jinkela_wire_2454),
        .b(new_Jinkela_wire_2455),
        .c(new_Jinkela_wire_2456)
    );

    bfr new_Jinkela_buffer_1532 (
        .din(_0315_),
        .dout(new_Jinkela_wire_2496)
    );

    spl4L new_Jinkela_splitter_374 (
        .a(_0792_),
        .d(new_Jinkela_wire_2507),
        .e(new_Jinkela_wire_2508),
        .b(new_Jinkela_wire_2509),
        .c(new_Jinkela_wire_2510)
    );

    bfr new_Jinkela_buffer_1500 (
        .din(new_Jinkela_wire_2460),
        .dout(new_Jinkela_wire_2461)
    );

    bfr new_Jinkela_buffer_1502 (
        .din(new_Jinkela_wire_2462),
        .dout(new_Jinkela_wire_2463)
    );

    bfr new_Jinkela_buffer_1539 (
        .din(_0002_),
        .dout(new_Jinkela_wire_2506)
    );

    bfr new_Jinkela_buffer_1540 (
        .din(new_Jinkela_wire_2510),
        .dout(new_Jinkela_wire_2511)
    );

    bfr new_Jinkela_buffer_1503 (
        .din(new_Jinkela_wire_2463),
        .dout(new_Jinkela_wire_2464)
    );

    bfr new_Jinkela_buffer_1504 (
        .din(new_Jinkela_wire_2464),
        .dout(new_Jinkela_wire_2465)
    );

    bfr new_Jinkela_buffer_1533 (
        .din(new_Jinkela_wire_2496),
        .dout(new_Jinkela_wire_2497)
    );

    bfr new_Jinkela_buffer_1505 (
        .din(new_Jinkela_wire_2465),
        .dout(new_Jinkela_wire_2466)
    );

    bfr new_Jinkela_buffer_1542 (
        .din(_0334_),
        .dout(new_Jinkela_wire_2513)
    );

    spl3L new_Jinkela_splitter_372 (
        .a(new_Jinkela_wire_2466),
        .d(new_Jinkela_wire_2467),
        .b(new_Jinkela_wire_2468),
        .c(new_Jinkela_wire_2469)
    );

    bfr new_Jinkela_buffer_1534 (
        .din(new_Jinkela_wire_2497),
        .dout(new_Jinkela_wire_2498)
    );

    bfr new_Jinkela_buffer_1506 (
        .din(new_Jinkela_wire_2469),
        .dout(new_Jinkela_wire_2470)
    );

    bfr new_Jinkela_buffer_1535 (
        .din(new_Jinkela_wire_2498),
        .dout(new_Jinkela_wire_2499)
    );

    bfr new_Jinkela_buffer_1507 (
        .din(new_Jinkela_wire_2470),
        .dout(new_Jinkela_wire_2471)
    );

    bfr new_Jinkela_buffer_1508 (
        .din(new_Jinkela_wire_2471),
        .dout(new_Jinkela_wire_2472)
    );

    spl3L new_Jinkela_splitter_373 (
        .a(new_Jinkela_wire_2499),
        .d(new_Jinkela_wire_2500),
        .b(new_Jinkela_wire_2501),
        .c(new_Jinkela_wire_2502)
    );

    bfr new_Jinkela_buffer_1509 (
        .din(new_Jinkela_wire_2472),
        .dout(new_Jinkela_wire_2473)
    );

    bfr new_Jinkela_buffer_1510 (
        .din(new_Jinkela_wire_2473),
        .dout(new_Jinkela_wire_2474)
    );

    bfr new_Jinkela_buffer_1536 (
        .din(new_Jinkela_wire_2502),
        .dout(new_Jinkela_wire_2503)
    );

    bfr new_Jinkela_buffer_1511 (
        .din(new_Jinkela_wire_2474),
        .dout(new_Jinkela_wire_2475)
    );

    bfr new_Jinkela_buffer_1541 (
        .din(new_Jinkela_wire_2511),
        .dout(new_Jinkela_wire_2512)
    );

    bfr new_Jinkela_buffer_1512 (
        .din(new_Jinkela_wire_2475),
        .dout(new_Jinkela_wire_2476)
    );

    bfr new_Jinkela_buffer_1537 (
        .din(new_Jinkela_wire_2503),
        .dout(new_Jinkela_wire_2504)
    );

    bfr new_Jinkela_buffer_1513 (
        .din(new_Jinkela_wire_2476),
        .dout(new_Jinkela_wire_2477)
    );

    spl2 new_Jinkela_splitter_380 (
        .a(_0066_),
        .b(new_Jinkela_wire_2551),
        .c(new_Jinkela_wire_2552)
    );

    spl2 new_Jinkela_splitter_386 (
        .a(new_Jinkela_wire_2572),
        .b(new_Jinkela_wire_2573),
        .c(new_Jinkela_wire_2574)
    );

    bfr new_Jinkela_buffer_1514 (
        .din(new_Jinkela_wire_2477),
        .dout(new_Jinkela_wire_2478)
    );

    bfr new_Jinkela_buffer_1538 (
        .din(new_Jinkela_wire_2504),
        .dout(new_Jinkela_wire_2505)
    );

    bfr new_Jinkela_buffer_1515 (
        .din(new_Jinkela_wire_2478),
        .dout(new_Jinkela_wire_2479)
    );

    spl2 new_Jinkela_splitter_385 (
        .a(_0563_),
        .b(new_Jinkela_wire_2571),
        .c(new_Jinkela_wire_2572)
    );

    bfr new_Jinkela_buffer_1577 (
        .din(_0261_),
        .dout(new_Jinkela_wire_2575)
    );

    bfr new_Jinkela_buffer_1516 (
        .din(new_Jinkela_wire_2479),
        .dout(new_Jinkela_wire_2480)
    );

    bfr new_Jinkela_buffer_583 (
        .din(_0730_),
        .dout(new_Jinkela_wire_1025)
    );

    and_bb _0824_ (
        .a(new_Jinkela_wire_2939),
        .b(new_Jinkela_wire_2645),
        .c(_0797_)
    );

    or_bb _1541_ (
        .a(_0711_),
        .b(new_Jinkela_wire_3087),
        .c(_0712_)
    );

    bfr new_Jinkela_buffer_557 (
        .din(new_Jinkela_wire_994),
        .dout(new_Jinkela_wire_995)
    );

    and_bi _0825_ (
        .a(new_Jinkela_wire_3323),
        .b(new_Jinkela_wire_800),
        .c(_0000_)
    );

    or_bb _1542_ (
        .a(new_Jinkela_wire_2823),
        .b(_0710_),
        .c(_0713_)
    );

    bfr new_Jinkela_buffer_570 (
        .din(new_Jinkela_wire_1009),
        .dout(new_Jinkela_wire_1010)
    );

    bfr new_Jinkela_buffer_565 (
        .din(new_Jinkela_wire_1002),
        .dout(new_Jinkela_wire_1003)
    );

    inv _0826_ (
        .din(new_Jinkela_wire_253),
        .dout(_0001_)
    );

    or_bb _1543_ (
        .a(_0713_),
        .b(new_Jinkela_wire_1208),
        .c(_0714_)
    );

    bfr new_Jinkela_buffer_558 (
        .din(new_Jinkela_wire_995),
        .dout(new_Jinkela_wire_996)
    );

    and_ii _0827_ (
        .a(new_Jinkela_wire_509),
        .b(new_Jinkela_wire_477),
        .c(_0002_)
    );

    or_bb _1544_ (
        .a(new_Jinkela_wire_1889),
        .b(new_Jinkela_wire_585),
        .c(_0715_)
    );

    or_bb _0828_ (
        .a(new_Jinkela_wire_2506),
        .b(new_Jinkela_wire_1141),
        .c(_0003_)
    );

    and_bi _1545_ (
        .a(new_Jinkela_wire_406),
        .b(new_Jinkela_wire_2352),
        .c(_0717_)
    );

    bfr new_Jinkela_buffer_559 (
        .din(new_Jinkela_wire_996),
        .dout(new_Jinkela_wire_997)
    );

    and_bi _0829_ (
        .a(new_Jinkela_wire_3229),
        .b(new_Jinkela_wire_1181),
        .c(_0004_)
    );

    and_bi _1546_ (
        .a(new_Jinkela_wire_2035),
        .b(_0717_),
        .c(_0718_)
    );

    bfr new_Jinkela_buffer_566 (
        .din(new_Jinkela_wire_1003),
        .dout(new_Jinkela_wire_1004)
    );

    or_bb _0830_ (
        .a(_0004_),
        .b(new_Jinkela_wire_1792),
        .c(_0005_)
    );

    and_bi _1547_ (
        .a(new_Jinkela_wire_1946),
        .b(new_Jinkela_wire_1116),
        .c(_0719_)
    );

    bfr new_Jinkela_buffer_560 (
        .din(new_Jinkela_wire_997),
        .dout(new_Jinkela_wire_998)
    );

    and_bi _0831_ (
        .a(new_Jinkela_wire_3093),
        .b(_0005_),
        .c(new_net_1481)
    );

    or_bb _1548_ (
        .a(_0719_),
        .b(new_Jinkela_wire_2316),
        .c(_0720_)
    );

    or_bb _0832_ (
        .a(new_Jinkela_wire_779),
        .b(new_Jinkela_wire_511),
        .c(_0006_)
    );

    and_bi _1549_ (
        .a(_0718_),
        .b(_0720_),
        .c(_0721_)
    );

    bfr new_Jinkela_buffer_561 (
        .din(new_Jinkela_wire_998),
        .dout(new_Jinkela_wire_999)
    );

    and_bb _0833_ (
        .a(new_Jinkela_wire_780),
        .b(new_Jinkela_wire_510),
        .c(_0007_)
    );

    or_bb _1550_ (
        .a(new_Jinkela_wire_2214),
        .b(new_Jinkela_wire_2776),
        .c(_0722_)
    );

    bfr new_Jinkela_buffer_571 (
        .din(new_Jinkela_wire_1010),
        .dout(new_Jinkela_wire_1011)
    );

    bfr new_Jinkela_buffer_567 (
        .din(new_Jinkela_wire_1004),
        .dout(new_Jinkela_wire_1005)
    );

    and_bi _0834_ (
        .a(_0006_),
        .b(_0007_),
        .c(_0008_)
    );

    or_bb _1551_ (
        .a(_0722_),
        .b(new_Jinkela_wire_1091),
        .c(_0723_)
    );

    bfr new_Jinkela_buffer_562 (
        .din(new_Jinkela_wire_999),
        .dout(new_Jinkela_wire_1000)
    );

    and_bi _0835_ (
        .a(new_Jinkela_wire_255),
        .b(new_Jinkela_wire_478),
        .c(_0009_)
    );

    or_bb _1552_ (
        .a(new_Jinkela_wire_2754),
        .b(new_Jinkela_wire_2174),
        .c(_0724_)
    );

    and_bi _0836_ (
        .a(new_Jinkela_wire_474),
        .b(new_Jinkela_wire_256),
        .c(_0010_)
    );

    and_bi _1553_ (
        .a(new_Jinkela_wire_1438),
        .b(_0724_),
        .c(_0725_)
    );

    spl2 new_Jinkela_splitter_172 (
        .a(_0207_),
        .b(new_Jinkela_wire_1031),
        .c(new_Jinkela_wire_1032)
    );

    spl2 new_Jinkela_splitter_170 (
        .a(new_Jinkela_wire_1005),
        .b(new_Jinkela_wire_1006),
        .c(new_Jinkela_wire_1007)
    );

    and_ii _0837_ (
        .a(_0010_),
        .b(_0009_),
        .c(_0011_)
    );

    and_bi _1554_ (
        .a(new_Jinkela_wire_965),
        .b(_0725_),
        .c(_0726_)
    );

    bfr new_Jinkela_buffer_568 (
        .din(new_Jinkela_wire_1007),
        .dout(new_Jinkela_wire_1008)
    );

    or_bi _0838_ (
        .a(new_Jinkela_wire_2723),
        .b(new_Jinkela_wire_1515),
        .c(_0012_)
    );

    and_bi _1555_ (
        .a(new_Jinkela_wire_1914),
        .b(_0726_),
        .c(_0728_)
    );

    bfr new_Jinkela_buffer_581 (
        .din(new_Jinkela_wire_1020),
        .dout(new_Jinkela_wire_1021)
    );

    and_bi _0839_ (
        .a(new_Jinkela_wire_2722),
        .b(new_Jinkela_wire_1514),
        .c(_0013_)
    );

    or_bb _1556_ (
        .a(_0728_),
        .b(new_Jinkela_wire_1349),
        .c(_0729_)
    );

    bfr new_Jinkela_buffer_572 (
        .din(new_Jinkela_wire_1011),
        .dout(new_Jinkela_wire_1012)
    );

    and_bi _0840_ (
        .a(_0012_),
        .b(_0013_),
        .c(_0014_)
    );

    and_bi _1557_ (
        .a(_0701_),
        .b(new_Jinkela_wire_2756),
        .c(_0730_)
    );

    bfr new_Jinkela_buffer_589 (
        .din(_0353_),
        .dout(new_Jinkela_wire_1035)
    );

    and_bi _0841_ (
        .a(new_Jinkela_wire_37),
        .b(new_Jinkela_wire_169),
        .c(_0015_)
    );

    or_bb _1558_ (
        .a(new_Jinkela_wire_1030),
        .b(_0700_),
        .c(_0731_)
    );

    bfr new_Jinkela_buffer_573 (
        .din(new_Jinkela_wire_1012),
        .dout(new_Jinkela_wire_1013)
    );

    and_bi _0842_ (
        .a(new_Jinkela_wire_170),
        .b(new_Jinkela_wire_35),
        .c(_0016_)
    );

    or_bb _1559_ (
        .a(new_Jinkela_wire_1351),
        .b(_0699_),
        .c(new_net_7)
    );

    bfr new_Jinkela_buffer_584 (
        .din(new_Jinkela_wire_1025),
        .dout(new_Jinkela_wire_1026)
    );

    bfr new_Jinkela_buffer_582 (
        .din(new_Jinkela_wire_1021),
        .dout(new_Jinkela_wire_1022)
    );

    and_ii _0843_ (
        .a(_0016_),
        .b(_0015_),
        .c(_0017_)
    );

    or_bb _1560_ (
        .a(new_Jinkela_wire_1768),
        .b(new_Jinkela_wire_2797),
        .c(_0732_)
    );

    bfr new_Jinkela_buffer_574 (
        .din(new_Jinkela_wire_1013),
        .dout(new_Jinkela_wire_1014)
    );

    and_bi _0847_ (
        .a(new_Jinkela_wire_1148),
        .b(new_Jinkela_wire_1270),
        .c(_0021_)
    );

    or_bb _1561_ (
        .a(new_Jinkela_wire_948),
        .b(new_Jinkela_wire_1277),
        .c(_0733_)
    );

    and_bi _0848_ (
        .a(new_Jinkela_wire_1269),
        .b(new_Jinkela_wire_1147),
        .c(_0022_)
    );

    or_bb _1562_ (
        .a(new_Jinkela_wire_2113),
        .b(new_Jinkela_wire_1414),
        .c(_0734_)
    );

    bfr new_Jinkela_buffer_575 (
        .din(new_Jinkela_wire_1014),
        .dout(new_Jinkela_wire_1015)
    );

    and_ii _0849_ (
        .a(_0022_),
        .b(_0021_),
        .c(_0023_)
    );

    and_ii _1563_ (
        .a(_0734_),
        .b(new_Jinkela_wire_909),
        .c(_0735_)
    );

    spl2 new_Jinkela_splitter_171 (
        .a(new_Jinkela_wire_1022),
        .b(new_Jinkela_wire_1023),
        .c(new_Jinkela_wire_1024)
    );

    or_bb _0850_ (
        .a(new_Jinkela_wire_1331),
        .b(new_Jinkela_wire_1869),
        .c(_0024_)
    );

    inv _1564_ (
        .din(new_Jinkela_wire_2009),
        .dout(new_net_1479)
    );

    bfr new_Jinkela_buffer_576 (
        .din(new_Jinkela_wire_1015),
        .dout(new_Jinkela_wire_1016)
    );

    and_bb _0851_ (
        .a(new_Jinkela_wire_1330),
        .b(new_Jinkela_wire_1868),
        .c(_0025_)
    );

    and_bi _1565_ (
        .a(new_Jinkela_wire_390),
        .b(new_Jinkela_wire_911),
        .c(_0737_)
    );

    and_bi _0852_ (
        .a(_0024_),
        .b(_0025_),
        .c(new_net_1477)
    );

    or_bi _1566_ (
        .a(new_Jinkela_wire_2008),
        .b(new_Jinkela_wire_145),
        .c(_0738_)
    );

    bfr new_Jinkela_buffer_577 (
        .din(new_Jinkela_wire_1016),
        .dout(new_Jinkela_wire_1017)
    );

    and_bb _0853_ (
        .a(new_Jinkela_wire_194),
        .b(new_Jinkela_wire_268),
        .c(_0026_)
    );

    or_bb _1567_ (
        .a(_0738_),
        .b(new_Jinkela_wire_3234),
        .c(new_net_1473)
    );

    spl2 new_Jinkela_splitter_173 (
        .a(new_Jinkela_wire_1032),
        .b(new_Jinkela_wire_1033),
        .c(new_Jinkela_wire_1034)
    );

    and_ii _0854_ (
        .a(new_Jinkela_wire_2006),
        .b(new_Jinkela_wire_2307),
        .c(_0027_)
    );

    and_bb _1568_ (
        .a(new_Jinkela_wire_2288),
        .b(new_Jinkela_wire_3164),
        .c(_0739_)
    );

    bfr new_Jinkela_buffer_578 (
        .din(new_Jinkela_wire_1017),
        .dout(new_Jinkela_wire_1018)
    );

    or_bb _0855_ (
        .a(new_Jinkela_wire_574),
        .b(new_Jinkela_wire_740),
        .c(_0028_)
    );

    and_bi _1569_ (
        .a(new_Jinkela_wire_910),
        .b(new_Jinkela_wire_3025),
        .c(_0740_)
    );

    bfr new_Jinkela_buffer_585 (
        .din(new_Jinkela_wire_1026),
        .dout(new_Jinkela_wire_1027)
    );

    spl3L new_Jinkela_splitter_174 (
        .a(_0245_),
        .d(new_Jinkela_wire_1036),
        .b(new_Jinkela_wire_1037),
        .c(new_Jinkela_wire_1038)
    );

    and_bb _0856_ (
        .a(new_Jinkela_wire_575),
        .b(new_Jinkela_wire_739),
        .c(_0029_)
    );

    and_bb _1570_ (
        .a(new_Jinkela_wire_2899),
        .b(new_Jinkela_wire_3272),
        .c(_0741_)
    );

    bfr new_Jinkela_buffer_579 (
        .din(new_Jinkela_wire_1018),
        .dout(new_Jinkela_wire_1019)
    );

    and_bi _0857_ (
        .a(new_Jinkela_wire_3134),
        .b(new_Jinkela_wire_2388),
        .c(_0030_)
    );

    or_bi _1571_ (
        .a(new_Jinkela_wire_2273),
        .b(new_Jinkela_wire_1413),
        .c(_0742_)
    );

    bfr new_Jinkela_buffer_586 (
        .din(new_Jinkela_wire_1027),
        .dout(new_Jinkela_wire_1028)
    );

    or_bi _0858_ (
        .a(new_Jinkela_wire_2779),
        .b(new_Jinkela_wire_1353),
        .c(_0031_)
    );

    and_bb _1572_ (
        .a(new_Jinkela_wire_1769),
        .b(new_Jinkela_wire_2798),
        .c(_0743_)
    );

    spl2 new_Jinkela_splitter_175 (
        .a(_0070_),
        .b(new_Jinkela_wire_1039),
        .c(new_Jinkela_wire_1040)
    );

    and_bi _0859_ (
        .a(new_Jinkela_wire_2780),
        .b(new_Jinkela_wire_1352),
        .c(_0032_)
    );

    or_bi _1573_ (
        .a(new_Jinkela_wire_1399),
        .b(new_Jinkela_wire_942),
        .c(_0744_)
    );

    bfr new_Jinkela_buffer_587 (
        .din(new_Jinkela_wire_1028),
        .dout(new_Jinkela_wire_1029)
    );

    and_bi _0860_ (
        .a(_0031_),
        .b(_0032_),
        .c(_0033_)
    );

    and_bb _1574_ (
        .a(new_Jinkela_wire_2657),
        .b(new_Jinkela_wire_1417),
        .c(_0745_)
    );

    bfr new_Jinkela_buffer_598 (
        .din(_0444_),
        .dout(new_Jinkela_wire_1069)
    );

    and_bi _0861_ (
        .a(new_Jinkela_wire_212),
        .b(new_Jinkela_wire_326),
        .c(_0034_)
    );

    and_bi _1575_ (
        .a(new_Jinkela_wire_1276),
        .b(new_Jinkela_wire_1926),
        .c(_0747_)
    );

    bfr new_Jinkela_buffer_588 (
        .din(new_Jinkela_wire_1029),
        .dout(new_Jinkela_wire_1030)
    );

    and_bi _0862_ (
        .a(new_Jinkela_wire_329),
        .b(new_Jinkela_wire_213),
        .c(_0035_)
    );

    and_ii _1576_ (
        .a(new_Jinkela_wire_1497),
        .b(new_Jinkela_wire_1522),
        .c(_0748_)
    );

    and_ii _0863_ (
        .a(_0035_),
        .b(_0034_),
        .c(_0036_)
    );

    and_bb _1577_ (
        .a(new_Jinkela_wire_1496),
        .b(new_Jinkela_wire_1521),
        .c(_0749_)
    );

    and_ii _0864_ (
        .a(new_Jinkela_wire_707),
        .b(new_Jinkela_wire_280),
        .c(_0037_)
    );

    or_bb _1578_ (
        .a(_0749_),
        .b(_0748_),
        .c(_0750_)
    );

    bfr new_Jinkela_buffer_599 (
        .din(new_Jinkela_wire_1069),
        .dout(new_Jinkela_wire_1070)
    );

    and_bb _0865_ (
        .a(new_Jinkela_wire_706),
        .b(new_Jinkela_wire_279),
        .c(_0038_)
    );

    or_bb _1579_ (
        .a(new_Jinkela_wire_2828),
        .b(new_Jinkela_wire_3257),
        .c(_0751_)
    );

    spl2 new_Jinkela_splitter_176 (
        .a(new_Jinkela_wire_1040),
        .b(new_Jinkela_wire_1041),
        .c(new_Jinkela_wire_1046)
    );

    spl4L new_Jinkela_splitter_177 (
        .a(new_Jinkela_wire_1041),
        .d(new_Jinkela_wire_1042),
        .e(new_Jinkela_wire_1043),
        .b(new_Jinkela_wire_1044),
        .c(new_Jinkela_wire_1045)
    );

    and_ii _0866_ (
        .a(_0038_),
        .b(_0037_),
        .c(_0039_)
    );

    and_bb _1580_ (
        .a(new_Jinkela_wire_2827),
        .b(new_Jinkela_wire_3256),
        .c(_0752_)
    );

    and_ii _0867_ (
        .a(new_Jinkela_wire_1674),
        .b(new_Jinkela_wire_1708),
        .c(_0040_)
    );

    and_bi _1581_ (
        .a(_0751_),
        .b(_0752_),
        .c(_0753_)
    );

    spl4L new_Jinkela_splitter_178 (
        .a(new_Jinkela_wire_1046),
        .d(new_Jinkela_wire_1047),
        .e(new_Jinkela_wire_1048),
        .b(new_Jinkela_wire_1049),
        .c(new_Jinkela_wire_1050)
    );

    bfr new_Jinkela_buffer_600 (
        .din(_0540_),
        .dout(new_Jinkela_wire_1071)
    );

    and_bb _0868_ (
        .a(new_Jinkela_wire_1673),
        .b(new_Jinkela_wire_1707),
        .c(_0041_)
    );

    or_bb _1582_ (
        .a(new_Jinkela_wire_1490),
        .b(new_Jinkela_wire_1672),
        .c(_0754_)
    );

    bfr new_Jinkela_buffer_590 (
        .din(_0059_),
        .dout(new_Jinkela_wire_1051)
    );

    bfr new_Jinkela_buffer_1543 (
        .din(new_Jinkela_wire_2513),
        .dout(new_Jinkela_wire_2514)
    );

    bfr new_Jinkela_buffer_1517 (
        .din(new_Jinkela_wire_2480),
        .dout(new_Jinkela_wire_2481)
    );

    bfr new_Jinkela_buffer_1948 (
        .din(new_Jinkela_wire_3113),
        .dout(new_Jinkela_wire_3114)
    );

    bfr new_Jinkela_buffer_1570 (
        .din(new_Jinkela_wire_2552),
        .dout(new_Jinkela_wire_2553)
    );

    bfr new_Jinkela_buffer_1972 (
        .din(new_Jinkela_wire_3140),
        .dout(new_Jinkela_wire_3141)
    );

    bfr new_Jinkela_buffer_1518 (
        .din(new_Jinkela_wire_2481),
        .dout(new_Jinkela_wire_2482)
    );

    bfr new_Jinkela_buffer_1949 (
        .din(new_Jinkela_wire_3114),
        .dout(new_Jinkela_wire_3115)
    );

    bfr new_Jinkela_buffer_1544 (
        .din(new_Jinkela_wire_2514),
        .dout(new_Jinkela_wire_2515)
    );

    bfr new_Jinkela_buffer_1519 (
        .din(new_Jinkela_wire_2482),
        .dout(new_Jinkela_wire_2483)
    );

    bfr new_Jinkela_buffer_1994 (
        .din(new_Jinkela_wire_3165),
        .dout(new_Jinkela_wire_3166)
    );

    bfr new_Jinkela_buffer_1950 (
        .din(new_Jinkela_wire_3115),
        .dout(new_Jinkela_wire_3116)
    );

    bfr new_Jinkela_buffer_1578 (
        .din(_0515_),
        .dout(new_Jinkela_wire_2576)
    );

    bfr new_Jinkela_buffer_1973 (
        .din(new_Jinkela_wire_3141),
        .dout(new_Jinkela_wire_3142)
    );

    bfr new_Jinkela_buffer_1520 (
        .din(new_Jinkela_wire_2483),
        .dout(new_Jinkela_wire_2484)
    );

    bfr new_Jinkela_buffer_1951 (
        .din(new_Jinkela_wire_3116),
        .dout(new_Jinkela_wire_3117)
    );

    bfr new_Jinkela_buffer_1545 (
        .din(new_Jinkela_wire_2515),
        .dout(new_Jinkela_wire_2516)
    );

    bfr new_Jinkela_buffer_2007 (
        .din(_0432_),
        .dout(new_Jinkela_wire_3181)
    );

    bfr new_Jinkela_buffer_1521 (
        .din(new_Jinkela_wire_2484),
        .dout(new_Jinkela_wire_2485)
    );

    bfr new_Jinkela_buffer_1995 (
        .din(new_Jinkela_wire_3166),
        .dout(new_Jinkela_wire_3167)
    );

    bfr new_Jinkela_buffer_1952 (
        .din(new_Jinkela_wire_3117),
        .dout(new_Jinkela_wire_3118)
    );

    bfr new_Jinkela_buffer_1579 (
        .din(new_Jinkela_wire_2576),
        .dout(new_Jinkela_wire_2577)
    );

    bfr new_Jinkela_buffer_1974 (
        .din(new_Jinkela_wire_3142),
        .dout(new_Jinkela_wire_3143)
    );

    bfr new_Jinkela_buffer_1522 (
        .din(new_Jinkela_wire_2485),
        .dout(new_Jinkela_wire_2486)
    );

    bfr new_Jinkela_buffer_1953 (
        .din(new_Jinkela_wire_3118),
        .dout(new_Jinkela_wire_3119)
    );

    bfr new_Jinkela_buffer_1546 (
        .din(new_Jinkela_wire_2516),
        .dout(new_Jinkela_wire_2517)
    );

    bfr new_Jinkela_buffer_1523 (
        .din(new_Jinkela_wire_2486),
        .dout(new_Jinkela_wire_2487)
    );

    bfr new_Jinkela_buffer_1954 (
        .din(new_Jinkela_wire_3119),
        .dout(new_Jinkela_wire_3120)
    );

    bfr new_Jinkela_buffer_1572 (
        .din(new_Jinkela_wire_2554),
        .dout(new_Jinkela_wire_2555)
    );

    bfr new_Jinkela_buffer_1975 (
        .din(new_Jinkela_wire_3143),
        .dout(new_Jinkela_wire_3144)
    );

    bfr new_Jinkela_buffer_1524 (
        .din(new_Jinkela_wire_2487),
        .dout(new_Jinkela_wire_2488)
    );

    bfr new_Jinkela_buffer_1955 (
        .din(new_Jinkela_wire_3120),
        .dout(new_Jinkela_wire_3121)
    );

    bfr new_Jinkela_buffer_2005 (
        .din(_0519_),
        .dout(new_Jinkela_wire_3179)
    );

    bfr new_Jinkela_buffer_1525 (
        .din(new_Jinkela_wire_2488),
        .dout(new_Jinkela_wire_2489)
    );

    bfr new_Jinkela_buffer_1996 (
        .din(new_Jinkela_wire_3167),
        .dout(new_Jinkela_wire_3168)
    );

    bfr new_Jinkela_buffer_1956 (
        .din(new_Jinkela_wire_3121),
        .dout(new_Jinkela_wire_3122)
    );

    bfr new_Jinkela_buffer_1548 (
        .din(new_Jinkela_wire_2518),
        .dout(new_Jinkela_wire_2519)
    );

    bfr new_Jinkela_buffer_1976 (
        .din(new_Jinkela_wire_3144),
        .dout(new_Jinkela_wire_3145)
    );

    bfr new_Jinkela_buffer_1526 (
        .din(new_Jinkela_wire_2489),
        .dout(new_Jinkela_wire_2490)
    );

    bfr new_Jinkela_buffer_1957 (
        .din(new_Jinkela_wire_3122),
        .dout(new_Jinkela_wire_3123)
    );

    bfr new_Jinkela_buffer_1547 (
        .din(new_Jinkela_wire_2517),
        .dout(new_Jinkela_wire_2518)
    );

    bfr new_Jinkela_buffer_1527 (
        .din(new_Jinkela_wire_2490),
        .dout(new_Jinkela_wire_2491)
    );

    bfr new_Jinkela_buffer_2012 (
        .din(_0596_),
        .dout(new_Jinkela_wire_3188)
    );

    bfr new_Jinkela_buffer_1958 (
        .din(new_Jinkela_wire_3123),
        .dout(new_Jinkela_wire_3124)
    );

    bfr new_Jinkela_buffer_1977 (
        .din(new_Jinkela_wire_3145),
        .dout(new_Jinkela_wire_3146)
    );

    bfr new_Jinkela_buffer_1528 (
        .din(new_Jinkela_wire_2491),
        .dout(new_Jinkela_wire_2492)
    );

    bfr new_Jinkela_buffer_1959 (
        .din(new_Jinkela_wire_3124),
        .dout(new_Jinkela_wire_3125)
    );

    bfr new_Jinkela_buffer_1571 (
        .din(new_Jinkela_wire_2553),
        .dout(new_Jinkela_wire_2554)
    );

    bfr new_Jinkela_buffer_2006 (
        .din(new_Jinkela_wire_3179),
        .dout(new_Jinkela_wire_3180)
    );

    bfr new_Jinkela_buffer_1529 (
        .din(new_Jinkela_wire_2492),
        .dout(new_Jinkela_wire_2493)
    );

    bfr new_Jinkela_buffer_1997 (
        .din(new_Jinkela_wire_3168),
        .dout(new_Jinkela_wire_3169)
    );

    bfr new_Jinkela_buffer_1960 (
        .din(new_Jinkela_wire_3125),
        .dout(new_Jinkela_wire_3126)
    );

    bfr new_Jinkela_buffer_1550 (
        .din(new_Jinkela_wire_2520),
        .dout(new_Jinkela_wire_2521)
    );

    bfr new_Jinkela_buffer_1581 (
        .din(new_Jinkela_wire_2580),
        .dout(new_Jinkela_wire_2581)
    );

    bfr new_Jinkela_buffer_1978 (
        .din(new_Jinkela_wire_3146),
        .dout(new_Jinkela_wire_3147)
    );

    bfr new_Jinkela_buffer_1530 (
        .din(new_Jinkela_wire_2493),
        .dout(new_Jinkela_wire_2494)
    );

    bfr new_Jinkela_buffer_1961 (
        .din(new_Jinkela_wire_3126),
        .dout(new_Jinkela_wire_3127)
    );

    bfr new_Jinkela_buffer_1549 (
        .din(new_Jinkela_wire_2519),
        .dout(new_Jinkela_wire_2520)
    );

    bfr new_Jinkela_buffer_1531 (
        .din(new_Jinkela_wire_2494),
        .dout(new_Jinkela_wire_2495)
    );

    bfr new_Jinkela_buffer_1979 (
        .din(new_Jinkela_wire_3147),
        .dout(new_Jinkela_wire_3148)
    );

    bfr new_Jinkela_buffer_1580 (
        .din(_0594_),
        .dout(new_Jinkela_wire_2580)
    );

    bfr new_Jinkela_buffer_1573 (
        .din(new_Jinkela_wire_2555),
        .dout(new_Jinkela_wire_2556)
    );

    bfr new_Jinkela_buffer_2008 (
        .din(new_Jinkela_wire_3181),
        .dout(new_Jinkela_wire_3182)
    );

    bfr new_Jinkela_buffer_1998 (
        .din(new_Jinkela_wire_3169),
        .dout(new_Jinkela_wire_3170)
    );

    spl2 new_Jinkela_splitter_387 (
        .a(_0375_),
        .b(new_Jinkela_wire_2578),
        .c(new_Jinkela_wire_2579)
    );

    bfr new_Jinkela_buffer_1980 (
        .din(new_Jinkela_wire_3148),
        .dout(new_Jinkela_wire_3149)
    );

    bfr new_Jinkela_buffer_1552 (
        .din(new_Jinkela_wire_2522),
        .dout(new_Jinkela_wire_2523)
    );

    bfr new_Jinkela_buffer_1551 (
        .din(new_Jinkela_wire_2521),
        .dout(new_Jinkela_wire_2522)
    );

    bfr new_Jinkela_buffer_1981 (
        .din(new_Jinkela_wire_3149),
        .dout(new_Jinkela_wire_3150)
    );

    bfr new_Jinkela_buffer_1574 (
        .din(new_Jinkela_wire_2556),
        .dout(new_Jinkela_wire_2557)
    );

    spl4L new_Jinkela_splitter_454 (
        .a(_0117_),
        .d(new_Jinkela_wire_3190),
        .e(new_Jinkela_wire_3191),
        .b(new_Jinkela_wire_3192),
        .c(new_Jinkela_wire_3193)
    );

    bfr new_Jinkela_buffer_1553 (
        .din(new_Jinkela_wire_2523),
        .dout(new_Jinkela_wire_2524)
    );

    bfr new_Jinkela_buffer_1999 (
        .din(new_Jinkela_wire_3170),
        .dout(new_Jinkela_wire_3171)
    );

    bfr new_Jinkela_buffer_1982 (
        .din(new_Jinkela_wire_3150),
        .dout(new_Jinkela_wire_3151)
    );

    bfr new_Jinkela_buffer_1583 (
        .din(_0577_),
        .dout(new_Jinkela_wire_2583)
    );

    bfr new_Jinkela_buffer_1554 (
        .din(new_Jinkela_wire_2524),
        .dout(new_Jinkela_wire_2525)
    );

    bfr new_Jinkela_buffer_1983 (
        .din(new_Jinkela_wire_3151),
        .dout(new_Jinkela_wire_3152)
    );

    bfr new_Jinkela_buffer_1575 (
        .din(new_Jinkela_wire_2557),
        .dout(new_Jinkela_wire_2558)
    );

    bfr new_Jinkela_buffer_1555 (
        .din(new_Jinkela_wire_2525),
        .dout(new_Jinkela_wire_2526)
    );

    bfr new_Jinkela_buffer_2000 (
        .din(new_Jinkela_wire_3171),
        .dout(new_Jinkela_wire_3172)
    );

    bfr new_Jinkela_buffer_1984 (
        .din(new_Jinkela_wire_3152),
        .dout(new_Jinkela_wire_3153)
    );

    spl4L new_Jinkela_splitter_388 (
        .a(_0223_),
        .d(new_Jinkela_wire_2584),
        .e(new_Jinkela_wire_2585),
        .b(new_Jinkela_wire_2586),
        .c(new_Jinkela_wire_2587)
    );

    bfr new_Jinkela_buffer_1556 (
        .din(new_Jinkela_wire_2526),
        .dout(new_Jinkela_wire_2527)
    );

    bfr new_Jinkela_buffer_2015 (
        .din(_0310_),
        .dout(new_Jinkela_wire_3195)
    );

    bfr new_Jinkela_buffer_1985 (
        .din(new_Jinkela_wire_3153),
        .dout(new_Jinkela_wire_3154)
    );

    bfr new_Jinkela_buffer_150 (
        .din(new_Jinkela_wire_224),
        .dout(new_Jinkela_wire_225)
    );

    bfr new_Jinkela_buffer_164 (
        .din(new_Jinkela_wire_260),
        .dout(new_Jinkela_wire_261)
    );

    bfr new_Jinkela_buffer_151 (
        .din(new_Jinkela_wire_225),
        .dout(new_Jinkela_wire_226)
    );

    spl2 new_Jinkela_splitter_41 (
        .a(G18),
        .b(new_Jinkela_wire_290),
        .c(new_Jinkela_wire_291)
    );

    bfr new_Jinkela_buffer_152 (
        .din(new_Jinkela_wire_226),
        .dout(new_Jinkela_wire_227)
    );

    bfr new_Jinkela_buffer_157 (
        .din(new_Jinkela_wire_239),
        .dout(new_Jinkela_wire_240)
    );

    bfr new_Jinkela_buffer_153 (
        .din(new_Jinkela_wire_227),
        .dout(new_Jinkela_wire_228)
    );

    spl3L new_Jinkela_splitter_29 (
        .a(new_Jinkela_wire_236),
        .d(new_Jinkela_wire_237),
        .b(new_Jinkela_wire_238),
        .c(new_Jinkela_wire_239)
    );

    spl2 new_Jinkela_splitter_35 (
        .a(new_Jinkela_wire_258),
        .b(new_Jinkela_wire_259),
        .c(new_Jinkela_wire_260)
    );

    spl2 new_Jinkela_splitter_27 (
        .a(new_Jinkela_wire_228),
        .b(new_Jinkela_wire_229),
        .c(new_Jinkela_wire_230)
    );

    bfr new_Jinkela_buffer_154 (
        .din(new_Jinkela_wire_230),
        .dout(new_Jinkela_wire_231)
    );

    bfr new_Jinkela_buffer_158 (
        .din(new_Jinkela_wire_240),
        .dout(new_Jinkela_wire_241)
    );

    bfr new_Jinkela_buffer_171 (
        .din(G46),
        .dout(new_Jinkela_wire_274)
    );

    spl2 new_Jinkela_splitter_30 (
        .a(new_Jinkela_wire_241),
        .b(new_Jinkela_wire_242),
        .c(new_Jinkela_wire_243)
    );

    bfr new_Jinkela_buffer_159 (
        .din(new_Jinkela_wire_243),
        .dout(new_Jinkela_wire_244)
    );

    spl4L new_Jinkela_splitter_38 (
        .a(G14),
        .d(new_Jinkela_wire_275),
        .e(new_Jinkela_wire_276),
        .b(new_Jinkela_wire_277),
        .c(new_Jinkela_wire_278)
    );

    bfr new_Jinkela_buffer_184 (
        .din(G32),
        .dout(new_Jinkela_wire_302)
    );

    bfr new_Jinkela_buffer_167 (
        .din(new_Jinkela_wire_269),
        .dout(new_Jinkela_wire_270)
    );

    bfr new_Jinkela_buffer_168 (
        .din(new_Jinkela_wire_270),
        .dout(new_Jinkela_wire_271)
    );

    spl2 new_Jinkela_splitter_31 (
        .a(new_Jinkela_wire_244),
        .b(new_Jinkela_wire_245),
        .c(new_Jinkela_wire_246)
    );

    spl2 new_Jinkela_splitter_32 (
        .a(new_Jinkela_wire_246),
        .b(new_Jinkela_wire_247),
        .c(new_Jinkela_wire_248)
    );

    bfr new_Jinkela_buffer_165 (
        .din(new_Jinkela_wire_261),
        .dout(new_Jinkela_wire_262)
    );

    bfr new_Jinkela_buffer_160 (
        .din(new_Jinkela_wire_248),
        .dout(new_Jinkela_wire_249)
    );

    bfr new_Jinkela_buffer_176 (
        .din(new_Jinkela_wire_291),
        .dout(new_Jinkela_wire_292)
    );

    bfr new_Jinkela_buffer_166 (
        .din(new_Jinkela_wire_262),
        .dout(new_Jinkela_wire_263)
    );

    bfr new_Jinkela_buffer_161 (
        .din(new_Jinkela_wire_249),
        .dout(new_Jinkela_wire_250)
    );

    bfr new_Jinkela_buffer_162 (
        .din(new_Jinkela_wire_250),
        .dout(new_Jinkela_wire_251)
    );

    spl3L new_Jinkela_splitter_40 (
        .a(new_Jinkela_wire_282),
        .d(new_Jinkela_wire_283),
        .b(new_Jinkela_wire_284),
        .c(new_Jinkela_wire_285)
    );

    spl4L new_Jinkela_splitter_39 (
        .a(new_Jinkela_wire_278),
        .d(new_Jinkela_wire_279),
        .e(new_Jinkela_wire_280),
        .b(new_Jinkela_wire_281),
        .c(new_Jinkela_wire_282)
    );

    bfr new_Jinkela_buffer_169 (
        .din(new_Jinkela_wire_271),
        .dout(new_Jinkela_wire_272)
    );

    bfr new_Jinkela_buffer_170 (
        .din(new_Jinkela_wire_272),
        .dout(new_Jinkela_wire_273)
    );

    bfr new_Jinkela_buffer_172 (
        .din(new_Jinkela_wire_285),
        .dout(new_Jinkela_wire_286)
    );

    spl3L new_Jinkela_splitter_45 (
        .a(G42),
        .d(new_Jinkela_wire_310),
        .b(new_Jinkela_wire_311),
        .c(new_Jinkela_wire_312)
    );

    bfr new_Jinkela_buffer_177 (
        .din(new_Jinkela_wire_292),
        .dout(new_Jinkela_wire_293)
    );

    bfr new_Jinkela_buffer_173 (
        .din(new_Jinkela_wire_286),
        .dout(new_Jinkela_wire_287)
    );

    spl4L new_Jinkela_splitter_43 (
        .a(new_Jinkela_wire_302),
        .d(new_Jinkela_wire_303),
        .e(new_Jinkela_wire_304),
        .b(new_Jinkela_wire_305),
        .c(new_Jinkela_wire_306)
    );

    bfr new_Jinkela_buffer_174 (
        .din(new_Jinkela_wire_287),
        .dout(new_Jinkela_wire_288)
    );

    spl3L new_Jinkela_splitter_47 (
        .a(G11),
        .d(new_Jinkela_wire_323),
        .b(new_Jinkela_wire_324),
        .c(new_Jinkela_wire_327)
    );

    bfr new_Jinkela_buffer_178 (
        .din(new_Jinkela_wire_293),
        .dout(new_Jinkela_wire_294)
    );

    bfr new_Jinkela_buffer_175 (
        .din(new_Jinkela_wire_288),
        .dout(new_Jinkela_wire_289)
    );

    spl2 new_Jinkela_splitter_44 (
        .a(new_Jinkela_wire_306),
        .b(new_Jinkela_wire_307),
        .c(new_Jinkela_wire_308)
    );

    bfr new_Jinkela_buffer_179 (
        .din(new_Jinkela_wire_294),
        .dout(new_Jinkela_wire_295)
    );

    and_ii _1205_ (
        .a(new_Jinkela_wire_2551),
        .b(new_Jinkela_wire_649),
        .c(_0376_)
    );

    or_bb _1206_ (
        .a(_0376_),
        .b(new_Jinkela_wire_2946),
        .c(_0377_)
    );

    and_bi _1207_ (
        .a(new_Jinkela_wire_2760),
        .b(new_Jinkela_wire_1746),
        .c(_0378_)
    );

    or_bb _1208_ (
        .a(new_Jinkela_wire_1243),
        .b(new_Jinkela_wire_2579),
        .c(_0379_)
    );

    or_bb _1209_ (
        .a(_0379_),
        .b(new_Jinkela_wire_2446),
        .c(_0380_)
    );

    and_bi _1210_ (
        .a(new_Jinkela_wire_247),
        .b(new_Jinkela_wire_2353),
        .c(_0381_)
    );

    inv _1211_ (
        .din(new_Jinkela_wire_419),
        .dout(_0382_)
    );

    inv _1212_ (
        .din(new_Jinkela_wire_210),
        .dout(_0383_)
    );

    and_bi _1213_ (
        .a(new_Jinkela_wire_926),
        .b(new_Jinkela_wire_2428),
        .c(_0384_)
    );

    or_bb _1214_ (
        .a(new_Jinkela_wire_1918),
        .b(new_Jinkela_wire_3091),
        .c(_0385_)
    );

    or_bb _1215_ (
        .a(_0385_),
        .b(new_Jinkela_wire_2383),
        .c(_0386_)
    );

    or_bb _1216_ (
        .a(_0386_),
        .b(_0380_),
        .c(_0387_)
    );

    or_bb _1217_ (
        .a(new_Jinkela_wire_3046),
        .b(_0371_),
        .c(_0388_)
    );

    or_bi _1218_ (
        .a(new_Jinkela_wire_1127),
        .b(new_Jinkela_wire_765),
        .c(_0389_)
    );

    and_bi _1219_ (
        .a(new_Jinkela_wire_471),
        .b(new_Jinkela_wire_2357),
        .c(_0390_)
    );

    and_bi _1220_ (
        .a(new_Jinkela_wire_400),
        .b(new_Jinkela_wire_1738),
        .c(_0391_)
    );

    or_bb _1221_ (
        .a(new_Jinkela_wire_1166),
        .b(_0390_),
        .c(_0392_)
    );

    and_bi _1222_ (
        .a(new_Jinkela_wire_2637),
        .b(_0392_),
        .c(_0393_)
    );

    and_bi _1223_ (
        .a(new_Jinkela_wire_672),
        .b(new_Jinkela_wire_1118),
        .c(_0394_)
    );

    or_bb _1224_ (
        .a(_0394_),
        .b(new_Jinkela_wire_455),
        .c(_0395_)
    );

    and_bi _1225_ (
        .a(new_Jinkela_wire_507),
        .b(new_Jinkela_wire_2998),
        .c(_0396_)
    );

    and_bi _1226_ (
        .a(new_Jinkela_wire_299),
        .b(new_Jinkela_wire_1882),
        .c(_0397_)
    );

    and_bi _1227_ (
        .a(new_Jinkela_wire_568),
        .b(new_Jinkela_wire_180),
        .c(_0398_)
    );

    and_ii _1228_ (
        .a(new_Jinkela_wire_1188),
        .b(new_Jinkela_wire_2425),
        .c(_0399_)
    );

    or_bb _1229_ (
        .a(_0399_),
        .b(_0397_),
        .c(_0400_)
    );

    or_bb _1230_ (
        .a(new_Jinkela_wire_968),
        .b(_0396_),
        .c(_0401_)
    );

    or_bb _1231_ (
        .a(_0401_),
        .b(new_Jinkela_wire_845),
        .c(_0402_)
    );

    and_bi _1232_ (
        .a(new_Jinkela_wire_2786),
        .b(_0402_),
        .c(_0403_)
    );

    and_bi _1233_ (
        .a(_0388_),
        .b(_0403_),
        .c(_0404_)
    );

    and_bi _1234_ (
        .a(new_Jinkela_wire_1911),
        .b(_0404_),
        .c(_0405_)
    );

    and_bi _1235_ (
        .a(new_Jinkela_wire_2648),
        .b(new_Jinkela_wire_644),
        .c(_0406_)
    );

    inv _1236_ (
        .din(new_Jinkela_wire_1439),
        .dout(_0407_)
    );

    or_bb _1237_ (
        .a(new_Jinkela_wire_1344),
        .b(_0405_),
        .c(_0408_)
    );

    and_bi _1238_ (
        .a(_0357_),
        .b(new_Jinkela_wire_2380),
        .c(_0409_)
    );

    or_bb _1239_ (
        .a(new_Jinkela_wire_1262),
        .b(_0355_),
        .c(_0410_)
    );

    or_bb _1240_ (
        .a(_0410_),
        .b(new_Jinkela_wire_1035),
        .c(new_net_1)
    );

    and_bi _1241_ (
        .a(new_Jinkela_wire_2086),
        .b(new_Jinkela_wire_2501),
        .c(_0411_)
    );

    or_bb _1242_ (
        .a(new_Jinkela_wire_1024),
        .b(new_Jinkela_wire_2034),
        .c(_0412_)
    );

    or_ii _1243_ (
        .a(new_Jinkela_wire_1023),
        .b(new_Jinkela_wire_2033),
        .c(_0413_)
    );

    or_ii _1244_ (
        .a(_0413_),
        .b(_0412_),
        .c(_0414_)
    );

    or_bb _1245_ (
        .a(new_Jinkela_wire_2927),
        .b(new_Jinkela_wire_2107),
        .c(_0415_)
    );

    and_ii _1246_ (
        .a(new_Jinkela_wire_391),
        .b(new_Jinkela_wire_290),
        .c(_0416_)
    );

    bfr new_Jinkela_buffer_524 (
        .din(new_Jinkela_wire_945),
        .dout(new_Jinkela_wire_946)
    );

    bfr new_Jinkela_buffer_495 (
        .din(new_Jinkela_wire_888),
        .dout(new_Jinkela_wire_889)
    );

    bfr new_Jinkela_buffer_2013 (
        .din(new_Jinkela_wire_3188),
        .dout(new_Jinkela_wire_3189)
    );

    bfr new_Jinkela_buffer_2001 (
        .din(new_Jinkela_wire_3172),
        .dout(new_Jinkela_wire_3173)
    );

    bfr new_Jinkela_buffer_1986 (
        .din(new_Jinkela_wire_3154),
        .dout(new_Jinkela_wire_3155)
    );

    bfr new_Jinkela_buffer_530 (
        .din(new_Jinkela_wire_954),
        .dout(new_Jinkela_wire_955)
    );

    bfr new_Jinkela_buffer_496 (
        .din(new_Jinkela_wire_889),
        .dout(new_Jinkela_wire_890)
    );

    spl2 new_Jinkela_splitter_453 (
        .a(new_Jinkela_wire_3182),
        .b(new_Jinkela_wire_3183),
        .c(new_Jinkela_wire_3184)
    );

    bfr new_Jinkela_buffer_529 (
        .din(new_Jinkela_wire_950),
        .dout(new_Jinkela_wire_951)
    );

    bfr new_Jinkela_buffer_1987 (
        .din(new_Jinkela_wire_3155),
        .dout(new_Jinkela_wire_3156)
    );

    bfr new_Jinkela_buffer_525 (
        .din(new_Jinkela_wire_946),
        .dout(new_Jinkela_wire_947)
    );

    bfr new_Jinkela_buffer_497 (
        .din(new_Jinkela_wire_890),
        .dout(new_Jinkela_wire_891)
    );

    bfr new_Jinkela_buffer_2002 (
        .din(new_Jinkela_wire_3173),
        .dout(new_Jinkela_wire_3174)
    );

    bfr new_Jinkela_buffer_1988 (
        .din(new_Jinkela_wire_3156),
        .dout(new_Jinkela_wire_3157)
    );

    spl3L new_Jinkela_splitter_166 (
        .a(_0214_),
        .d(new_Jinkela_wire_962),
        .b(new_Jinkela_wire_963),
        .c(new_Jinkela_wire_964)
    );

    bfr new_Jinkela_buffer_526 (
        .din(new_Jinkela_wire_947),
        .dout(new_Jinkela_wire_948)
    );

    bfr new_Jinkela_buffer_2009 (
        .din(new_Jinkela_wire_3184),
        .dout(new_Jinkela_wire_3185)
    );

    bfr new_Jinkela_buffer_1989 (
        .din(new_Jinkela_wire_3157),
        .dout(new_Jinkela_wire_3158)
    );

    bfr new_Jinkela_buffer_2003 (
        .din(new_Jinkela_wire_3174),
        .dout(new_Jinkela_wire_3175)
    );

    bfr new_Jinkela_buffer_535 (
        .din(_0714_),
        .dout(new_Jinkela_wire_965)
    );

    bfr new_Jinkela_buffer_1990 (
        .din(new_Jinkela_wire_3158),
        .dout(new_Jinkela_wire_3159)
    );

    bfr new_Jinkela_buffer_531 (
        .din(new_Jinkela_wire_955),
        .dout(new_Jinkela_wire_956)
    );

    bfr new_Jinkela_buffer_536 (
        .din(_0400_),
        .dout(new_Jinkela_wire_966)
    );

    bfr new_Jinkela_buffer_1991 (
        .din(new_Jinkela_wire_3159),
        .dout(new_Jinkela_wire_3160)
    );

    bfr new_Jinkela_buffer_532 (
        .din(new_Jinkela_wire_956),
        .dout(new_Jinkela_wire_957)
    );

    bfr new_Jinkela_buffer_2014 (
        .din(new_Jinkela_wire_3193),
        .dout(new_Jinkela_wire_3194)
    );

    bfr new_Jinkela_buffer_539 (
        .din(_0508_),
        .dout(new_Jinkela_wire_969)
    );

    bfr new_Jinkela_buffer_1992 (
        .din(new_Jinkela_wire_3160),
        .dout(new_Jinkela_wire_3161)
    );

    bfr new_Jinkela_buffer_533 (
        .din(new_Jinkela_wire_957),
        .dout(new_Jinkela_wire_958)
    );

    bfr new_Jinkela_buffer_2010 (
        .din(new_Jinkela_wire_3185),
        .dout(new_Jinkela_wire_3186)
    );

    bfr new_Jinkela_buffer_537 (
        .din(new_Jinkela_wire_966),
        .dout(new_Jinkela_wire_967)
    );

    bfr new_Jinkela_buffer_1993 (
        .din(new_Jinkela_wire_3161),
        .dout(new_Jinkela_wire_3162)
    );

    bfr new_Jinkela_buffer_534 (
        .din(new_Jinkela_wire_958),
        .dout(new_Jinkela_wire_959)
    );

    spl3L new_Jinkela_splitter_457 (
        .a(_0319_),
        .d(new_Jinkela_wire_3208),
        .b(new_Jinkela_wire_3209),
        .c(new_Jinkela_wire_3210)
    );

    spl2 new_Jinkela_splitter_167 (
        .a(_0305_),
        .b(new_Jinkela_wire_970),
        .c(new_Jinkela_wire_972)
    );

    bfr new_Jinkela_buffer_2019 (
        .din(_0567_),
        .dout(new_Jinkela_wire_3204)
    );

    bfr new_Jinkela_buffer_541 (
        .din(_0675_),
        .dout(new_Jinkela_wire_977)
    );

    bfr new_Jinkela_buffer_2011 (
        .din(new_Jinkela_wire_3186),
        .dout(new_Jinkela_wire_3187)
    );

    bfr new_Jinkela_buffer_538 (
        .din(new_Jinkela_wire_967),
        .dout(new_Jinkela_wire_968)
    );

    spl3L new_Jinkela_splitter_456 (
        .a(_0545_),
        .d(new_Jinkela_wire_3200),
        .b(new_Jinkela_wire_3201),
        .c(new_Jinkela_wire_3202)
    );

    bfr new_Jinkela_buffer_551 (
        .din(_0151_),
        .dout(new_Jinkela_wire_987)
    );

    bfr new_Jinkela_buffer_2016 (
        .din(new_Jinkela_wire_3195),
        .dout(new_Jinkela_wire_3196)
    );

    bfr new_Jinkela_buffer_540 (
        .din(new_Jinkela_wire_970),
        .dout(new_Jinkela_wire_971)
    );

    spl4L new_Jinkela_splitter_168 (
        .a(new_Jinkela_wire_972),
        .d(new_Jinkela_wire_973),
        .e(new_Jinkela_wire_974),
        .b(new_Jinkela_wire_975),
        .c(new_Jinkela_wire_976)
    );

    bfr new_Jinkela_buffer_2018 (
        .din(new_Jinkela_wire_3202),
        .dout(new_Jinkela_wire_3203)
    );

    bfr new_Jinkela_buffer_549 (
        .din(_0046_),
        .dout(new_Jinkela_wire_985)
    );

    bfr new_Jinkela_buffer_2017 (
        .din(new_Jinkela_wire_3196),
        .dout(new_Jinkela_wire_3197)
    );

    bfr new_Jinkela_buffer_2020 (
        .din(new_Jinkela_wire_3204),
        .dout(new_Jinkela_wire_3205)
    );

    bfr new_Jinkela_buffer_553 (
        .din(_0615_),
        .dout(new_Jinkela_wire_991)
    );

    spl2 new_Jinkela_splitter_455 (
        .a(new_Jinkela_wire_3197),
        .b(new_Jinkela_wire_3198),
        .c(new_Jinkela_wire_3199)
    );

    bfr new_Jinkela_buffer_542 (
        .din(new_Jinkela_wire_977),
        .dout(new_Jinkela_wire_978)
    );

    bfr new_Jinkela_buffer_543 (
        .din(new_Jinkela_wire_978),
        .dout(new_Jinkela_wire_979)
    );

    bfr new_Jinkela_buffer_2030 (
        .din(_0628_),
        .dout(new_Jinkela_wire_3226)
    );

    bfr new_Jinkela_buffer_2025 (
        .din(_0562_),
        .dout(new_Jinkela_wire_3215)
    );

    bfr new_Jinkela_buffer_550 (
        .din(new_Jinkela_wire_985),
        .dout(new_Jinkela_wire_986)
    );

    bfr new_Jinkela_buffer_544 (
        .din(new_Jinkela_wire_979),
        .dout(new_Jinkela_wire_980)
    );

    bfr new_Jinkela_buffer_2021 (
        .din(new_Jinkela_wire_3205),
        .dout(new_Jinkela_wire_3206)
    );

    bfr new_Jinkela_buffer_552 (
        .din(new_Jinkela_wire_987),
        .dout(new_Jinkela_wire_988)
    );

    spl2 new_Jinkela_splitter_459 (
        .a(_0068_),
        .b(new_Jinkela_wire_3216),
        .c(new_Jinkela_wire_3218)
    );

    bfr new_Jinkela_buffer_545 (
        .din(new_Jinkela_wire_980),
        .dout(new_Jinkela_wire_981)
    );

    bfr new_Jinkela_buffer_2022 (
        .din(new_Jinkela_wire_3206),
        .dout(new_Jinkela_wire_3207)
    );

    bfr new_Jinkela_buffer_563 (
        .din(_0439_),
        .dout(new_Jinkela_wire_1001)
    );

    bfr new_Jinkela_buffer_2023 (
        .din(new_Jinkela_wire_3210),
        .dout(new_Jinkela_wire_3211)
    );

    bfr new_Jinkela_buffer_2027 (
        .din(new_Jinkela_wire_3222),
        .dout(new_Jinkela_wire_3223)
    );

    bfr new_Jinkela_buffer_546 (
        .din(new_Jinkela_wire_981),
        .dout(new_Jinkela_wire_982)
    );

    bfr new_Jinkela_buffer_2024 (
        .din(new_Jinkela_wire_3211),
        .dout(new_Jinkela_wire_3212)
    );

    bfr new_Jinkela_buffer_569 (
        .din(_0497_),
        .dout(new_Jinkela_wire_1009)
    );

    bfr new_Jinkela_buffer_547 (
        .din(new_Jinkela_wire_982),
        .dout(new_Jinkela_wire_983)
    );

    bfr new_Jinkela_buffer_2026 (
        .din(new_Jinkela_wire_3216),
        .dout(new_Jinkela_wire_3217)
    );

    spl4L new_Jinkela_splitter_460 (
        .a(new_Jinkela_wire_3218),
        .d(new_Jinkela_wire_3219),
        .e(new_Jinkela_wire_3220),
        .b(new_Jinkela_wire_3221),
        .c(new_Jinkela_wire_3222)
    );

    bfr new_Jinkela_buffer_554 (
        .din(new_Jinkela_wire_991),
        .dout(new_Jinkela_wire_992)
    );

    spl2 new_Jinkela_splitter_458 (
        .a(new_Jinkela_wire_3212),
        .b(new_Jinkela_wire_3213),
        .c(new_Jinkela_wire_3214)
    );

    spl2 new_Jinkela_splitter_169 (
        .a(new_Jinkela_wire_988),
        .b(new_Jinkela_wire_989),
        .c(new_Jinkela_wire_990)
    );

    bfr new_Jinkela_buffer_548 (
        .din(new_Jinkela_wire_983),
        .dout(new_Jinkela_wire_984)
    );

    bfr new_Jinkela_buffer_2032 (
        .din(_0633_),
        .dout(new_Jinkela_wire_3228)
    );

    bfr new_Jinkela_buffer_555 (
        .din(new_Jinkela_wire_992),
        .dout(new_Jinkela_wire_993)
    );

    bfr new_Jinkela_buffer_2031 (
        .din(new_Jinkela_wire_3226),
        .dout(new_Jinkela_wire_3227)
    );

    bfr new_Jinkela_buffer_580 (
        .din(_0411_),
        .dout(new_Jinkela_wire_1020)
    );

    spl4L new_Jinkela_splitter_461 (
        .a(_0000_),
        .d(new_Jinkela_wire_3229),
        .e(new_Jinkela_wire_3230),
        .b(new_Jinkela_wire_3231),
        .c(new_Jinkela_wire_3232)
    );

    bfr new_Jinkela_buffer_564 (
        .din(new_Jinkela_wire_1001),
        .dout(new_Jinkela_wire_1002)
    );

    bfr new_Jinkela_buffer_2033 (
        .din(_0737_),
        .dout(new_Jinkela_wire_3233)
    );

    bfr new_Jinkela_buffer_556 (
        .din(new_Jinkela_wire_993),
        .dout(new_Jinkela_wire_994)
    );

    bfr new_Jinkela_buffer_2028 (
        .din(new_Jinkela_wire_3223),
        .dout(new_Jinkela_wire_3224)
    );

    bfr new_Jinkela_buffer_185 (
        .din(new_Jinkela_wire_308),
        .dout(new_Jinkela_wire_309)
    );

    bfr new_Jinkela_buffer_180 (
        .din(new_Jinkela_wire_295),
        .dout(new_Jinkela_wire_296)
    );

    spl2 new_Jinkela_splitter_48 (
        .a(new_Jinkela_wire_324),
        .b(new_Jinkela_wire_325),
        .c(new_Jinkela_wire_326)
    );

    bfr new_Jinkela_buffer_181 (
        .din(new_Jinkela_wire_296),
        .dout(new_Jinkela_wire_297)
    );

    spl2 new_Jinkela_splitter_53 (
        .a(G48),
        .b(new_Jinkela_wire_343),
        .c(new_Jinkela_wire_344)
    );

    bfr new_Jinkela_buffer_182 (
        .din(new_Jinkela_wire_297),
        .dout(new_Jinkela_wire_298)
    );

    bfr new_Jinkela_buffer_186 (
        .din(new_Jinkela_wire_312),
        .dout(new_Jinkela_wire_313)
    );

    spl2 new_Jinkela_splitter_42 (
        .a(new_Jinkela_wire_298),
        .b(new_Jinkela_wire_299),
        .c(new_Jinkela_wire_300)
    );

    bfr new_Jinkela_buffer_183 (
        .din(new_Jinkela_wire_300),
        .dout(new_Jinkela_wire_301)
    );

    bfr new_Jinkela_buffer_187 (
        .din(new_Jinkela_wire_313),
        .dout(new_Jinkela_wire_314)
    );

    spl4L new_Jinkela_splitter_49 (
        .a(new_Jinkela_wire_327),
        .d(new_Jinkela_wire_328),
        .e(new_Jinkela_wire_329),
        .b(new_Jinkela_wire_330),
        .c(new_Jinkela_wire_331)
    );

    bfr new_Jinkela_buffer_188 (
        .din(new_Jinkela_wire_314),
        .dout(new_Jinkela_wire_315)
    );

    bfr new_Jinkela_buffer_199 (
        .din(new_Jinkela_wire_344),
        .dout(new_Jinkela_wire_345)
    );

    bfr new_Jinkela_buffer_189 (
        .din(new_Jinkela_wire_315),
        .dout(new_Jinkela_wire_316)
    );

    spl2 new_Jinkela_splitter_50 (
        .a(new_Jinkela_wire_331),
        .b(new_Jinkela_wire_332),
        .c(new_Jinkela_wire_333)
    );

    bfr new_Jinkela_buffer_190 (
        .din(new_Jinkela_wire_316),
        .dout(new_Jinkela_wire_317)
    );

    spl2 new_Jinkela_splitter_54 (
        .a(G22),
        .b(new_Jinkela_wire_391),
        .c(new_Jinkela_wire_392)
    );

    bfr new_Jinkela_buffer_191 (
        .din(new_Jinkela_wire_317),
        .dout(new_Jinkela_wire_318)
    );

    bfr new_Jinkela_buffer_200 (
        .din(new_Jinkela_wire_345),
        .dout(new_Jinkela_wire_346)
    );

    bfr new_Jinkela_buffer_192 (
        .din(new_Jinkela_wire_318),
        .dout(new_Jinkela_wire_319)
    );

    spl2 new_Jinkela_splitter_59 (
        .a(G4),
        .b(new_Jinkela_wire_407),
        .c(new_Jinkela_wire_410)
    );

    spl2 new_Jinkela_splitter_46 (
        .a(new_Jinkela_wire_319),
        .b(new_Jinkela_wire_320),
        .c(new_Jinkela_wire_321)
    );

    bfr new_Jinkela_buffer_193 (
        .din(new_Jinkela_wire_321),
        .dout(new_Jinkela_wire_322)
    );

    bfr new_Jinkela_buffer_250 (
        .din(new_Jinkela_wire_407),
        .dout(new_Jinkela_wire_408)
    );

    bfr new_Jinkela_buffer_194 (
        .din(new_Jinkela_wire_333),
        .dout(new_Jinkela_wire_334)
    );

    bfr new_Jinkela_buffer_201 (
        .din(new_Jinkela_wire_346),
        .dout(new_Jinkela_wire_347)
    );

    spl2 new_Jinkela_splitter_51 (
        .a(new_Jinkela_wire_334),
        .b(new_Jinkela_wire_335),
        .c(new_Jinkela_wire_336)
    );

    bfr new_Jinkela_buffer_195 (
        .din(new_Jinkela_wire_336),
        .dout(new_Jinkela_wire_337)
    );

    bfr new_Jinkela_buffer_260 (
        .din(G17),
        .dout(new_Jinkela_wire_461)
    );

    bfr new_Jinkela_buffer_261 (
        .din(new_Jinkela_wire_461),
        .dout(new_Jinkela_wire_462)
    );

    bfr new_Jinkela_buffer_202 (
        .din(new_Jinkela_wire_347),
        .dout(new_Jinkela_wire_348)
    );

    spl2 new_Jinkela_splitter_52 (
        .a(new_Jinkela_wire_337),
        .b(new_Jinkela_wire_338),
        .c(new_Jinkela_wire_339)
    );

    bfr new_Jinkela_buffer_196 (
        .din(new_Jinkela_wire_339),
        .dout(new_Jinkela_wire_340)
    );

    bfr new_Jinkela_buffer_245 (
        .din(new_Jinkela_wire_395),
        .dout(new_Jinkela_wire_396)
    );

    bfr new_Jinkela_buffer_203 (
        .din(new_Jinkela_wire_348),
        .dout(new_Jinkela_wire_349)
    );

    bfr new_Jinkela_buffer_197 (
        .din(new_Jinkela_wire_340),
        .dout(new_Jinkela_wire_341)
    );

    spl3L new_Jinkela_splitter_55 (
        .a(new_Jinkela_wire_392),
        .d(new_Jinkela_wire_393),
        .b(new_Jinkela_wire_394),
        .c(new_Jinkela_wire_395)
    );

    bfr new_Jinkela_buffer_198 (
        .din(new_Jinkela_wire_341),
        .dout(new_Jinkela_wire_342)
    );

    bfr new_Jinkela_buffer_204 (
        .din(new_Jinkela_wire_349),
        .dout(new_Jinkela_wire_350)
    );

    bfr new_Jinkela_buffer_268 (
        .din(new_Jinkela_wire_473),
        .dout(new_Jinkela_wire_474)
    );

    spl4L new_Jinkela_splitter_60 (
        .a(new_Jinkela_wire_410),
        .d(new_Jinkela_wire_411),
        .e(new_Jinkela_wire_416),
        .b(new_Jinkela_wire_421),
        .c(new_Jinkela_wire_426)
    );

    bfr new_Jinkela_buffer_205 (
        .din(new_Jinkela_wire_350),
        .dout(new_Jinkela_wire_351)
    );

    and_ii _0869_ (
        .a(_0041_),
        .b(_0040_),
        .c(_0042_)
    );

    and_bb _1583_ (
        .a(new_Jinkela_wire_1491),
        .b(new_Jinkela_wire_1671),
        .c(_0755_)
    );

    or_bb _0870_ (
        .a(new_Jinkela_wire_1930),
        .b(new_Jinkela_wire_1626),
        .c(_0043_)
    );

    and_bi _1584_ (
        .a(_0754_),
        .b(_0755_),
        .c(new_net_1469)
    );

    and_bb _0871_ (
        .a(new_Jinkela_wire_1929),
        .b(new_Jinkela_wire_1625),
        .c(_0044_)
    );

    and_bi _1585_ (
        .a(new_Jinkela_wire_2309),
        .b(new_Jinkela_wire_3135),
        .c(new_net_1467)
    );

    and_bi _0872_ (
        .a(_0043_),
        .b(_0044_),
        .c(new_net_1463)
    );

    and_bi _1586_ (
        .a(new_Jinkela_wire_2313),
        .b(new_Jinkela_wire_1724),
        .c(new_net_1471)
    );

    and_bi _0873_ (
        .a(new_Jinkela_wire_160),
        .b(new_Jinkela_wire_2509),
        .c(_0045_)
    );

    and_bi _1587_ (
        .a(new_Jinkela_wire_2943),
        .b(new_Jinkela_wire_2647),
        .c(_0757_)
    );

    or_bb _0874_ (
        .a(new_Jinkela_wire_3304),
        .b(new_Jinkela_wire_582),
        .c(_0046_)
    );

    and_bi _1588_ (
        .a(new_Jinkela_wire_2891),
        .b(new_Jinkela_wire_626),
        .c(_0758_)
    );

    and_bi _0875_ (
        .a(new_Jinkela_wire_154),
        .b(new_Jinkela_wire_599),
        .c(_0047_)
    );

    or_bb _1589_ (
        .a(_0758_),
        .b(new_Jinkela_wire_1227),
        .c(new_net_1483)
    );

    or_ii _0876_ (
        .a(new_Jinkela_wire_793),
        .b(new_Jinkela_wire_589),
        .c(_0048_)
    );

    or_ii _1590_ (
        .a(new_Jinkela_wire_953),
        .b(new_Jinkela_wire_2315),
        .c(_0759_)
    );

    or_ii _0877_ (
        .a(new_Jinkela_wire_597),
        .b(new_Jinkela_wire_157),
        .c(_0049_)
    );

    and_bi _1591_ (
        .a(new_Jinkela_wire_2073),
        .b(new_Jinkela_wire_952),
        .c(_0760_)
    );

    and_bi _0878_ (
        .a(new_Jinkela_wire_433),
        .b(_0049_),
        .c(_0050_)
    );

    and_bi _1592_ (
        .a(_0759_),
        .b(_0760_),
        .c(_0761_)
    );

    or_bi _0879_ (
        .a(_0050_),
        .b(new_Jinkela_wire_1466),
        .c(_0051_)
    );

    and_bi _1593_ (
        .a(new_Jinkela_wire_973),
        .b(new_Jinkela_wire_2751),
        .c(_0762_)
    );

    and_ii _0880_ (
        .a(new_Jinkela_wire_3311),
        .b(new_Jinkela_wire_3261),
        .c(_0052_)
    );

    and_bi _1594_ (
        .a(new_Jinkela_wire_2710),
        .b(new_Jinkela_wire_905),
        .c(_0763_)
    );

    and_bi _0881_ (
        .a(new_Jinkela_wire_586),
        .b(new_Jinkela_wire_2167),
        .c(_0053_)
    );

    and_bi _1595_ (
        .a(new_Jinkela_wire_904),
        .b(new_Jinkela_wire_2711),
        .c(_0765_)
    );

    and_bi _0882_ (
        .a(new_Jinkela_wire_986),
        .b(_0053_),
        .c(_0054_)
    );

    and_ii _1596_ (
        .a(_0765_),
        .b(_0763_),
        .c(_0766_)
    );

    and_bi _0883_ (
        .a(new_Jinkela_wire_2306),
        .b(new_Jinkela_wire_578),
        .c(_0055_)
    );

    or_ii _1597_ (
        .a(new_Jinkela_wire_3013),
        .b(new_Jinkela_wire_1235),
        .c(_0767_)
    );

    or_bb _0884_ (
        .a(_0055_),
        .b(new_Jinkela_wire_2948),
        .c(_0056_)
    );

    or_bb _1598_ (
        .a(new_Jinkela_wire_3012),
        .b(new_Jinkela_wire_1234),
        .c(_0768_)
    );

    or_bb _0885_ (
        .a(new_Jinkela_wire_444),
        .b(new_Jinkela_wire_161),
        .c(_0057_)
    );

    or_ii _1599_ (
        .a(_0768_),
        .b(_0767_),
        .c(_0769_)
    );

    and_bi _0886_ (
        .a(new_Jinkela_wire_495),
        .b(new_Jinkela_wire_1280),
        .c(_0058_)
    );

    and_ii _1600_ (
        .a(new_Jinkela_wire_795),
        .b(new_Jinkela_wire_588),
        .c(_0770_)
    );

    inv _0887_ (
        .din(new_Jinkela_wire_264),
        .dout(_0059_)
    );

    or_bb _1601_ (
        .a(new_Jinkela_wire_1863),
        .b(new_Jinkela_wire_3322),
        .c(_0771_)
    );

    or_bi _0888_ (
        .a(new_Jinkela_wire_162),
        .b(new_Jinkela_wire_432),
        .c(_0060_)
    );

    and_bi _1602_ (
        .a(_0769_),
        .b(new_Jinkela_wire_1979),
        .c(_0772_)
    );

    and_bi _0889_ (
        .a(new_Jinkela_wire_1056),
        .b(new_Jinkela_wire_3332),
        .c(_0061_)
    );

    or_bi _1603_ (
        .a(new_Jinkela_wire_199),
        .b(new_Jinkela_wire_576),
        .c(_0773_)
    );

    or_bb _0890_ (
        .a(_0061_),
        .b(new_Jinkela_wire_1728),
        .c(_0062_)
    );

    and_ii _1604_ (
        .a(new_Jinkela_wire_3137),
        .b(new_Jinkela_wire_2777),
        .c(_0774_)
    );

    and_bi _0891_ (
        .a(new_Jinkela_wire_2733),
        .b(_0062_),
        .c(_0063_)
    );

    and_bi _1605_ (
        .a(new_Jinkela_wire_1371),
        .b(_0774_),
        .c(_0776_)
    );

    and_bi _0892_ (
        .a(new_Jinkela_wire_3319),
        .b(_0063_),
        .c(_0064_)
    );

    and_bi _1606_ (
        .a(new_Jinkela_wire_1867),
        .b(_0776_),
        .c(_0777_)
    );

    or_bb _0893_ (
        .a(_0064_),
        .b(_0054_),
        .c(_0065_)
    );

    or_ii _1607_ (
        .a(new_Jinkela_wire_2644),
        .b(new_Jinkela_wire_2392),
        .c(_0778_)
    );

    or_bb _0894_ (
        .a(new_Jinkela_wire_561),
        .b(new_Jinkela_wire_0),
        .c(_0066_)
    );

    and_bi _1608_ (
        .a(new_Jinkela_wire_806),
        .b(_0778_),
        .c(_0779_)
    );

    or_bb _0895_ (
        .a(new_Jinkela_wire_535),
        .b(new_Jinkela_wire_633),
        .c(_0067_)
    );

    or_bb _1609_ (
        .a(new_Jinkela_wire_3288),
        .b(_0777_),
        .c(_0780_)
    );

    and_bi _0896_ (
        .a(new_Jinkela_wire_3291),
        .b(new_Jinkela_wire_598),
        .c(_0068_)
    );

    or_bb _1610_ (
        .a(new_Jinkela_wire_2868),
        .b(_0772_),
        .c(new_net_1485)
    );

    and_bb _0897_ (
        .a(new_Jinkela_wire_420),
        .b(new_Jinkela_wire_538),
        .c(_0069_)
    );

    or_ii _1611_ (
        .a(new_Jinkela_wire_1668),
        .b(new_Jinkela_wire_94),
        .c(_0781_)
    );

    or_bb _0898_ (
        .a(new_Jinkela_wire_1284),
        .b(new_Jinkela_wire_1465),
        .c(_0070_)
    );

    and_ii _1612_ (
        .a(new_Jinkela_wire_1667),
        .b(new_Jinkela_wire_93),
        .c(_0782_)
    );

    or_ii _0899_ (
        .a(new_Jinkela_wire_1039),
        .b(new_Jinkela_wire_560),
        .c(_0071_)
    );

    or_bi _1613_ (
        .a(_0782_),
        .b(new_Jinkela_wire_2264),
        .c(_0783_)
    );

    and_bi _0900_ (
        .a(new_Jinkela_wire_3225),
        .b(new_Jinkela_wire_2166),
        .c(_0072_)
    );

    and_bi _1614_ (
        .a(new_Jinkela_wire_3036),
        .b(_0783_),
        .c(_0784_)
    );

    or_bi _0901_ (
        .a(new_Jinkela_wire_3217),
        .b(new_Jinkela_wire_43),
        .c(_0073_)
    );

    or_ii _1615_ (
        .a(new_Jinkela_wire_1272),
        .b(new_Jinkela_wire_1494),
        .c(_0786_)
    );

    or_bb _0902_ (
        .a(new_Jinkela_wire_790),
        .b(new_Jinkela_wire_414),
        .c(_0074_)
    );

    or_bb _1616_ (
        .a(new_Jinkela_wire_1271),
        .b(new_Jinkela_wire_1495),
        .c(_0787_)
    );

    and_bi _0903_ (
        .a(new_Jinkela_wire_632),
        .b(new_Jinkela_wire_3034),
        .c(_0075_)
    );

    or_ii _1617_ (
        .a(_0787_),
        .b(_0786_),
        .c(G3539)
    );

    or_bi _0904_ (
        .a(new_Jinkela_wire_428),
        .b(new_Jinkela_wire_742),
        .c(_0076_)
    );

    or_ii _0905_ (
        .a(new_Jinkela_wire_750),
        .b(new_Jinkela_wire_423),
        .c(_0077_)
    );

    or_ii _0906_ (
        .a(new_Jinkela_wire_1398),
        .b(new_Jinkela_wire_2639),
        .c(_0078_)
    );

    or_bb _0907_ (
        .a(_0078_),
        .b(_0075_),
        .c(_0079_)
    );

    and_bi _0908_ (
        .a(new_Jinkela_wire_1329),
        .b(_0079_),
        .c(_0080_)
    );

    and_bi _0909_ (
        .a(new_Jinkela_wire_1042),
        .b(_0080_),
        .c(_0081_)
    );

    or_bb _0910_ (
        .a(new_Jinkela_wire_2457),
        .b(new_Jinkela_wire_838),
        .c(_0082_)
    );

    bfr new_Jinkela_buffer_0 (
        .din(new_Jinkela_wire_1),
        .dout(new_Jinkela_wire_2)
    );

    spl2 new_Jinkela_splitter_0 (
        .a(G25),
        .b(new_Jinkela_wire_0),
        .c(new_Jinkela_wire_1)
    );

    spl2 new_Jinkela_splitter_1 (
        .a(G47),
        .b(new_Jinkela_wire_3),
        .c(new_Jinkela_wire_4)
    );

    bfr new_Jinkela_buffer_26 (
        .din(G30),
        .dout(new_Jinkela_wire_34)
    );

    spl2 new_Jinkela_splitter_9 (
        .a(G3),
        .b(new_Jinkela_wire_146),
        .c(new_Jinkela_wire_150)
    );

    bfr new_Jinkela_buffer_1 (
        .din(new_Jinkela_wire_4),
        .dout(new_Jinkela_wire_5)
    );

    bfr new_Jinkela_buffer_2 (
        .din(new_Jinkela_wire_5),
        .dout(new_Jinkela_wire_6)
    );

    spl2 new_Jinkela_splitter_7 (
        .a(G27),
        .b(new_Jinkela_wire_95),
        .c(new_Jinkela_wire_96)
    );

    spl2 new_Jinkela_splitter_4 (
        .a(new_Jinkela_wire_38),
        .b(new_Jinkela_wire_39),
        .c(new_Jinkela_wire_40)
    );

    bfr new_Jinkela_buffer_3 (
        .din(new_Jinkela_wire_6),
        .dout(new_Jinkela_wire_7)
    );

    bfr new_Jinkela_buffer_30 (
        .din(new_Jinkela_wire_45),
        .dout(new_Jinkela_wire_46)
    );

    bfr new_Jinkela_buffer_4 (
        .din(new_Jinkela_wire_7),
        .dout(new_Jinkela_wire_8)
    );

    bfr new_Jinkela_buffer_5 (
        .din(new_Jinkela_wire_8),
        .dout(new_Jinkela_wire_9)
    );

    bfr new_Jinkela_buffer_27 (
        .din(new_Jinkela_wire_40),
        .dout(new_Jinkela_wire_41)
    );

    bfr new_Jinkela_buffer_6 (
        .din(new_Jinkela_wire_9),
        .dout(new_Jinkela_wire_10)
    );

    bfr new_Jinkela_buffer_29 (
        .din(G50),
        .dout(new_Jinkela_wire_45)
    );

    spl4L new_Jinkela_splitter_3 (
        .a(new_Jinkela_wire_34),
        .d(new_Jinkela_wire_35),
        .e(new_Jinkela_wire_36),
        .b(new_Jinkela_wire_37),
        .c(new_Jinkela_wire_38)
    );

    bfr new_Jinkela_buffer_474 (
        .din(new_Jinkela_wire_867),
        .dout(new_Jinkela_wire_868)
    );

    bfr new_Jinkela_buffer_520 (
        .din(_0470_),
        .dout(new_Jinkela_wire_938)
    );

    bfr new_Jinkela_buffer_475 (
        .din(new_Jinkela_wire_868),
        .dout(new_Jinkela_wire_869)
    );

    bfr new_Jinkela_buffer_476 (
        .din(new_Jinkela_wire_869),
        .dout(new_Jinkela_wire_870)
    );

    bfr new_Jinkela_buffer_513 (
        .din(new_Jinkela_wire_921),
        .dout(new_Jinkela_wire_922)
    );

    bfr new_Jinkela_buffer_512 (
        .din(new_Jinkela_wire_920),
        .dout(new_Jinkela_wire_921)
    );

    bfr new_Jinkela_buffer_477 (
        .din(new_Jinkela_wire_870),
        .dout(new_Jinkela_wire_871)
    );

    spl2 new_Jinkela_splitter_161 (
        .a(_0082_),
        .b(new_Jinkela_wire_936),
        .c(new_Jinkela_wire_937)
    );

    spl2 new_Jinkela_splitter_163 (
        .a(_0732_),
        .b(new_Jinkela_wire_942),
        .c(new_Jinkela_wire_943)
    );

    bfr new_Jinkela_buffer_478 (
        .din(new_Jinkela_wire_871),
        .dout(new_Jinkela_wire_872)
    );

    spl2 new_Jinkela_splitter_158 (
        .a(new_Jinkela_wire_922),
        .b(new_Jinkela_wire_923),
        .c(new_Jinkela_wire_924)
    );

    bfr new_Jinkela_buffer_521 (
        .din(new_Jinkela_wire_938),
        .dout(new_Jinkela_wire_939)
    );

    bfr new_Jinkela_buffer_479 (
        .din(new_Jinkela_wire_872),
        .dout(new_Jinkela_wire_873)
    );

    bfr new_Jinkela_buffer_480 (
        .din(new_Jinkela_wire_873),
        .dout(new_Jinkela_wire_874)
    );

    bfr new_Jinkela_buffer_514 (
        .din(new_Jinkela_wire_924),
        .dout(new_Jinkela_wire_925)
    );

    bfr new_Jinkela_buffer_481 (
        .din(new_Jinkela_wire_874),
        .dout(new_Jinkela_wire_875)
    );

    bfr new_Jinkela_buffer_482 (
        .din(new_Jinkela_wire_875),
        .dout(new_Jinkela_wire_876)
    );

    spl2 new_Jinkela_splitter_162 (
        .a(_0327_),
        .b(new_Jinkela_wire_940),
        .c(new_Jinkela_wire_941)
    );

    bfr new_Jinkela_buffer_483 (
        .din(new_Jinkela_wire_876),
        .dout(new_Jinkela_wire_877)
    );

    spl3L new_Jinkela_splitter_159 (
        .a(new_Jinkela_wire_925),
        .d(new_Jinkela_wire_926),
        .b(new_Jinkela_wire_927),
        .c(new_Jinkela_wire_928)
    );

    bfr new_Jinkela_buffer_484 (
        .din(new_Jinkela_wire_877),
        .dout(new_Jinkela_wire_878)
    );

    bfr new_Jinkela_buffer_485 (
        .din(new_Jinkela_wire_878),
        .dout(new_Jinkela_wire_879)
    );

    bfr new_Jinkela_buffer_515 (
        .din(new_Jinkela_wire_928),
        .dout(new_Jinkela_wire_929)
    );

    bfr new_Jinkela_buffer_486 (
        .din(new_Jinkela_wire_879),
        .dout(new_Jinkela_wire_880)
    );

    bfr new_Jinkela_buffer_527 (
        .din(_0638_),
        .dout(new_Jinkela_wire_949)
    );

    bfr new_Jinkela_buffer_487 (
        .din(new_Jinkela_wire_880),
        .dout(new_Jinkela_wire_881)
    );

    bfr new_Jinkela_buffer_516 (
        .din(new_Jinkela_wire_929),
        .dout(new_Jinkela_wire_930)
    );

    bfr new_Jinkela_buffer_488 (
        .din(new_Jinkela_wire_881),
        .dout(new_Jinkela_wire_882)
    );

    bfr new_Jinkela_buffer_522 (
        .din(new_Jinkela_wire_943),
        .dout(new_Jinkela_wire_944)
    );

    bfr new_Jinkela_buffer_489 (
        .din(new_Jinkela_wire_882),
        .dout(new_Jinkela_wire_883)
    );

    bfr new_Jinkela_buffer_517 (
        .din(new_Jinkela_wire_930),
        .dout(new_Jinkela_wire_931)
    );

    bfr new_Jinkela_buffer_490 (
        .din(new_Jinkela_wire_883),
        .dout(new_Jinkela_wire_884)
    );

    spl3L new_Jinkela_splitter_164 (
        .a(_0321_),
        .d(new_Jinkela_wire_952),
        .b(new_Jinkela_wire_953),
        .c(new_Jinkela_wire_954)
    );

    spl2 new_Jinkela_splitter_165 (
        .a(_0328_),
        .b(new_Jinkela_wire_960),
        .c(new_Jinkela_wire_961)
    );

    bfr new_Jinkela_buffer_491 (
        .din(new_Jinkela_wire_884),
        .dout(new_Jinkela_wire_885)
    );

    bfr new_Jinkela_buffer_518 (
        .din(new_Jinkela_wire_931),
        .dout(new_Jinkela_wire_932)
    );

    bfr new_Jinkela_buffer_492 (
        .din(new_Jinkela_wire_885),
        .dout(new_Jinkela_wire_886)
    );

    bfr new_Jinkela_buffer_528 (
        .din(new_Jinkela_wire_949),
        .dout(new_Jinkela_wire_950)
    );

    bfr new_Jinkela_buffer_523 (
        .din(new_Jinkela_wire_944),
        .dout(new_Jinkela_wire_945)
    );

    bfr new_Jinkela_buffer_493 (
        .din(new_Jinkela_wire_886),
        .dout(new_Jinkela_wire_887)
    );

    bfr new_Jinkela_buffer_494 (
        .din(new_Jinkela_wire_887),
        .dout(new_Jinkela_wire_888)
    );

    bfr new_Jinkela_buffer_2046 (
        .din(_0511_),
        .dout(new_Jinkela_wire_3248)
    );

    bfr new_Jinkela_buffer_2029 (
        .din(new_Jinkela_wire_3224),
        .dout(new_Jinkela_wire_3225)
    );

    bfr new_Jinkela_buffer_2035 (
        .din(_0325_),
        .dout(new_Jinkela_wire_3235)
    );

    bfr new_Jinkela_buffer_2034 (
        .din(new_Jinkela_wire_3233),
        .dout(new_Jinkela_wire_3234)
    );

    spl2 new_Jinkela_splitter_463 (
        .a(_0160_),
        .b(new_Jinkela_wire_3254),
        .c(new_Jinkela_wire_3255)
    );

    bfr new_Jinkela_buffer_2036 (
        .din(new_Jinkela_wire_3235),
        .dout(new_Jinkela_wire_3236)
    );

    spl2 new_Jinkela_splitter_464 (
        .a(_0742_),
        .b(new_Jinkela_wire_3256),
        .c(new_Jinkela_wire_3257)
    );

    bfr new_Jinkela_buffer_2047 (
        .din(new_Jinkela_wire_3248),
        .dout(new_Jinkela_wire_3249)
    );

    bfr new_Jinkela_buffer_2037 (
        .din(new_Jinkela_wire_3236),
        .dout(new_Jinkela_wire_3237)
    );

    spl2 new_Jinkela_splitter_462 (
        .a(new_Jinkela_wire_3237),
        .b(new_Jinkela_wire_3238),
        .c(new_Jinkela_wire_3239)
    );

    bfr new_Jinkela_buffer_2038 (
        .din(new_Jinkela_wire_3239),
        .dout(new_Jinkela_wire_3240)
    );

    bfr new_Jinkela_buffer_2048 (
        .din(new_Jinkela_wire_3249),
        .dout(new_Jinkela_wire_3250)
    );

    bfr new_Jinkela_buffer_2039 (
        .din(new_Jinkela_wire_3240),
        .dout(new_Jinkela_wire_3241)
    );

    bfr new_Jinkela_buffer_2049 (
        .din(new_Jinkela_wire_3250),
        .dout(new_Jinkela_wire_3251)
    );

    bfr new_Jinkela_buffer_2040 (
        .din(new_Jinkela_wire_3241),
        .dout(new_Jinkela_wire_3242)
    );

    spl2 new_Jinkela_splitter_465 (
        .a(_0047_),
        .b(new_Jinkela_wire_3258),
        .c(new_Jinkela_wire_3259)
    );

    bfr new_Jinkela_buffer_2041 (
        .din(new_Jinkela_wire_3242),
        .dout(new_Jinkela_wire_3243)
    );

    bfr new_Jinkela_buffer_2050 (
        .din(new_Jinkela_wire_3251),
        .dout(new_Jinkela_wire_3252)
    );

    bfr new_Jinkela_buffer_2042 (
        .din(new_Jinkela_wire_3243),
        .dout(new_Jinkela_wire_3244)
    );

    bfr new_Jinkela_buffer_2054 (
        .din(_0358_),
        .dout(new_Jinkela_wire_3262)
    );

    bfr new_Jinkela_buffer_2043 (
        .din(new_Jinkela_wire_3244),
        .dout(new_Jinkela_wire_3245)
    );

    bfr new_Jinkela_buffer_2052 (
        .din(new_Jinkela_wire_3259),
        .dout(new_Jinkela_wire_3260)
    );

    bfr new_Jinkela_buffer_2051 (
        .din(new_Jinkela_wire_3252),
        .dout(new_Jinkela_wire_3253)
    );

    bfr new_Jinkela_buffer_2044 (
        .din(new_Jinkela_wire_3245),
        .dout(new_Jinkela_wire_3246)
    );

    bfr new_Jinkela_buffer_2055 (
        .din(new_net_3),
        .dout(new_Jinkela_wire_3263)
    );

    bfr new_Jinkela_buffer_2045 (
        .din(new_Jinkela_wire_3246),
        .dout(new_Jinkela_wire_3247)
    );

    spl3L new_Jinkela_splitter_467 (
        .a(_0631_),
        .d(new_Jinkela_wire_3285),
        .b(new_Jinkela_wire_3286),
        .c(new_Jinkela_wire_3287)
    );

    bfr new_Jinkela_buffer_2053 (
        .din(new_Jinkela_wire_3260),
        .dout(new_Jinkela_wire_3261)
    );

    bfr new_Jinkela_buffer_2074 (
        .din(_0779_),
        .dout(new_Jinkela_wire_3288)
    );

    bfr new_Jinkela_buffer_2056 (
        .din(new_Jinkela_wire_3263),
        .dout(new_Jinkela_wire_3264)
    );

    bfr new_Jinkela_buffer_2075 (
        .din(_0523_),
        .dout(new_Jinkela_wire_3289)
    );

    bfr new_Jinkela_buffer_2057 (
        .din(new_Jinkela_wire_3264),
        .dout(new_Jinkela_wire_3265)
    );

    bfr new_Jinkela_buffer_2058 (
        .din(new_Jinkela_wire_3265),
        .dout(new_Jinkela_wire_3266)
    );

    bfr new_Jinkela_buffer_2077 (
        .din(_0067_),
        .dout(new_Jinkela_wire_3291)
    );

    bfr new_Jinkela_buffer_2076 (
        .din(new_Jinkela_wire_3289),
        .dout(new_Jinkela_wire_3290)
    );

    bfr new_Jinkela_buffer_2059 (
        .din(new_Jinkela_wire_3266),
        .dout(new_Jinkela_wire_3267)
    );

    bfr new_Jinkela_buffer_2078 (
        .din(_0637_),
        .dout(new_Jinkela_wire_3292)
    );

    bfr new_Jinkela_buffer_2060 (
        .din(new_Jinkela_wire_3267),
        .dout(new_Jinkela_wire_3268)
    );

    spl2 new_Jinkela_splitter_468 (
        .a(_0045_),
        .b(new_Jinkela_wire_3298),
        .c(new_Jinkela_wire_3303)
    );

    bfr new_Jinkela_buffer_2061 (
        .din(new_Jinkela_wire_3268),
        .dout(new_Jinkela_wire_3269)
    );

    bfr new_Jinkela_buffer_2084 (
        .din(_0491_),
        .dout(new_Jinkela_wire_3308)
    );

    bfr new_Jinkela_buffer_2079 (
        .din(new_Jinkela_wire_3292),
        .dout(new_Jinkela_wire_3293)
    );

    bfr new_Jinkela_buffer_2062 (
        .din(new_Jinkela_wire_3269),
        .dout(new_Jinkela_wire_3270)
    );

    and_ii _1247_ (
        .a(new_Jinkela_wire_1176),
        .b(new_Jinkela_wire_2427),
        .c(_0417_)
    );

    and_bi _1248_ (
        .a(new_Jinkela_wire_764),
        .b(new_Jinkela_wire_2348),
        .c(_0418_)
    );

    and_bi _1249_ (
        .a(new_Jinkela_wire_676),
        .b(new_Jinkela_wire_3006),
        .c(_0419_)
    );

    or_bb _1250_ (
        .a(_0419_),
        .b(new_Jinkela_wire_2728),
        .c(_0420_)
    );

    and_bi _1251_ (
        .a(new_Jinkela_wire_469),
        .b(new_Jinkela_wire_1881),
        .c(_0421_)
    );

    or_bb _1252_ (
        .a(new_Jinkela_wire_791),
        .b(new_Jinkela_wire_178),
        .c(_0422_)
    );

    and_bi _1253_ (
        .a(new_Jinkela_wire_1513),
        .b(new_Jinkela_wire_1129),
        .c(_0423_)
    );

    or_bb _1254_ (
        .a(_0423_),
        .b(new_Jinkela_wire_1917),
        .c(_0424_)
    );

    or_bi _1255_ (
        .a(new_Jinkela_wire_1751),
        .b(new_Jinkela_wire_497),
        .c(_0425_)
    );

    or_ii _1256_ (
        .a(_0425_),
        .b(new_Jinkela_wire_1288),
        .c(_0426_)
    );

    or_bb _1257_ (
        .a(new_Jinkela_wire_2962),
        .b(_0424_),
        .c(_0427_)
    );

    or_bb _1258_ (
        .a(new_Jinkela_wire_1762),
        .b(_0420_),
        .c(_0428_)
    );

    or_bb _1259_ (
        .a(_0428_),
        .b(new_Jinkela_wire_1576),
        .c(_0429_)
    );

    and_bi _1260_ (
        .a(new_Jinkela_wire_2769),
        .b(new_Jinkela_wire_3010),
        .c(_0430_)
    );

    and_bi _1261_ (
        .a(new_Jinkela_wire_552),
        .b(new_Jinkela_wire_2175),
        .c(_0431_)
    );

    and_bi _1262_ (
        .a(new_Jinkela_wire_1940),
        .b(new_Jinkela_wire_1740),
        .c(_0432_)
    );

    and_bi _1263_ (
        .a(new_Jinkela_wire_2399),
        .b(new_Jinkela_wire_2369),
        .c(_0433_)
    );

    or_bb _1264_ (
        .a(_0433_),
        .b(new_Jinkela_wire_3183),
        .c(_0434_)
    );

    and_bi _1265_ (
        .a(new_Jinkela_wire_927),
        .b(new_Jinkela_wire_1877),
        .c(_0435_)
    );

    and_bi _1266_ (
        .a(new_Jinkela_wire_1717),
        .b(new_Jinkela_wire_2417),
        .c(_0436_)
    );

    or_bb _1267_ (
        .a(new_Jinkela_wire_2317),
        .b(new_Jinkela_wire_2649),
        .c(_0437_)
    );

    or_bb _1268_ (
        .a(_0437_),
        .b(_0434_),
        .c(_0438_)
    );

    and_bi _1269_ (
        .a(new_Jinkela_wire_328),
        .b(new_Jinkela_wire_234),
        .c(_0439_)
    );

    and_ii _1270_ (
        .a(new_Jinkela_wire_1008),
        .b(new_Jinkela_wire_1136),
        .c(_0440_)
    );

    and_bi _1271_ (
        .a(new_Jinkela_wire_1062),
        .b(new_Jinkela_wire_2430),
        .c(_0441_)
    );

    or_bb _1272_ (
        .a(_0441_),
        .b(new_Jinkela_wire_452),
        .c(_0442_)
    );

    or_bb _1273_ (
        .a(new_Jinkela_wire_1088),
        .b(new_Jinkela_wire_2734),
        .c(_0443_)
    );

    or_bb _1274_ (
        .a(_0443_),
        .b(_0438_),
        .c(_0444_)
    );

    and_bi _1275_ (
        .a(_0431_),
        .b(new_Jinkela_wire_1070),
        .c(_0445_)
    );

    and_bi _1276_ (
        .a(_0429_),
        .b(_0445_),
        .c(_0446_)
    );

    and_bi _1277_ (
        .a(new_Jinkela_wire_1913),
        .b(_0446_),
        .c(_0447_)
    );

    or_bb _1278_ (
        .a(_0447_),
        .b(new_Jinkela_wire_1346),
        .c(_0448_)
    );

    and_bi _1279_ (
        .a(_0415_),
        .b(new_Jinkela_wire_1268),
        .c(_0449_)
    );

    and_bi _1280_ (
        .a(new_Jinkela_wire_1503),
        .b(new_Jinkela_wire_2024),
        .c(_0450_)
    );

    and_bi _1281_ (
        .a(new_Jinkela_wire_2077),
        .b(new_Jinkela_wire_2021),
        .c(_0451_)
    );

    and_bi _1282_ (
        .a(new_Jinkela_wire_1560),
        .b(_0451_),
        .c(_0452_)
    );

    and_bi _1283_ (
        .a(new_Jinkela_wire_2119),
        .b(new_Jinkela_wire_2458),
        .c(_0453_)
    );

    or_bb _1284_ (
        .a(_0453_),
        .b(new_Jinkela_wire_2549),
        .c(_0454_)
    );

    and_bb _1285_ (
        .a(new_Jinkela_wire_2505),
        .b(new_Jinkela_wire_2285),
        .c(_0455_)
    );

    and_ii _1286_ (
        .a(new_Jinkela_wire_2720),
        .b(new_Jinkela_wire_960),
        .c(_0456_)
    );

    or_bi _1287_ (
        .a(new_Jinkela_wire_900),
        .b(new_Jinkela_wire_2935),
        .c(_0457_)
    );

    and_bi _1288_ (
        .a(new_Jinkela_wire_901),
        .b(new_Jinkela_wire_2936),
        .c(_0458_)
    );

endmodule
