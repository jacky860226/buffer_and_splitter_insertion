module c880(N1, N8, N13, N17, N26, N29, N36, N42, N51, N55, N59, N68, N72, N73, N74, N75, N80, N85, N86, N87, N88, N89, N90, N91, N96, N101, N106, N111, N116, N121, N126, N130, N135, N138, N143, N146, N149, N152, N153, N156, N159, N165, N171, N177, N183, N189, N195, N201, N207, N210, N219, N228, N237, N246, N255, N259, N260, N261, N267, N268, N388, N389, N390, N391, N418, N419, N420, N421, N422, N423, N446, N447, N448, N449, N450, N767, N768, N850, N863, N864, N865, N866, N874, N878, N879, N880);
	wire new_net_1907;
	wire new_net_1796;
	wire new_net_2032;
	wire new_net_1718;
	wire new_net_2074;
	wire new_net_217;
	wire new_net_2038;
	wire _009_;
	wire _093_;
	wire _177_;
	wire _219_;
	wire new_net_23;
	wire new_net_56;
	wire new_net_278;
	wire new_net_798;
	wire new_net_810;
	wire new_net_605;
	wire new_net_1441;
	wire new_net_1893;
	wire new_net_1236;
	wire new_net_2060;
	wire new_net_1933;
	wire new_net_159;
	wire new_net_210;
	wire new_net_396;
	wire new_net_454;
	wire new_net_1103;
	wire new_net_1365;
	wire new_net_1528;
	wire new_net_1839;
	wire new_net_1508;
	wire new_net_1968;
	wire new_net_1864;
	wire new_net_1501;
	wire new_net_1630;
	wire new_net_1517;
	wire new_net_226;
	wire _178_;
	wire _220_;
	wire _010_;
	wire _094_;
	wire new_net_40;
	wire new_net_193;
	wire new_net_699;
	wire new_net_408;
	wire new_net_1459;
	wire new_net_1636;
	wire new_net_1095;
	wire new_net_175;
	wire new_net_74;
	wire new_net_347;
	wire new_net_530;
	wire new_net_542;
	wire new_net_554;
	wire new_net_566;
	wire new_net_589;
	wire new_net_673;
	wire new_net_767;
	wire new_net_845;
	wire new_net_1364;
	wire new_net_1701;
	wire new_net_1536;
	wire new_net_1370;
	wire new_net_2028;
	wire _179_;
	wire _221_;
	wire _011_;
	wire _095_;
	wire new_net_6;
	wire new_net_57;
	wire new_net_108;
	wire new_net_606;
	wire new_net_297;
	wire new_net_572;
	wire new_net_2034;
	wire new_net_1473;
	wire new_net_1801;
	wire new_net_1222;
	wire new_net_1723;
	wire new_net_1435;
	wire new_net_1687;
	wire new_net_160;
	wire new_net_211;
	wire new_net_364;
	wire new_net_465;
	wire new_net_486;
	wire new_net_931;
	wire new_net_700;
	wire new_net_1043;
	wire new_net_1324;
	wire new_net_1518;
	wire new_net_1448;
	wire new_net_1570;
	wire new_net_1898;
	wire _012_;
	wire _096_;
	wire _180_;
	wire _222_;
	wire new_net_194;
	wire new_net_227;
	wire new_net_898;
	wire new_net_1250;
	wire new_net_1377;
	wire new_net_1389;
	wire new_net_2065;
	wire new_net_1296;
	wire new_net_1840;
	wire new_net_1783;
	wire new_net_811;
	wire new_net_24;
	wire new_net_75;
	wire new_net_279;
	wire new_net_348;
	wire new_net_789;
	wire new_net_799;
	wire new_net_1054;
	wire new_net_1179;
	wire new_net_1218;
	wire new_net_1519;
	wire new_net_1641;
	wire new_net_7;
	wire _013_;
	wire _097_;
	wire _181_;
	wire _223_;
	wire new_net_58;
	wire new_net_109;
	wire new_net_397;
	wire new_net_298;
	wire new_net_1219;
	wire new_net_1366;
	wire new_net_2024;
	wire new_net_1157;
	wire new_net_1244;
	wire new_net_41;
	wire new_net_365;
	wire new_net_455;
	wire new_net_1267;
	wire new_net_1382;
	wire new_net_1375;
	wire new_net_1460;
	wire new_net_1472;
	wire new_net_1649;
	wire new_net_1740;
	wire new_net_1912;
	wire new_net_1478;
	wire new_net_940;
	wire new_net_887;
	wire _014_;
	wire _098_;
	wire _182_;
	wire _224_;
	wire new_net_195;
	wire new_net_228;
	wire new_net_674;
	wire new_net_590;
	wire new_net_1562;
	wire new_net_1281;
	wire new_net_1279;
	wire new_net_1453;
	wire new_net_25;
	wire new_net_76;
	wire new_net_280;
	wire new_net_349;
	wire new_net_607;
	wire new_net_777;
	wire new_net_1114;
	wire new_net_1190;
	wire new_net_1413;
	wire new_net_2035;
	wire new_net_1575;
	wire new_net_1709;
	wire new_net_1869;
	wire new_net_161;
	wire new_net_932;
	wire _015_;
	wire _099_;
	wire new_net_8;
	wire _183_;
	wire _225_;
	wire new_net_59;
	wire new_net_110;
	wire new_net_701;
	wire new_net_1845;
	wire new_net_1762;
	wire new_net_1646;
	wire new_net_42;
	wire new_net_466;
	wire new_net_487;
	wire new_net_899;
	wire new_net_846;
	wire new_net_1075;
	wire new_net_1251;
	wire new_net_1262;
	wire new_net_1378;
	wire new_net_1390;
	wire new_net_778;
	wire _016_;
	wire _100_;
	wire _184_;
	wire _226_;
	wire new_net_790;
	wire new_net_800;
	wire new_net_812;
	wire new_net_1055;
	wire new_net_1180;
	wire new_net_1387;
	wire new_net_1917;
	wire new_net_26;
	wire new_net_281;
	wire new_net_299;
	wire new_net_350;
	wire new_net_405;
	wire new_net_439;
	wire new_net_597;
	wire new_net_1191;
	wire new_net_1355;
	wire new_net_1367;
	wire new_net_1485;
	wire new_net_1808;
	wire new_net_1739;
	wire new_net_1326;
	wire new_net_9;
	wire _017_;
	wire _101_;
	wire _185_;
	wire _227_;
	wire new_net_60;
	wire new_net_162;
	wire new_net_213;
	wire new_net_366;
	wire new_net_999;
	wire new_net_1254;
	wire new_net_1582;
	wire new_net_1172;
	wire new_net_1542;
	wire new_net_1714;
	wire new_net_675;
	wire new_net_532;
	wire new_net_591;
	wire new_net_769;
	wire new_net_544;
	wire new_net_43;
	wire new_net_196;
	wire new_net_229;
	wire new_net_456;
	wire new_net_556;
	wire new_net_1767;
	wire _186_;
	wire _228_;
	wire _018_;
	wire _102_;
	wire new_net_77;
	wire new_net_505;
	wire new_net_1104;
	wire new_net_1403;
	wire new_net_1414;
	wire new_net_1529;
	wire new_net_768;
	wire new_net_823;
	wire new_net_941;
	wire new_net_111;
	wire new_net_282;
	wire new_net_300;
	wire new_net_399;
	wire new_net_702;
	wire new_net_933;
	wire new_net_1105;
	wire new_net_1159;
	wire new_net_1170;
	wire new_net_1550;
	wire new_net_1135;
	wire new_net_852;
	wire new_net_1877;
	wire new_net_2007;
	wire new_net_1271;
	wire new_net_2044;
	wire new_net_888;
	wire new_net_367;
	wire new_net_900;
	wire _019_;
	wire _103_;
	wire _187_;
	wire _229_;
	wire new_net_10;
	wire new_net_163;
	wire new_net_847;
	wire new_net_1490;
	wire new_net_1813;
	wire new_net_1744;
	wire new_net_1612;
	wire new_net_779;
	wire new_net_791;
	wire new_net_801;
	wire new_net_0;
	wire new_net_197;
	wire new_net_230;
	wire new_net_425;
	wire new_net_467;
	wire new_net_488;
	wire new_net_813;
	wire new_net_1944;
	wire new_net_1788;
	wire new_net_574;
	wire new_net_1835;
	wire new_net_1259;
	wire new_net_1587;
	wire new_net_598;
	wire new_net_351;
	wire _020_;
	wire _104_;
	wire _188_;
	wire _230_;
	wire new_net_27;
	wire new_net_78;
	wire new_net_1076;
	wire new_net_1160;
	wire new_net_1313;
	wire new_net_1185;
	wire new_net_61;
	wire new_net_112;
	wire new_net_214;
	wire new_net_283;
	wire new_net_301;
	wire new_net_400;
	wire new_net_581;
	wire new_net_1000;
	wire new_net_1229;
	wire new_net_1462;
	wire new_net_870;
	wire new_net_1660;
	wire new_net_1119;
	wire new_net_1705;
	wire new_net_592;
	wire new_net_770;
	wire new_net_848;
	wire _021_;
	wire _105_;
	wire _189_;
	wire _231_;
	wire new_net_11;
	wire new_net_44;
	wire new_net_676;
	wire new_net_1671;
	wire new_net_1347;
	wire new_net_1555;
	wire new_net_1140;
	wire new_net_198;
	wire new_net_231;
	wire new_net_457;
	wire new_net_1102;
	wire new_net_1394;
	wire new_net_1415;
	wire new_net_1530;
	wire new_net_1882;
	wire new_net_1924;
	wire new_net_1994;
	wire new_net_2012;
	wire new_net_2049;
	wire new_net_1971;
	wire new_net_753;
	wire new_net_2018;
	wire new_net_1820;
	wire new_net_1940;
	wire _190_;
	wire _232_;
	wire _022_;
	wire _106_;
	wire new_net_28;
	wire new_net_79;
	wire new_net_352;
	wire new_net_411;
	wire new_net_934;
	wire new_net_703;
	wire new_net_1619;
	wire new_net_1749;
	wire new_net_1946;
	wire new_net_1126;
	wire new_net_1009;
	wire new_net_1793;
	wire new_net_901;
	wire new_net_62;
	wire new_net_113;
	wire new_net_164;
	wire new_net_215;
	wire new_net_284;
	wire new_net_368;
	wire new_net_889;
	wire new_net_1230;
	wire new_net_1253;
	wire new_net_1265;
	wire new_net_1594;
	wire new_net_1558;
	wire new_net_1523;
	wire new_net_792;
	wire new_net_802;
	wire new_net_814;
	wire _233_;
	wire _023_;
	wire _107_;
	wire _191_;
	wire new_net_12;
	wire new_net_45;
	wire new_net_780;
	wire new_net_1308;
	wire new_net_1779;
	wire new_net_722;
	wire new_net_1903;
	wire new_net_1665;
	wire new_net_232;
	wire new_net_468;
	wire new_net_489;
	wire new_net_599;
	wire new_net_1077;
	wire new_net_1161;
	wire new_net_1357;
	wire new_net_1520;
	wire new_net_1752;
	wire new_net_1972;
	wire new_net_652;
	wire new_net_582;
	wire _234_;
	wire _024_;
	wire _108_;
	wire _192_;
	wire new_net_302;
	wire new_net_1001;
	wire new_net_1463;
	wire new_net_1652;
	wire new_net_1743;
	wire new_net_1889;
	wire new_net_1399;
	wire new_net_1651;
	wire new_net_1887;
	wire new_net_1716;
	wire new_net_1936;
	wire new_net_2056;
	wire new_net_1929;
	wire new_net_2054;
	wire new_net_1976;
	wire new_net_1412;
	wire new_net_546;
	wire new_net_558;
	wire new_net_849;
	wire new_net_609;
	wire new_net_114;
	wire new_net_165;
	wire new_net_285;
	wire new_net_369;
	wire new_net_534;
	wire new_net_771;
	wire new_net_1497;
	wire new_net_1825;
	wire new_net_1624;
	wire new_net_1958;
	wire new_net_1513;
	wire new_net_1951;
	wire new_net_1753;
	wire new_net_1131;
	wire new_net_419;
	wire _025_;
	wire _109_;
	wire _193_;
	wire _235_;
	wire new_net_13;
	wire new_net_46;
	wire new_net_199;
	wire new_net_1416;
	wire new_net_1531;
	wire new_net_1360;
	wire new_net_935;
	wire new_net_704;
	wire new_net_29;
	wire new_net_80;
	wire new_net_233;
	wire new_net_353;
	wire new_net_458;
	wire new_net_1192;
	wire new_net_1328;
	wire new_net_1510;
	wire new_net_1697;
	wire new_net_1735;
	wire new_net_634;
	wire new_net_880;
	wire new_net_952;
	wire new_net_890;
	wire new_net_528;
	wire _194_;
	wire _236_;
	wire _026_;
	wire _110_;
	wire new_net_63;
	wire new_net_216;
	wire new_net_303;
	wire new_net_902;
	wire new_net_1908;
	wire new_net_1797;
	wire new_net_1719;
	wire new_net_2075;
	wire new_net_1683;
	wire new_net_2039;
	wire new_net_803;
	wire new_net_815;
	wire new_net_781;
	wire new_net_115;
	wire new_net_286;
	wire new_net_401;
	wire new_net_440;
	wire new_net_793;
	wire new_net_1046;
	wire new_net_1058;
	wire new_net_1586;
	wire new_net_1442;
	wire new_net_1566;
	wire new_net_1894;
	wire new_net_1237;
	wire new_net_1656;
	wire new_net_2061;
	wire new_net_418;
	wire new_net_600;
	wire _195_;
	wire _237_;
	wire _027_;
	wire _111_;
	wire new_net_47;
	wire new_net_200;
	wire new_net_764;
	wire new_net_1113;
	wire new_net_1502;
	wire new_net_819;
	wire new_net_1631;
	wire new_net_30;
	wire new_net_81;
	wire new_net_234;
	wire new_net_354;
	wire new_net_469;
	wire new_net_490;
	wire new_net_577;
	wire new_net_1002;
	wire new_net_1464;
	wire new_net_1653;
	wire new_net_1956;
	wire new_net_1637;
	wire new_net_296;
	wire new_net_1096;
	wire new_net_1065;
	wire new_net_573;
	wire new_net_850;
	wire new_net_610;
	wire new_net_370;
	wire new_net_772;
	wire _196_;
	wire _238_;
	wire _028_;
	wire _112_;
	wire new_net_64;
	wire new_net_1195;
	wire new_net_1027;
	wire new_net_1702;
	wire new_net_1371;
	wire new_net_2029;
	wire new_net_14;
	wire new_net_404;
	wire new_net_1106;
	wire new_net_1417;
	wire new_net_1532;
	wire new_net_212;
	wire new_net_596;
	wire new_net_1996;
	wire new_net_1474;
	wire new_net_1802;
	wire new_net_611;
	wire new_net_1223;
	wire new_net_1724;
	wire new_net_568;
	wire new_net_936;
	wire new_net_705;
	wire _239_;
	wire _029_;
	wire _113_;
	wire _197_;
	wire new_net_201;
	wire new_net_1173;
	wire new_net_1329;
	wire new_net_1688;
	wire new_net_663;
	wire new_net_242;
	wire new_net_1449;
	wire new_net_804;
	wire new_net_891;
	wire new_net_903;
	wire new_net_31;
	wire new_net_235;
	wire new_net_304;
	wire new_net_355;
	wire new_net_459;
	wire new_net_1116;
	wire new_net_1124;
	wire new_net_1232;
	wire new_net_1899;
	wire new_net_2066;
	wire new_net_1750;
	wire new_net_1774;
	wire new_net_1297;
	wire new_net_1422;
	wire _030_;
	wire _114_;
	wire _198_;
	wire _240_;
	wire new_net_116;
	wire new_net_167;
	wire new_net_677;
	wire new_net_782;
	wire new_net_287;
	wire new_net_794;
	wire new_net_1758;
	wire new_net_1319;
	wire new_net_1642;
	wire new_net_1101;
	wire new_net_15;
	wire new_net_48;
	wire new_net_601;
	wire new_net_1163;
	wire new_net_1194;
	wire new_net_1359;
	wire new_net_1522;
	wire new_net_1754;
	wire new_net_1974;
	wire new_net_2025;
	wire _031_;
	wire _115_;
	wire _199_;
	wire _241_;
	wire new_net_82;
	wire new_net_569;
	wire new_net_1003;
	wire new_net_1465;
	wire new_net_1654;
	wire new_net_1745;
	wire new_net_1383;
	wire new_net_1913;
	wire new_net_65;
	wire new_net_218;
	wire new_net_236;
	wire new_net_305;
	wire new_net_470;
	wire new_net_491;
	wire new_net_678;
	wire new_net_536;
	wire new_net_773;
	wire new_net_548;
	wire new_net_1479;
	wire new_net_1228;
	wire new_net_1729;
	wire new_net_1603;
	wire new_net_1693;
	wire new_net_1454;
	wire new_net_288;
	wire _032_;
	wire _116_;
	wire _200_;
	wire _242_;
	wire new_net_117;
	wire new_net_168;
	wire new_net_1107;
	wire new_net_1418;
	wire new_net_1997;
	wire new_net_1578;
	wire new_net_1576;
	wire new_net_1870;
	wire new_net_49;
	wire new_net_202;
	wire new_net_706;
	wire new_net_937;
	wire new_net_1084;
	wire new_net_1174;
	wire new_net_1330;
	wire new_net_1049;
	wire new_net_1512;
	wire new_net_1854;
	wire new_net_1763;
	wire new_net_1850;
	wire new_net_863;
	wire _007_;
	wire _033_;
	wire _117_;
	wire _201_;
	wire _243_;
	wire new_net_32;
	wire new_net_83;
	wire new_net_356;
	wire new_net_892;
	wire new_net_583;
	wire new_net_904;
	wire new_net_66;
	wire new_net_219;
	wire new_net_372;
	wire new_net_460;
	wire new_net_783;
	wire new_net_795;
	wire new_net_805;
	wire new_net_1048;
	wire new_net_1098;
	wire new_net_1117;
	wire new_net_1546;
	wire new_net_2003;
	wire new_net_1918;
	wire new_net_429;
	wire new_net_16;
	wire _202_;
	wire _244_;
	wire _034_;
	wire _118_;
	wire new_net_118;
	wire new_net_169;
	wire new_net_602;
	wire new_net_1164;
	wire new_net_1486;
	wire new_net_1809;
	wire new_net_1327;
	wire new_net_50;
	wire new_net_203;
	wire new_net_449;
	wire new_net_570;
	wire new_net_1004;
	wire new_net_1079;
	wire new_net_1466;
	wire new_net_1533;
	wire new_net_1655;
	wire new_net_1746;
	wire new_net_1784;
	wire new_net_1831;
	wire new_net_1255;
	wire new_net_1583;
	wire new_net_584;
	wire new_net_774;
	wire _035_;
	wire _119_;
	wire _203_;
	wire _245_;
	wire new_net_33;
	wire new_net_84;
	wire new_net_237;
	wire new_net_306;
	wire new_net_1715;
	wire new_net_1309;
	wire new_net_1056;
	wire new_net_1181;
	wire new_net_1770;
	wire new_net_1768;
	wire new_net_289;
	wire new_net_373;
	wire new_net_471;
	wire new_net_492;
	wire new_net_1059;
	wire new_net_1108;
	wire new_net_1419;
	wire new_net_1596;
	wire new_net_1855;
	wire new_net_1998;
	wire new_net_938;
	wire new_net_707;
	wire new_net_17;
	wire _036_;
	wire _120_;
	wire _204_;
	wire _246_;
	wire new_net_575;
	wire new_net_1175;
	wire new_net_1331;
	wire new_net_1551;
	wire new_net_1136;
	wire new_net_1878;
	wire new_net_2008;
	wire new_net_204;
	wire new_net_576;
	wire new_net_816;
	wire new_net_851;
	wire new_net_893;
	wire new_net_905;
	wire new_net_1234;
	wire new_net_1257;
	wire new_net_1272;
	wire new_net_1372;
	wire new_net_2045;
	wire new_net_2043;
	wire new_net_2014;
	wire new_net_1491;
	wire new_net_1814;
	wire new_net_1615;
	wire new_net_784;
	wire new_net_358;
	wire _037_;
	wire _121_;
	wire _205_;
	wire _247_;
	wire new_net_67;
	wire new_net_238;
	wire new_net_307;
	wire new_net_806;
	wire new_net_1537;
	wire new_net_1592;
	wire new_net_1789;
	wire new_net_1044;
	wire new_net_1590;
	wire new_net_119;
	wire new_net_170;
	wire new_net_290;
	wire new_net_374;
	wire new_net_461;
	wire new_net_603;
	wire new_net_1165;
	wire new_net_1196;
	wire new_net_1260;
	wire new_net_1361;
	wire new_net_1588;
	wire new_net_1316;
	wire new_net_1599;
	wire new_net_1060;
	wire new_net_1186;
	wire _206_;
	wire _248_;
	wire _038_;
	wire _122_;
	wire new_net_18;
	wire new_net_51;
	wire new_net_1005;
	wire new_net_1080;
	wire new_net_1467;
	wire new_net_1534;
	wire new_net_1775;
	wire new_net_381;
	wire new_net_876;
	wire new_net_1153;
	wire new_net_1661;
	wire new_net_1120;
	wire new_net_680;
	wire new_net_775;
	wire new_net_817;
	wire new_net_34;
	wire new_net_85;
	wire new_net_205;
	wire new_net_538;
	wire new_net_550;
	wire new_net_562;
	wire new_net_585;
	wire new_net_1991;
	wire new_net_1672;
	wire new_net_969;
	wire new_net_973;
	wire new_net_1348;
	wire _207_;
	wire _249_;
	wire _039_;
	wire _123_;
	wire new_net_68;
	wire new_net_221;
	wire new_net_359;
	wire new_net_308;
	wire new_net_1109;
	wire new_net_1420;
	wire new_net_1395;
	wire new_net_1883;
	wire new_net_1925;
	wire new_net_2013;
	wire new_net_2050;
	wire new_net_1199;
	wire new_net_1821;
	wire new_net_708;
	wire new_net_120;
	wire new_net_171;
	wire new_net_430;
	wire new_net_472;
	wire new_net_493;
	wire new_net_1176;
	wire new_net_1332;
	wire new_net_1514;
	wire new_net_1703;
	wire new_net_1941;
	wire new_net_1509;
	wire new_net_1947;
	wire new_net_1127;
	wire new_net_594;
	wire new_net_894;
	wire _208_;
	wire _250_;
	wire new_net_1;
	wire _040_;
	wire _124_;
	wire new_net_52;
	wire new_net_906;
	wire new_net_1235;
	wire new_net_1266;
	wire new_net_1595;
	wire new_net_1144;
	wire new_net_1356;
	wire new_net_1524;
	wire new_net_807;
	wire new_net_35;
	wire new_net_86;
	wire new_net_206;
	wire new_net_239;
	wire new_net_446;
	wire new_net_785;
	wire new_net_1050;
	wire new_net_1061;
	wire new_net_1100;
	wire new_net_1323;
	wire new_net_1780;
	wire new_net_524;
	wire new_net_1904;
	wire new_net_604;
	wire _041_;
	wire _125_;
	wire _209_;
	wire _251_;
	wire new_net_69;
	wire new_net_222;
	wire new_net_291;
	wire new_net_375;
	wire new_net_1166;
	wire new_net_1666;
	wire new_net_1677;
	wire new_net_19;
	wire new_net_121;
	wire new_net_172;
	wire new_net_462;
	wire new_net_942;
	wire new_net_1081;
	wire new_net_1468;
	wire new_net_1535;
	wire new_net_1657;
	wire new_net_1748;
	wire new_net_1890;
	wire new_net_1233;
	wire new_net_1888;
	wire new_net_1937;
	wire new_net_2057;
	wire new_net_1930;
	wire new_net_2055;
	wire new_net_776;
	wire new_net_818;
	wire new_net_853;
	wire new_net_614;
	wire _210_;
	wire _252_;
	wire _042_;
	wire _126_;
	wire new_net_2;
	wire new_net_586;
	wire new_net_1861;
	wire new_net_1977;
	wire new_net_1498;
	wire new_net_1826;
	wire new_net_1627;
	wire new_net_1171;
	wire new_net_1959;
	wire new_net_87;
	wire new_net_207;
	wire new_net_240;
	wire new_net_309;
	wire new_net_360;
	wire new_net_1110;
	wire new_net_1421;
	wire new_net_1598;
	wire new_net_1756;
	wire new_net_1847;
	wire new_net_1874;
	wire new_net_1999;
	wire _211_;
	wire _253_;
	wire _043_;
	wire _127_;
	wire new_net_292;
	wire new_net_376;
	wire new_net_709;
	wire new_net_1177;
	wire new_net_1333;
	wire new_net_1515;
	wire new_net_1111;
	wire new_net_1698;
	wire new_net_1736;
	wire new_net_1115;
	wire new_net_907;
	wire new_net_595;
	wire new_net_881;
	wire new_net_473;
	wire new_net_20;
	wire new_net_53;
	wire new_net_122;
	wire new_net_173;
	wire new_net_494;
	wire new_net_895;
	wire new_net_1909;
	wire new_net_1798;
	wire new_net_1720;
	wire new_net_2076;
	wire new_net_1684;
	wire new_net_2040;
	wire new_net_433;
	wire new_net_808;
	wire _212_;
	wire _254_;
	wire _044_;
	wire _128_;
	wire new_net_36;
	wire new_net_786;
	wire new_net_1051;
	wire new_net_1062;
	wire new_net_1443;
	wire new_net_1567;
	wire new_net_1895;
	wire new_net_70;
	wire new_net_223;
	wire new_net_310;
	wire new_net_361;
	wire new_net_1167;
	wire new_net_1363;
	wire new_net_1526;
	wire new_net_1837;
	wire new_net_1978;
	wire new_net_2062;
	wire new_net_1503;
	wire new_net_939;
	wire _213_;
	wire _255_;
	wire _045_;
	wire _129_;
	wire new_net_293;
	wire new_net_377;
	wire new_net_1082;
	wire new_net_1469;
	wire new_net_1658;
	wire new_net_1638;
	wire new_net_1846;
	wire new_net_1664;
	wire new_net_1097;
	wire new_net_1268;
	wire new_net_564;
	wire new_net_854;
	wire new_net_552;
	wire new_net_615;
	wire new_net_587;
	wire new_net_3;
	wire new_net_21;
	wire new_net_54;
	wire new_net_445;
	wire new_net_463;
	wire new_net_625;
	wire new_net_241;
	wire new_net_796;
	wire new_net_953;
	wire new_net_407;
	wire _214_;
	wire _256_;
	wire _046_;
	wire _130_;
	wire new_net_37;
	wire new_net_88;
	wire new_net_1379;
	wire new_net_2030;
	wire new_net_2036;
	wire new_net_1475;
	wire new_net_1803;
	wire new_net_71;
	wire new_net_224;
	wire new_net_311;
	wire new_net_441;
	wire new_net_612;
	wire new_net_710;
	wire new_net_1006;
	wire new_net_1178;
	wire new_net_1224;
	wire new_net_1334;
	wire new_net_1725;
	wire new_net_1689;
	wire new_net_664;
	wire new_net_985;
	wire new_net_294;
	wire new_net_896;
	wire _047_;
	wire _131_;
	wire _215_;
	wire _257_;
	wire new_net_123;
	wire new_net_174;
	wire new_net_908;
	wire new_net_378;
	wire new_net_1572;
	wire new_net_1900;
	wire new_net_1706;
	wire new_net_2067;
	wire new_net_1045;
	wire new_net_809;
	wire new_net_943;
	wire new_net_787;
	wire new_net_4;
	wire new_net_55;
	wire new_net_406;
	wire new_net_474;
	wire new_net_495;
	wire new_net_797;
	wire new_net_1052;
	wire new_net_1261;
	wire new_net_1842;
	wire new_net_1759;
	wire new_net_1556;
	wire new_net_1320;
	wire new_net_209;
	wire new_net_428;
	wire new_net_362;
	wire new_net_448;
	wire _048_;
	wire _132_;
	wire _216_;
	wire _258_;
	wire new_net_38;
	wire new_net_89;
	wire new_net_1368;
	wire new_net_257;
	wire new_net_72;
	wire new_net_225;
	wire new_net_312;
	wire new_net_437;
	wire new_net_681;
	wire new_net_1007;
	wire new_net_1083;
	wire new_net_1470;
	wire new_net_1659;
	wire new_net_1757;
	wire new_net_1384;
	wire new_net_1471;
	wire new_net_1914;
	wire new_net_1906;
	wire new_net_295;
	wire new_net_616;
	wire new_net_588;
	wire new_net_820;
	wire _049_;
	wire _133_;
	wire _217_;
	wire _259_;
	wire new_net_22;
	wire new_net_124;
	wire new_net_1482;
	wire new_net_1805;
	wire new_net_1480;
	wire new_net_1694;
	wire new_net_669;
	wire new_net_5;
	wire new_net_464;
	wire new_net_1112;
	wire new_net_1141;
	wire new_net_1423;
	wire new_net_1600;
	wire new_net_2002;
	wire new_net_2033;
	wire new_net_1455;
	wire new_net_1579;
	wire new_net_1078;
	wire new_net_1577;
	wire new_net_1711;
	wire new_net_402;
	wire new_net_363;
	wire new_net_243;
	wire new_net_711;
	wire new_net_682;
	wire _218_;
	wire _260_;
	wire _050_;
	wire _134_;
	wire new_net_39;
	wire new_net_1836;
	wire new_net_1764;
	wire new_net_1851;
	wire new_net_864;
	wire new_net_73;
	wire new_net_379;
	wire new_net_897;
	wire new_net_909;
	wire new_net_1168;
	wire new_net_1198;
	wire new_net_1238;
	wire new_net_1376;
	wire new_net_1388;
	wire new_net_1400;
	wire new_net_1563;
	wire new_net_1130;
	wire new_net_1547;
	wire new_net_1860;
	wire new_net_1132;
	wire new_net_1042;
	wire new_net_1342;
	wire _051_;
	wire _135_;
	wire _261_;
	wire new_net_944;
	wire new_net_734;
	wire new_net_866;
	wire new_net_1064;
	wire new_net_1122;
	wire new_net_1142;
	wire new_net_1269;
	wire new_net_1487;
	wire new_net_1810;
	wire new_net_1741;
	wire new_net_1609;
	wire new_net_2019;
	wire new_net_1952;
	wire new_net_475;
	wire new_net_496;
	wire new_net_517;
	wire new_net_1032;
	wire new_net_1980;
	wire new_net_1785;
	wire new_net_997;
	wire new_net_1832;
	wire new_net_1865;
	wire new_net_1256;
	wire new_net_1584;
	wire _052_;
	wire _262_;
	wire _136_;
	wire new_net_142;
	wire new_net_313;
	wire new_net_331;
	wire new_net_966;
	wire new_net_977;
	wire new_net_989;
	wire new_net_1008;
	wire new_net_1057;
	wire new_net_1182;
	wire new_net_1771;
	wire new_net_1769;
	wire new_net_1856;
	wire new_net_650;
	wire new_net_691;
	wire new_net_856;
	wire new_net_125;
	wire new_net_176;
	wire new_net_380;
	wire new_net_617;
	wire new_net_862;
	wire new_net_756;
	wire new_net_872;
	wire _263_;
	wire _053_;
	wire _137_;
	wire new_net_261;
	wire new_net_1014;
	wire new_net_1424;
	wire new_net_1436;
	wire new_net_1601;
	wire new_net_1613;
	wire new_net_1625;
	wire new_net_1227;
	wire new_net_1552;
	wire new_net_1873;
	wire new_net_1137;
	wire new_net_1391;
	wire new_net_1879;
	wire new_net_2009;
	wire new_net_2046;
	wire new_net_683;
	wire new_net_91;
	wire new_net_244;
	wire new_net_507;
	wire new_net_832;
	wire new_net_712;
	wire new_net_1336;
	wire new_net_1343;
	wire new_net_1858;
	wire new_net_1867;
	wire new_net_2015;
	wire new_net_1817;
	wire new_net_1246;
	wire new_net_1492;
	wire new_net_1815;
	wire _264_;
	wire _054_;
	wire _138_;
	wire new_net_314;
	wire new_net_910;
	wire new_net_1209;
	wire new_net_1239;
	wire new_net_1291;
	wire new_net_1303;
	wire new_net_1315;
	wire new_net_1284;
	wire new_net_1790;
	wire new_net_1591;
	wire new_net_1589;
	wire new_net_945;
	wire new_net_126;
	wire new_net_177;
	wire new_net_723;
	wire new_net_735;
	wire new_net_922;
	wire new_net_1123;
	wire new_net_1143;
	wire new_net_1270;
	wire new_net_1538;
	wire new_net_1187;
	wire _265_;
	wire _139_;
	wire _055_;
	wire new_net_262;
	wire new_net_442;
	wire new_net_1033;
	wire new_net_1776;
	wire new_net_1981;
	wire new_net_1662;
	wire new_net_1829;
	wire new_net_1121;
	wire new_net_593;
	wire new_net_92;
	wire new_net_143;
	wire new_net_245;
	wire new_net_332;
	wire new_net_476;
	wire new_net_497;
	wire new_net_518;
	wire new_net_967;
	wire new_net_978;
	wire new_net_990;
	wire new_net_1673;
	wire new_net_745;
	wire new_net_618;
	wire new_net_662;
	wire new_net_822;
	wire _056_;
	wire _266_;
	wire _140_;
	wire new_net_315;
	wire new_net_757;
	wire new_net_873;
	wire new_net_1396;
	wire new_net_1648;
	wire new_net_1884;
	wire new_net_1926;
	wire new_net_2051;
	wire new_net_1973;
	wire new_net_1200;
	wire new_net_1494;
	wire new_net_1822;
	wire new_net_178;
	wire new_net_923;
	wire new_net_1425;
	wire new_net_1437;
	wire new_net_1602;
	wire new_net_1614;
	wire new_net_1626;
	wire new_net_2004;
	wire new_net_1621;
	wire new_net_1948;
	wire new_net_1128;
	wire new_net_1214;
	wire new_net_1995;
	wire new_net_833;
	wire _267_;
	wire _057_;
	wire _141_;
	wire new_net_713;
	wire new_net_263;
	wire new_net_1344;
	wire new_net_2069;
	wire new_net_1145;
	wire new_net_1730;
	wire new_net_1560;
	wire new_net_1525;
	wire new_net_93;
	wire new_net_144;
	wire new_net_333;
	wire new_net_443;
	wire new_net_508;
	wire new_net_911;
	wire new_net_1210;
	wire new_net_1240;
	wire new_net_1292;
	wire new_net_1304;
	wire new_net_1781;
	wire new_net_1905;
	wire new_net_1247;
	wire new_net_1794;
	wire new_net_1667;
	wire new_net_724;
	wire new_net_736;
	wire _058_;
	wire _142_;
	wire _268_;
	wire new_net_127;
	wire new_net_316;
	wire new_net_382;
	wire new_net_946;
	wire new_net_1085;
	wire new_net_2072;
	wire new_net_1034;
	wire new_net_1439;
	wire new_net_1982;
	wire new_net_1891;
	wire new_net_2058;
	wire new_net_956;
	wire _143_;
	wire _059_;
	wire _269_;
	wire new_net_409;
	wire new_net_246;
	wire new_net_968;
	wire new_net_979;
	wire new_net_991;
	wire new_net_1010;
	wire new_net_1499;
	wire new_net_1506;
	wire new_net_1827;
	wire new_net_1862;
	wire new_net_1960;
	wire new_net_1953;
	wire new_net_1755;
	wire new_net_758;
	wire new_net_519;
	wire new_net_630;
	wire new_net_94;
	wire new_net_145;
	wire new_net_334;
	wire new_net_477;
	wire new_net_498;
	wire new_net_882;
	wire new_net_641;
	wire new_net_1875;
	wire new_net_1955;
	wire new_net_2000;
	wire new_net_383;
	wire _144_;
	wire _060_;
	wire _270_;
	wire new_net_128;
	wire new_net_179;
	wire new_net_924;
	wire new_net_692;
	wire new_net_1362;
	wire new_net_1426;
	wire new_net_1699;
	wire new_net_1737;
	wire new_net_2026;
	wire new_net_264;
	wire new_net_714;
	wire new_net_834;
	wire new_net_1073;
	wire new_net_1345;
	wire new_net_2070;
	wire new_net_1799;
	wire new_net_1220;
	wire new_net_1721;
	wire new_net_2077;
	wire new_net_1685;
	wire new_net_2041;
	wire new_net_912;
	wire _061_;
	wire _145_;
	wire _271_;
	wire new_net_247;
	wire new_net_410;
	wire new_net_1211;
	wire new_net_1241;
	wire new_net_1293;
	wire new_net_1305;
	wire new_net_1568;
	wire new_net_1896;
	wire new_net_737;
	wire new_net_693;
	wire new_net_509;
	wire new_net_95;
	wire new_net_146;
	wire new_net_317;
	wire new_net_421;
	wire new_net_947;
	wire new_net_725;
	wire new_net_970;
	wire new_net_1162;
	wire new_net_2063;
	wire new_net_1504;
	wire new_net_423;
	wire new_net_180;
	wire new_net_436;
	wire _062_;
	wire _146_;
	wire _272_;
	wire new_net_129;
	wire new_net_1035;
	wire new_net_1066;
	wire new_net_1282;
	wire new_net_1639;
	wire new_net_1287;
	wire new_net_1733;
	wire new_net_957;
	wire new_net_265;
	wire new_net_684;
	wire new_net_980;
	wire new_net_992;
	wire new_net_1011;
	wire new_net_1202;
	wire new_net_628;
	wire new_net_1438;
	wire new_net_1450;
	wire new_net_1197;
	wire new_net_1380;
	wire new_net_580;
	wire new_net_631;
	wire new_net_824;
	wire new_net_653;
	wire _063_;
	wire _147_;
	wire _273_;
	wire new_net_335;
	wire new_net_747;
	wire new_net_620;
	wire new_net_1910;
	wire new_net_1476;
	wire new_net_1804;
	wire new_net_613;
	wire new_net_1225;
	wire new_net_1726;
	wire new_net_318;
	wire new_net_384;
	wire new_net_478;
	wire new_net_499;
	wire new_net_925;
	wire new_net_1427;
	wire new_net_1604;
	wire new_net_1616;
	wire new_net_1628;
	wire new_net_2006;
	wire new_net_1690;
	wire new_net_1451;
	wire new_net_715;
	wire _064_;
	wire _148_;
	wire _274_;
	wire new_net_130;
	wire new_net_835;
	wire new_net_181;
	wire new_net_1346;
	wire new_net_1573;
	wire new_net_2071;
	wire new_net_403;
	wire new_net_1707;
	wire new_net_1992;
	wire new_net_1299;
	wire new_net_913;
	wire new_net_248;
	wire new_net_266;
	wire new_net_874;
	wire new_net_1016;
	wire new_net_1212;
	wire new_net_1242;
	wire new_net_1294;
	wire new_net_1306;
	wire new_net_1404;
	wire new_net_1843;
	wire new_net_1094;
	wire new_net_1760;
	wire new_net_1015;
	wire new_net_1644;
	wire new_net_694;
	wire new_net_948;
	wire new_net_147;
	wire new_net_336;
	wire new_net_726;
	wire _275_;
	wire _065_;
	wire _149_;
	wire new_net_96;
	wire new_net_738;
	wire new_net_319;
	wire new_net_385;
	wire new_net_510;
	wire new_net_1036;
	wire new_net_1067;
	wire new_net_1984;
	wire new_net_1385;
	wire new_net_1915;
	wire new_net_1483;
	wire new_net_1806;
	wire new_net_958;
	wire _276_;
	wire _066_;
	wire _150_;
	wire new_net_182;
	wire new_net_981;
	wire new_net_993;
	wire new_net_1025;
	wire new_net_1203;
	wire new_net_1317;
	wire new_net_1481;
	wire new_net_670;
	wire new_net_654;
	wire new_net_665;
	wire new_net_825;
	wire new_net_748;
	wire new_net_249;
	wire new_net_267;
	wire new_net_522;
	wire new_net_632;
	wire new_net_1559;
	wire new_net_1710;
	wire new_net_1252;
	wire new_net_1580;
	wire new_net_1208;
	wire new_net_1712;
	wire new_net_148;
	wire new_net_337;
	wire new_net_926;
	wire _067_;
	wire _277_;
	wire _151_;
	wire new_net_97;
	wire new_net_1053;
	wire new_net_1428;
	wire new_net_1605;
	wire new_net_1765;
	wire new_net_1852;
	wire new_net_865;
	wire new_net_1401;
	wire new_net_836;
	wire new_net_500;
	wire new_net_131;
	wire new_net_320;
	wire new_net_386;
	wire new_net_417;
	wire new_net_479;
	wire new_net_716;
	wire new_net_1146;
	wire new_net_1273;
	wire new_net_1564;
	wire new_net_1983;
	wire new_net_998;
	wire new_net_639;
	wire new_net_821;
	wire new_net_914;
	wire new_net_857;
	wire _068_;
	wire _278_;
	wire _152_;
	wire new_net_183;
	wire new_net_1017;
	wire new_net_1026;
	wire new_net_1213;
	wire new_net_1243;
	wire new_net_1548;
	wire new_net_1133;
	wire new_net_2005;
	wire new_net_746;
	wire new_net_1920;
	wire new_net_949;
	wire new_net_727;
	wire new_net_739;
	wire new_net_695;
	wire new_net_250;
	wire new_net_268;
	wire new_net_432;
	wire new_net_642;
	wire new_net_1086;
	wire new_net_1676;
	wire new_net_1488;
	wire new_net_1811;
	wire new_net_1742;
	wire new_net_2020;
	wire new_net_413;
	wire _279_;
	wire _069_;
	wire _153_;
	wire new_net_98;
	wire new_net_1037;
	wire new_net_1068;
	wire new_net_1125;
	wire new_net_1961;
	wire new_net_1985;
	wire new_net_1786;
	wire new_net_1833;
	wire new_net_1866;
	wire new_net_540;
	wire new_net_1585;
	wire new_net_579;
	wire new_net_685;
	wire new_net_959;
	wire new_net_132;
	wire new_net_321;
	wire new_net_511;
	wire new_net_982;
	wire new_net_994;
	wire new_net_1204;
	wire new_net_1318;
	wire new_net_1717;
	wire new_net_1311;
	wire new_net_571;
	wire new_net_1183;
	wire new_net_1772;
	wire new_net_655;
	wire new_net_858;
	wire new_net_749;
	wire new_net_666;
	wire new_net_633;
	wire _280_;
	wire _070_;
	wire _154_;
	wire new_net_643;
	wire new_net_826;
	wire new_net_1857;
	wire new_net_927;
	wire new_net_149;
	wire new_net_251;
	wire new_net_269;
	wire new_net_338;
	wire new_net_450;
	wire new_net_1087;
	wire new_net_730;
	wire new_net_1405;
	wire new_net_1429;
	wire new_net_90;
	wire new_net_608;
	wire new_net_1553;
	wire new_net_1138;
	wire new_net_855;
	wire new_net_1392;
	wire new_net_1880;
	wire new_net_1897;
	wire new_net_686;
	wire new_net_837;
	wire new_net_843;
	wire new_net_717;
	wire _281_;
	wire _155_;
	wire _071_;
	wire new_net_99;
	wire new_net_387;
	wire new_net_1274;
	wire new_net_1922;
	wire new_net_2010;
	wire new_net_2047;
	wire new_net_1969;
	wire new_net_751;
	wire new_net_2016;
	wire new_net_1818;
	wire new_net_371;
	wire new_net_1938;
	wire new_net_1493;
	wire new_net_1816;
	wire new_net_480;
	wire new_net_501;
	wire new_net_875;
	wire new_net_915;
	wire new_net_133;
	wire new_net_184;
	wire new_net_322;
	wire new_net_435;
	wire new_net_986;
	wire new_net_1018;
	wire new_net_1539;
	wire new_net_1617;
	wire new_net_1747;
	wire new_net_1791;
	wire _072_;
	wire _282_;
	wire _156_;
	wire new_net_760;
	wire new_net_728;
	wire new_net_883;
	wire new_net_696;
	wire new_net_740;
	wire new_net_950;
	wire new_net_621;
	wire new_net_1263;
	wire new_net_1521;
	wire _091_;
	wire new_net_1188;
	wire new_net_150;
	wire new_net_252;
	wire new_net_339;
	wire new_net_427;
	wire new_net_1069;
	wire new_net_1962;
	wire new_net_1986;
	wire new_net_1777;
	wire new_net_1901;
	wire new_net_1663;
	wire new_net_2068;
	wire _283_;
	wire _073_;
	wire _157_;
	wire new_net_388;
	wire new_net_867;
	wire new_net_960;
	wire new_net_971;
	wire new_net_983;
	wire new_net_995;
	wire new_net_1205;
	wire new_net_2031;
	wire new_net_1674;
	wire new_net_656;
	wire new_net_859;
	wire new_net_134;
	wire new_net_185;
	wire new_net_323;
	wire new_net_512;
	wire new_net_750;
	wire new_net_622;
	wire new_net_667;
	wire new_net_761;
	wire new_net_1350;
	wire new_net_1397;
	wire new_net_1885;
	wire new_net_1934;
	wire new_net_1927;
	wire new_net_2052;
	wire new_net_1283;
	wire new_net_1201;
	wire new_net_1495;
	wire _284_;
	wire _074_;
	wire _158_;
	wire new_net_270;
	wire new_net_424;
	wire new_net_1088;
	wire new_net_1406;
	wire new_net_1430;
	wire new_net_1540;
	wire new_net_1607;
	wire new_net_1823;
	wire new_net_1511;
	wire new_net_1949;
	wire new_net_1751;
	wire new_net_1129;
	wire new_net_1871;
	wire new_net_100;
	wire new_net_151;
	wire new_net_253;
	wire new_net_687;
	wire new_net_718;
	wire new_net_838;
	wire new_net_1147;
	wire new_net_1275;
	wire new_net_1337;
	wire new_net_1349;
	wire new_net_166;
	wire new_net_1731;
	wire new_net_1561;
	wire new_net_1358;
	wire _285_;
	wire _159_;
	wire _075_;
	wire new_net_447;
	wire new_net_916;
	wire new_net_1019;
	wire new_net_1028;
	wire new_net_1154;
	wire new_net_1215;
	wire new_net_1285;
	wire new_net_1695;
	wire new_net_1704;
	wire new_net_729;
	wire new_net_135;
	wire new_net_186;
	wire new_net_324;
	wire new_net_481;
	wire new_net_502;
	wire new_net_697;
	wire new_net_741;
	wire new_net_951;
	wire new_net_1678;
	wire new_net_1668;
	wire new_net_1795;
	wire new_net_2073;
	wire new_net_2037;
	wire new_net_1679;
	wire _160_;
	wire _076_;
	wire _286_;
	wire new_net_271;
	wire new_net_340;
	wire new_net_1070;
	wire new_net_1148;
	wire new_net_1963;
	wire new_net_1987;
	wire new_net_1440;
	wire new_net_1571;
	wire new_net_1892;
	wire new_net_2059;
	wire new_net_1932;
	wire new_net_101;
	wire new_net_254;
	wire new_net_389;
	wire new_net_868;
	wire new_net_961;
	wire new_net_884;
	wire new_net_972;
	wire new_net_984;
	wire new_net_996;
	wire new_net_1206;
	wire new_net_1288;
	wire new_net_1979;
	wire new_net_1507;
	wire new_net_1863;
	wire new_net_1500;
	wire new_net_1828;
	wire new_net_1629;
	wire new_net_762;
	wire new_net_877;
	wire _077_;
	wire _161_;
	wire new_net_860;
	wire new_net_645;
	wire new_net_828;
	wire new_net_623;
	wire new_net_668;
	wire new_net_657;
	wire new_net_1189;
	wire new_net_1516;
	wire new_net_1954;
	wire new_net_1876;
	wire new_net_2001;
	wire new_net_1354;
	wire new_net_438;
	wire new_net_513;
	wire new_net_1089;
	wire new_net_1407;
	wire new_net_1431;
	wire new_net_1541;
	wire new_net_1608;
	wire new_net_1620;
	wire new_net_1632;
	wire new_net_1193;
	wire new_net_1700;
	wire new_net_1841;
	wire new_net_1738;
	wire new_net_679;
	wire new_net_1369;
	wire new_net_2027;
	wire new_net_1461;
	wire new_net_839;
	wire _078_;
	wire _162_;
	wire new_net_152;
	wire new_net_272;
	wire new_net_341;
	wire new_net_719;
	wire new_net_688;
	wire new_net_1276;
	wire new_net_1338;
	wire new_net_1800;
	wire new_net_1221;
	wire new_net_1722;
	wire new_net_390;
	wire new_net_917;
	wire new_net_1020;
	wire new_net_1029;
	wire new_net_1155;
	wire new_net_1216;
	wire new_net_1245;
	wire new_net_1286;
	wire new_net_1298;
	wire new_net_1310;
	wire new_net_1686;
	wire new_net_2042;
	wire new_net_1447;
	wire new_net_1569;
	wire new_net_742;
	wire new_net_431;
	wire new_net_698;
	wire _079_;
	wire _163_;
	wire new_net_136;
	wire new_net_187;
	wire new_net_414;
	wire new_net_325;
	wire new_net_578;
	wire new_net_2064;
	wire new_net_1295;
	wire new_net_1505;
	wire new_net_451;
	wire new_net_482;
	wire new_net_503;
	wire new_net_1038;
	wire new_net_1071;
	wire new_net_1149;
	wire new_net_1964;
	wire new_net_1988;
	wire new_net_1640;
	wire new_net_1848;
	wire new_net_1099;
	wire new_net_273;
	wire new_net_342;
	wire new_net_885;
	wire new_net_962;
	wire _080_;
	wire _164_;
	wire new_net_102;
	wire new_net_153;
	wire new_net_434;
	wire new_net_255;
	wire new_net_629;
	wire new_net_2023;
	wire new_net_763;
	wire new_net_878;
	wire new_net_635;
	wire new_net_391;
	wire new_net_526;
	wire new_net_646;
	wire new_net_829;
	wire new_net_658;
	wire new_net_752;
	wire new_net_624;
	wire new_net_1374;
	wire new_net_1381;
	wire new_net_1911;
	wire new_net_1477;
	wire new_net_326;
	wire _081_;
	wire _165_;
	wire new_net_137;
	wire new_net_188;
	wire new_net_426;
	wire new_net_1090;
	wire new_net_1226;
	wire new_net_1408;
	wire new_net_1432;
	wire new_net_1727;
	wire new_net_1280;
	wire new_net_1691;
	wire new_net_1278;
	wire new_net_1452;
	wire new_net_720;
	wire new_net_416;
	wire new_net_514;
	wire new_net_689;
	wire new_net_840;
	wire new_net_1039;
	wire new_net_1277;
	wire new_net_1339;
	wire new_net_1351;
	wire new_net_1942;
	wire new_net_1574;
	wire new_net_1708;
	wire new_net_1868;
	wire new_net_1993;
	wire new_net_1169;
	wire new_net_1300;
	wire new_net_918;
	wire _082_;
	wire _166_;
	wire new_net_103;
	wire new_net_154;
	wire new_net_256;
	wire new_net_1021;
	wire new_net_1030;
	wire new_net_1047;
	wire new_net_1156;
	wire new_net_1844;
	wire new_net_1761;
	wire new_net_743;
	wire new_net_731;
	wire new_net_1207;
	wire new_net_1321;
	wire new_net_1645;
	wire new_net_1680;
	wire new_net_1692;
	wire new_net_1919;
	wire new_net_1931;
	wire new_net_2022;
	wire _167_;
	wire _083_;
	wire new_net_327;
	wire new_net_1012;
	wire new_net_1072;
	wire new_net_1150;
	wire new_net_1965;
	wire new_net_1989;
	wire new_net_1386;
	wire new_net_1916;
	wire new_net_963;
	wire new_net_274;
	wire new_net_343;
	wire new_net_483;
	wire new_net_504;
	wire new_net_974;
	wire new_net_1444;
	wire new_net_1456;
	wire new_net_1484;
	wire new_net_1633;
	wire new_net_1807;
	wire new_net_1373;
	wire new_net_1606;
	wire new_net_1325;
	wire new_net_392;
	wire new_net_636;
	wire new_net_647;
	wire new_net_928;
	wire new_net_520;
	wire new_net_659;
	wire _168_;
	wire _000_;
	wire _084_;
	wire new_net_155;
	wire new_net_1782;
	wire new_net_1457;
	wire new_net_1581;
	wire new_net_1643;
	wire new_net_138;
	wire new_net_189;
	wire new_net_1091;
	wire new_net_1217;
	wire new_net_1409;
	wire new_net_1433;
	wire new_net_1307;
	wire new_net_1543;
	wire new_net_1610;
	wire new_net_1622;
	wire new_net_1713;
	wire new_net_1838;
	wire new_net_1766;
	wire new_net_1853;
	wire new_net_721;
	wire new_net_690;
	wire _001_;
	wire _085_;
	wire _169_;
	wire new_net_841;
	wire new_net_1040;
	wire new_net_1340;
	wire new_net_1352;
	wire new_net_1402;
	wire new_net_1565;
	wire new_net_1411;
	wire new_net_515;
	wire new_net_869;
	wire new_net_919;
	wire new_net_104;
	wire new_net_275;
	wire new_net_344;
	wire new_net_415;
	wire new_net_452;
	wire new_net_640;
	wire new_net_1022;
	wire _175_;
	wire new_net_1549;
	wire new_net_1134;
	wire new_net_393;
	wire new_net_732;
	wire _002_;
	wire _086_;
	wire _170_;
	wire new_net_156;
	wire new_net_258;
	wire new_net_1322;
	wire new_net_1669;
	wire new_net_1681;
	wire new_net_1921;
	wire new_net_1489;
	wire new_net_1812;
	wire new_net_1728;
	wire new_net_139;
	wire new_net_190;
	wire new_net_328;
	wire new_net_1151;
	wire new_net_1966;
	wire new_net_1990;
	wire new_net_2021;
	wire new_net_1943;
	wire new_net_1787;
	wire new_net_1834;
	wire new_net_444;
	wire _171_;
	wire _003_;
	wire _087_;
	wire new_net_412;
	wire new_net_964;
	wire new_net_975;
	wire new_net_987;
	wire new_net_1258;
	wire new_net_1445;
	wire new_net_1312;
	wire new_net_1597;
	wire new_net_1849;
	wire new_net_1184;
	wire new_net_626;
	wire new_net_671;
	wire new_net_637;
	wire new_net_660;
	wire new_net_754;
	wire new_net_648;
	wire new_net_765;
	wire new_net_105;
	wire new_net_276;
	wire new_net_484;
	wire new_net_1773;
	wire new_net_1118;
	wire new_net_420;
	wire _004_;
	wire _088_;
	wire _172_;
	wire new_net_1092;
	wire new_net_1410;
	wire new_net_1434;
	wire new_net_1545;
	wire new_net_1611;
	wire new_net_1623;
	wire new_net_644;
	wire new_net_827;
	wire new_net_788;
	wire new_net_1554;
	wire new_net_929;
	wire new_net_191;
	wire new_net_329;
	wire new_net_357;
	wire new_net_842;
	wire new_net_1041;
	wire new_net_1139;
	wire new_net_1341;
	wire new_net_1353;
	wire new_net_1393;
	wire new_net_1881;
	wire new_net_1923;
	wire new_net_2011;
	wire new_net_2048;
	wire new_net_1970;
	wire new_net_2017;
	wire new_net_1819;
	wire new_net_1939;
	wire new_net_920;
	wire new_net_345;
	wire _005_;
	wire _089_;
	wire _173_;
	wire new_net_1023;
	wire new_net_1158;
	wire new_net_1248;
	wire new_net_1289;
	wire new_net_1301;
	wire new_net_1618;
	wire new_net_1830;
	wire new_net_1945;
	wire new_net_1335;
	wire new_net_1792;
	wire new_net_516;
	wire new_net_733;
	wire new_net_106;
	wire new_net_157;
	wire new_net_259;
	wire new_net_394;
	wire new_net_453;
	wire new_net_560;
	wire new_net_1670;
	wire new_net_1682;
	wire new_net_1264;
	wire new_net_1593;
	wire new_net_1557;
	wire new_net_830;
	wire _006_;
	wire _090_;
	wire _174_;
	wire new_net_140;
	wire new_net_422;
	wire new_net_1063;
	wire new_net_1074;
	wire new_net_1152;
	wire new_net_1967;
	wire new_net_1778;
	wire new_net_1902;
	wire new_net_965;
	wire new_net_976;
	wire new_net_208;
	wire new_net_988;
	wire new_net_1013;
	wire new_net_1446;
	wire new_net_1458;
	wire new_net_1544;
	wire new_net_1635;
	wire new_net_1647;
	wire new_net_1675;
	wire new_net_651;
	wire new_net_661;
	wire new_net_755;
	wire new_net_627;
	wire new_net_672;
	wire new_net_871;
	wire new_net_766;
	wire new_net_638;
	wire new_net_277;
	wire new_net_346;
	wire new_net_649;
	wire new_net_1231;
	wire new_net_1398;
	wire new_net_1650;
	wire new_net_1886;
	wire new_net_1935;
	wire new_net_1928;
	wire new_net_759;
	wire new_net_2053;
	wire new_net_1975;
	wire new_net_844;
	wire new_net_955;
	wire new_net_107;
	wire new_net_158;
	wire new_net_260;
	wire new_net_395;
	wire new_net_485;
	wire new_net_506;
	wire new_net_744;
	wire new_net_1093;
	wire new_net_1496;
	wire new_net_1859;
	wire new_net_1824;
	wire new_net_398;
	wire new_net_1957;
	wire new_net_1950;
	wire new_net_831;
	wire new_net_930;
	wire new_net_192;
	wire new_net_330;
	wire new_net_954;
	wire _176_;
	wire _008_;
	wire _092_;
	wire new_net_141;
	wire new_net_1031;
	wire new_net_1872;
	wire new_net_1634;
	wire new_net_619;
	wire new_net_1732;
	wire new_net_861;
	wire new_net_879;
	wire new_net_886;
	wire new_net_921;
	wire new_net_1024;
	wire new_net_1249;
	wire new_net_1290;
	wire new_net_1302;
	wire new_net_1314;
	wire new_net_1527;
	wire new_net_1696;
	wire new_net_1734;
	input N1;
	input N101;
	input N106;
	input N111;
	input N116;
	input N121;
	input N126;
	input N13;
	input N130;
	input N135;
	input N138;
	input N143;
	input N146;
	input N149;
	input N152;
	input N153;
	input N156;
	input N159;
	input N165;
	input N17;
	input N171;
	input N177;
	input N183;
	input N189;
	input N195;
	input N201;
	input N207;
	input N210;
	input N219;
	input N228;
	input N237;
	input N246;
	input N255;
	input N259;
	input N26;
	input N260;
	input N261;
	input N267;
	input N268;
	input N29;
	input N36;
	input N42;
	input N51;
	input N55;
	input N59;
	input N68;
	input N72;
	input N73;
	input N74;
	input N75;
	input N8;
	input N80;
	input N85;
	input N86;
	input N87;
	input N88;
	input N89;
	input N90;
	input N91;
	input N96;
	output N388;
	output N389;
	output N390;
	output N391;
	output N418;
	output N419;
	output N420;
	output N421;
	output N422;
	output N423;
	output N446;
	output N447;
	output N448;
	output N449;
	output N450;
	output N767;
	output N768;
	output N850;
	output N863;
	output N864;
	output N865;
	output N866;
	output N874;
	output N878;
	output N879;
	output N880;

	or_bi _287_ (
		.a(new_net_202),
		.b(new_net_70),
		.c(_274_)
	);

	and_bi _288_ (
		.a(new_net_207),
		.b(new_net_76),
		.c(_275_)
	);

	and_bi _289_ (
		.a(_274_),
		.b(_275_),
		.c(_276_)
	);

	or_ii _290_ (
		.a(new_net_448),
		.b(new_net_108),
		.c(_277_)
	);

	or_bi _291_ (
		.a(new_net_343),
		.b(new_net_389),
		.c(_278_)
	);

	and_bb _292_ (
		.a(new_net_449),
		.b(new_net_44),
		.c(_279_)
	);

	or_bi _293_ (
		.a(new_net_356),
		.b(new_net_370),
		.c(_280_)
	);

	or_bb _294_ (
		.a(_280_),
		.b(new_net_450),
		.c(_281_)
	);

	inv _295_ (
		.din(new_net_204),
		.dout(_282_)
	);

	or_ii _296_ (
		.a(new_net_47),
		.b(new_net_138),
		.c(_283_)
	);

	or_bb _297_ (
		.a(new_net_27),
		.b(new_net_1),
		.c(_284_)
	);

	or_ii _298_ (
		.a(new_net_391),
		.b(new_net_74),
		.c(_285_)
	);

	or_ii _299_ (
		.a(new_net_187),
		.b(new_net_109),
		.c(_286_)
	);

	or_bb _300_ (
		.a(new_net_85),
		.b(_285_),
		.c(_000_)
	);

	and_bi _301_ (
		.a(_284_),
		.b(_000_),
		.c(_001_)
	);

	and_bi _302_ (
		.a(_281_),
		.b(new_net_451),
		.c(_002_)
	);

	or_bi _303_ (
		.a(new_net_291),
		.b(new_net_143),
		.c(_003_)
	);

	or_bb _304_ (
		.a(new_net_371),
		.b(new_net_358),
		.c(_004_)
	);

	or_bi _305_ (
		.a(new_net_330),
		.b(new_net_24),
		.c(_005_)
	);

	and_bi _306_ (
		.a(new_net_392),
		.b(new_net_347),
		.c(_006_)
	);

	and_bb _307_ (
		.a(new_net_309),
		.b(new_net_452),
		.c(_007_)
	);

	inv _308_ (
		.din(new_net_212),
		.dout(_008_)
	);

	or_ii _309_ (
		.a(new_net_139),
		.b(new_net_48),
		.c(_009_)
	);

	or_bb _310_ (
		.a(new_net_14),
		.b(new_net_394),
		.c(_010_)
	);

	or_bb _311_ (
		.a(new_net_453),
		.b(new_net_359),
		.c(_011_)
	);

	and_bi _312_ (
		.a(new_net_75),
		.b(new_net_29),
		.c(_012_)
	);

	and_bi _313_ (
		.a(new_net_454),
		.b(new_net_51),
		.c(_013_)
	);

	or_bb _314_ (
		.a(new_net_96),
		.b(new_net_455),
		.c(_014_)
	);

	or_bb _315_ (
		.a(_014_),
		.b(_006_),
		.c(_015_)
	);

	and_bi _316_ (
		.a(_003_),
		.b(_015_),
		.c(_016_)
	);

	or_bi _317_ (
		.a(new_net_111),
		.b(new_net_149),
		.c(_017_)
	);

	and_bi _318_ (
		.a(new_net_115),
		.b(new_net_150),
		.c(_018_)
	);

	and_bi _319_ (
		.a(new_net_164),
		.b(new_net_184),
		.c(_019_)
	);

	and_bi _320_ (
		.a(new_net_26),
		.b(new_net_52),
		.c(_020_)
	);

	and_bi _321_ (
		.a(_020_),
		.b(new_net_30),
		.c(_021_)
	);

	and_bi _322_ (
		.a(new_net_157),
		.b(new_net_296),
		.c(_022_)
	);

	and_bi _323_ (
		.a(new_net_71),
		.b(new_net_331),
		.c(_023_)
	);

	and_bi _324_ (
		.a(new_net_110),
		.b(_023_),
		.c(_024_)
	);

	and_bi _325_ (
		.a(new_net_328),
		.b(new_net_313),
		.c(_025_)
	);

	or_bb _326_ (
		.a(_025_),
		.b(new_net_456),
		.c(_026_)
	);

	and_ii _327_ (
		.a(_026_),
		.b(new_net_255),
		.c(_027_)
	);

	and_bi _328_ (
		.a(new_net_134),
		.b(new_net_372),
		.c(_028_)
	);

	and_bi _329_ (
		.a(new_net_374),
		.b(new_net_132),
		.c(_029_)
	);

	or_bi _330_ (
		.a(new_net_316),
		.b(new_net_345),
		.c(_030_)
	);

	and_bi _331_ (
		.a(new_net_170),
		.b(new_net_292),
		.c(_031_)
	);

	or_bb _332_ (
		.a(_031_),
		.b(new_net_258),
		.c(_032_)
	);

	and_bi _333_ (
		.a(_030_),
		.b(_032_),
		.c(_033_)
	);

	and_bi _334_ (
		.a(new_net_154),
		.b(new_net_67),
		.c(_034_)
	);

	or_bi _335_ (
		.a(new_net_153),
		.b(new_net_69),
		.c(_035_)
	);

	inv _336_ (
		.din(new_net_166),
		.dout(_036_)
	);

	or_bi _337_ (
		.a(new_net_315),
		.b(new_net_368),
		.c(_037_)
	);

	and_bi _338_ (
		.a(new_net_192),
		.b(new_net_295),
		.c(_038_)
	);

	or_bb _339_ (
		.a(_038_),
		.b(new_net_257),
		.c(_039_)
	);

	and_bi _340_ (
		.a(_037_),
		.b(_039_),
		.c(_040_)
	);

	or_bb _341_ (
		.a(new_net_189),
		.b(new_net_123),
		.c(_041_)
	);

	or_ii _342_ (
		.a(new_net_190),
		.b(new_net_124),
		.c(_042_)
	);

	or_bi _343_ (
		.a(new_net_314),
		.b(new_net_393),
		.c(_043_)
	);

	and_bi _344_ (
		.a(new_net_226),
		.b(new_net_297),
		.c(_044_)
	);

	or_bb _345_ (
		.a(_044_),
		.b(new_net_256),
		.c(_045_)
	);

	and_bi _346_ (
		.a(_043_),
		.b(_045_),
		.c(_046_)
	);

	and_bi _347_ (
		.a(new_net_325),
		.b(new_net_179),
		.c(_047_)
	);

	inv _348_ (
		.din(new_net_397),
		.dout(_048_)
	);

	and_bi _349_ (
		.a(new_net_180),
		.b(new_net_327),
		.c(_049_)
	);

	and_bi _350_ (
		.a(new_net_364),
		.b(new_net_381),
		.c(_050_)
	);

	or_bb _351_ (
		.a(_050_),
		.b(new_net_351),
		.c(_051_)
	);

	and_bi _352_ (
		.a(new_net_239),
		.b(new_net_16),
		.c(_052_)
	);

	and_bi _353_ (
		.a(new_net_223),
		.b(_052_),
		.c(_053_)
	);

	or_bi _354_ (
		.a(new_net_53),
		.b(new_net_102),
		.c(_054_)
	);

	and_bi _355_ (
		.a(_054_),
		.b(new_net_82),
		.c(_055_)
	);

	or_bb _356_ (
		.a(new_net_88),
		.b(new_net_399),
		.c(_056_)
	);

	and_bi _357_ (
		.a(_056_),
		.b(new_net_384),
		.c(_057_)
	);

	or_ii _358_ (
		.a(new_net_140),
		.b(new_net_266),
		.c(_058_)
	);

	and_bi _359_ (
		.a(_058_),
		.b(new_net_279),
		.c(_059_)
	);

	and_bi _360_ (
		.a(new_net_210),
		.b(_059_),
		.c(_060_)
	);

	and_bi _361_ (
		.a(new_net_264),
		.b(new_net_211),
		.c(_061_)
	);

	and_bi _362_ (
		.a(new_net_457),
		.b(new_net_142),
		.c(_062_)
	);

	inv _363_ (
		.din(new_net_302),
		.dout(_063_)
	);

	and_bi _364_ (
		.a(new_net_186),
		.b(new_net_251),
		.c(_064_)
	);

	and_bi _365_ (
		.a(new_net_317),
		.b(new_net_151),
		.c(_065_)
	);

	or_ii _366_ (
		.a(new_net_246),
		.b(new_net_25),
		.c(_066_)
	);

	and_ii _367_ (
		.a(new_net_458),
		.b(new_net_87),
		.c(_067_)
	);

	or_ii _368_ (
		.a(new_net_61),
		.b(new_net_46),
		.c(_068_)
	);

	and_bb _369_ (
		.a(new_net_459),
		.b(new_net_203),
		.c(_069_)
	);

	or_ii _370_ (
		.a(_069_),
		.b(new_net_460),
		.c(_070_)
	);

	and_ii _371_ (
		.a(_070_),
		.b(new_net_360),
		.c(_071_)
	);

	or_ii _372_ (
		.a(new_net_461),
		.b(new_net_332),
		.c(_072_)
	);

	and_bi _373_ (
		.a(new_net_112),
		.b(new_net_6),
		.c(_073_)
	);

	and_bb _374_ (
		.a(new_net_232),
		.b(new_net_127),
		.c(_074_)
	);

	or_bb _375_ (
		.a(new_net_462),
		.b(_073_),
		.c(_075_)
	);

	or_bb _376_ (
		.a(new_net_463),
		.b(_065_),
		.c(_076_)
	);

	or_bb _377_ (
		.a(new_net_464),
		.b(_064_),
		.c(_077_)
	);

	or_bb _378_ (
		.a(new_net_465),
		.b(_062_),
		.c(_078_)
	);

	or_bb _379_ (
		.a(new_net_466),
		.b(_060_),
		.c(new_net_542)
	);

	or_bi _380_ (
		.a(new_net_298),
		.b(new_net_104),
		.c(_079_)
	);

	and_bi _381_ (
		.a(new_net_329),
		.b(new_net_348),
		.c(_080_)
	);

	and_bb _382_ (
		.a(new_net_312),
		.b(new_net_188),
		.c(_081_)
	);

	or_bb _383_ (
		.a(new_net_467),
		.b(new_net_99),
		.c(_082_)
	);

	or_bb _384_ (
		.a(_082_),
		.b(_080_),
		.c(_083_)
	);

	and_bi _385_ (
		.a(_079_),
		.b(_083_),
		.c(_084_)
	);

	and_bi _386_ (
		.a(new_net_39),
		.b(new_net_241),
		.c(_085_)
	);

	and_bi _387_ (
		.a(new_net_242),
		.b(new_net_38),
		.c(_086_)
	);

	and_ii _388_ (
		.a(new_net_289),
		.b(new_net_274),
		.c(_087_)
	);

	or_bi _389_ (
		.a(new_net_293),
		.b(new_net_119),
		.c(_088_)
	);

	and_bi _390_ (
		.a(new_net_346),
		.b(new_net_349),
		.c(_089_)
	);

	and_bb _391_ (
		.a(new_net_310),
		.b(new_net_390),
		.c(_090_)
	);

	or_bb _392_ (
		.a(new_net_468),
		.b(new_net_97),
		.c(_091_)
	);

	or_bb _393_ (
		.a(_091_),
		.b(_089_),
		.c(_092_)
	);

	and_bi _394_ (
		.a(_088_),
		.b(_092_),
		.c(_093_)
	);

	and_bi _395_ (
		.a(new_net_56),
		.b(new_net_19),
		.c(_094_)
	);

	and_bi _396_ (
		.a(new_net_20),
		.b(new_net_60),
		.c(_095_)
	);

	or_bi _397_ (
		.a(new_net_294),
		.b(new_net_128),
		.c(_096_)
	);

	and_bi _398_ (
		.a(new_net_369),
		.b(new_net_350),
		.c(_097_)
	);

	and_bb _399_ (
		.a(new_net_311),
		.b(new_net_72),
		.c(_098_)
	);

	or_bb _400_ (
		.a(new_net_469),
		.b(new_net_98),
		.c(_099_)
	);

	or_bb _401_ (
		.a(_099_),
		.b(_097_),
		.c(_100_)
	);

	and_bi _402_ (
		.a(_096_),
		.b(_100_),
		.c(_101_)
	);

	and_bi _403_ (
		.a(new_net_91),
		.b(new_net_161),
		.c(_102_)
	);

	and_bi _404_ (
		.a(new_net_163),
		.b(new_net_94),
		.c(_103_)
	);

	or_bi _405_ (
		.a(new_net_141),
		.b(new_net_165),
		.c(_104_)
	);

	and_bi _406_ (
		.a(_104_),
		.b(new_net_185),
		.c(_105_)
	);

	or_bb _407_ (
		.a(new_net_261),
		.b(new_net_218),
		.c(_106_)
	);

	and_bi _408_ (
		.a(_106_),
		.b(new_net_176),
		.c(_107_)
	);

	or_bb _409_ (
		.a(new_net_299),
		.b(new_net_63),
		.c(_108_)
	);

	and_bi _410_ (
		.a(_108_),
		.b(new_net_41),
		.c(_109_)
	);

	or_bi _411_ (
		.a(new_net_306),
		.b(new_net_340),
		.c(_110_)
	);

	inv _412_ (
		.din(new_net_268),
		.dout(_111_)
	);

	and_bi _413_ (
		.a(new_net_307),
		.b(new_net_341),
		.c(_112_)
	);

	or_bb _414_ (
		.a(_112_),
		.b(new_net_375),
		.c(_113_)
	);

	and_bi _415_ (
		.a(new_net_470),
		.b(_113_),
		.c(_114_)
	);

	and_bb _416_ (
		.a(new_net_308),
		.b(new_net_284),
		.c(_115_)
	);

	and_bi _417_ (
		.a(new_net_276),
		.b(new_net_249),
		.c(_116_)
	);

	and_bi _418_ (
		.a(new_net_322),
		.b(new_net_243),
		.c(_117_)
	);

	and_bi _419_ (
		.a(new_net_37),
		.b(new_net_8),
		.c(_118_)
	);

	and_bb _420_ (
		.a(new_net_233),
		.b(new_net_31),
		.c(_119_)
	);

	or_bb _421_ (
		.a(new_net_471),
		.b(_118_),
		.c(_120_)
	);

	or_bb _422_ (
		.a(new_net_472),
		.b(_117_),
		.c(_121_)
	);

	or_bb _423_ (
		.a(new_net_473),
		.b(_116_),
		.c(_122_)
	);

	or_bb _424_ (
		.a(new_net_474),
		.b(_115_),
		.c(_123_)
	);

	or_bb _425_ (
		.a(new_net_475),
		.b(_114_),
		.c(N878)
	);

	and_ii _426_ (
		.a(new_net_64),
		.b(new_net_43),
		.c(_124_)
	);

	or_bi _427_ (
		.a(new_net_300),
		.b(new_net_196),
		.c(_125_)
	);

	and_bi _428_ (
		.a(new_net_301),
		.b(new_net_197),
		.c(_126_)
	);

	or_bb _429_ (
		.a(_126_),
		.b(new_net_377),
		.c(_127_)
	);

	and_bi _430_ (
		.a(new_net_476),
		.b(_127_),
		.c(_128_)
	);

	and_bb _431_ (
		.a(new_net_198),
		.b(new_net_281),
		.c(_129_)
	);

	and_bi _432_ (
		.a(new_net_42),
		.b(new_net_253),
		.c(_130_)
	);

	and_bi _433_ (
		.a(new_net_318),
		.b(new_net_21),
		.c(_131_)
	);

	and_bb _434_ (
		.a(new_net_229),
		.b(new_net_106),
		.c(_132_)
	);

	and_bi _435_ (
		.a(new_net_59),
		.b(new_net_11),
		.c(_133_)
	);

	or_bb _436_ (
		.a(_133_),
		.b(new_net_477),
		.c(_134_)
	);

	or_bb _437_ (
		.a(new_net_478),
		.b(_131_),
		.c(_135_)
	);

	or_bb _438_ (
		.a(new_net_479),
		.b(_130_),
		.c(_136_)
	);

	or_bb _439_ (
		.a(new_net_480),
		.b(_129_),
		.c(_137_)
	);

	or_bb _440_ (
		.a(new_net_481),
		.b(_128_),
		.c(new_net_548)
	);

	and_ii _441_ (
		.a(new_net_219),
		.b(new_net_178),
		.c(_138_)
	);

	or_bi _442_ (
		.a(new_net_263),
		.b(new_net_77),
		.c(_139_)
	);

	and_bi _443_ (
		.a(new_net_262),
		.b(new_net_79),
		.c(_140_)
	);

	or_bb _444_ (
		.a(_140_),
		.b(new_net_378),
		.c(_141_)
	);

	and_bi _445_ (
		.a(new_net_482),
		.b(_141_),
		.c(_142_)
	);

	and_bb _446_ (
		.a(new_net_78),
		.b(new_net_280),
		.c(_143_)
	);

	and_bi _447_ (
		.a(new_net_177),
		.b(new_net_252),
		.c(_144_)
	);

	and_bi _448_ (
		.a(new_net_319),
		.b(new_net_162),
		.c(_145_)
	);

	and_bb _449_ (
		.a(new_net_234),
		.b(new_net_121),
		.c(_146_)
	);

	and_bi _450_ (
		.a(new_net_93),
		.b(new_net_7),
		.c(_147_)
	);

	or_bb _451_ (
		.a(_147_),
		.b(new_net_483),
		.c(_148_)
	);

	or_bb _452_ (
		.a(new_net_484),
		.b(_145_),
		.c(_149_)
	);

	or_bb _453_ (
		.a(new_net_485),
		.b(_144_),
		.c(_150_)
	);

	or_bb _454_ (
		.a(new_net_486),
		.b(_143_),
		.c(_151_)
	);

	or_bb _455_ (
		.a(new_net_487),
		.b(_142_),
		.c(new_net_532)
	);

	and_ii _456_ (
		.a(new_net_400),
		.b(new_net_386),
		.c(_152_)
	);

	and_bi _457_ (
		.a(new_net_90),
		.b(new_net_353),
		.c(_153_)
	);

	and_bi _458_ (
		.a(new_net_354),
		.b(new_net_89),
		.c(_154_)
	);

	or_bb _459_ (
		.a(_154_),
		.b(_153_),
		.c(_155_)
	);

	and_bi _460_ (
		.a(new_net_265),
		.b(_155_),
		.c(_156_)
	);

	and_bb _461_ (
		.a(new_net_355),
		.b(new_net_285),
		.c(_157_)
	);

	and_bi _462_ (
		.a(new_net_385),
		.b(new_net_248),
		.c(_158_)
	);

	and_bi _463_ (
		.a(new_net_323),
		.b(new_net_373),
		.c(_159_)
	);

	and_bi _464_ (
		.a(new_net_131),
		.b(new_net_9),
		.c(_160_)
	);

	and_bb _465_ (
		.a(new_net_235),
		.b(new_net_146),
		.c(_161_)
	);

	or_bb _466_ (
		.a(new_net_488),
		.b(_160_),
		.c(_162_)
	);

	or_bb _467_ (
		.a(new_net_489),
		.b(_159_),
		.c(_163_)
	);

	or_bb _468_ (
		.a(new_net_490),
		.b(_158_),
		.c(_164_)
	);

	or_bb _469_ (
		.a(new_net_491),
		.b(_157_),
		.c(_165_)
	);

	or_bb _470_ (
		.a(new_net_492),
		.b(_156_),
		.c(new_net_564)
	);

	and_bi _471_ (
		.a(new_net_103),
		.b(new_net_84),
		.c(_166_)
	);

	and_bi _472_ (
		.a(new_net_55),
		.b(new_net_199),
		.c(_167_)
	);

	and_bi _473_ (
		.a(new_net_200),
		.b(new_net_54),
		.c(_168_)
	);

	or_bb _474_ (
		.a(_168_),
		.b(_167_),
		.c(_169_)
	);

	and_bi _475_ (
		.a(new_net_267),
		.b(_169_),
		.c(_170_)
	);

	and_bb _476_ (
		.a(new_net_201),
		.b(new_net_282),
		.c(_171_)
	);

	and_bi _477_ (
		.a(new_net_83),
		.b(new_net_254),
		.c(_172_)
	);

	and_bi _478_ (
		.a(new_net_320),
		.b(new_net_68),
		.c(_173_)
	);

	and_bi _479_ (
		.a(new_net_155),
		.b(new_net_12),
		.c(_174_)
	);

	and_bb _480_ (
		.a(new_net_230),
		.b(new_net_160),
		.c(_175_)
	);

	and_bb _481_ (
		.a(new_net_493),
		.b(new_net_335),
		.c(_176_)
	);

	or_bb _482_ (
		.a(new_net_494),
		.b(_175_),
		.c(_177_)
	);

	or_bb _483_ (
		.a(new_net_495),
		.b(_174_),
		.c(_178_)
	);

	or_bb _484_ (
		.a(new_net_496),
		.b(_173_),
		.c(_179_)
	);

	or_bb _485_ (
		.a(new_net_497),
		.b(_172_),
		.c(_180_)
	);

	or_bb _486_ (
		.a(new_net_498),
		.b(_171_),
		.c(_181_)
	);

	or_bb _487_ (
		.a(new_net_499),
		.b(_170_),
		.c(new_net_530)
	);

	and_ii _488_ (
		.a(new_net_383),
		.b(new_net_352),
		.c(_182_)
	);

	or_ii _489_ (
		.a(new_net_116),
		.b(new_net_398),
		.c(_183_)
	);

	and_bi _490_ (
		.a(new_net_365),
		.b(new_net_117),
		.c(_184_)
	);

	or_bb _491_ (
		.a(_184_),
		.b(new_net_376),
		.c(_185_)
	);

	and_bi _492_ (
		.a(new_net_500),
		.b(_185_),
		.c(_186_)
	);

	and_bb _493_ (
		.a(new_net_118),
		.b(new_net_286),
		.c(_187_)
	);

	and_bi _494_ (
		.a(new_net_382),
		.b(new_net_250),
		.c(_188_)
	);

	and_bi _495_ (
		.a(new_net_324),
		.b(new_net_326),
		.c(_189_)
	);

	and_bi _496_ (
		.a(new_net_182),
		.b(new_net_10),
		.c(_190_)
	);

	and_bb _497_ (
		.a(new_net_501),
		.b(new_net_337),
		.c(_191_)
	);

	and_bb _498_ (
		.a(new_net_231),
		.b(new_net_195),
		.c(_192_)
	);

	or_bb _499_ (
		.a(_192_),
		.b(new_net_502),
		.c(_193_)
	);

	or_bb _500_ (
		.a(new_net_503),
		.b(_190_),
		.c(_194_)
	);

	or_bb _501_ (
		.a(new_net_504),
		.b(_189_),
		.c(_195_)
	);

	or_bb _502_ (
		.a(new_net_505),
		.b(_188_),
		.c(_196_)
	);

	or_bb _503_ (
		.a(new_net_506),
		.b(_187_),
		.c(_197_)
	);

	or_bb _504_ (
		.a(new_net_507),
		.b(_186_),
		.c(new_net_544)
	);

	and_bb _505_ (
		.a(new_net_240),
		.b(new_net_224),
		.c(_198_)
	);

	and_bi _506_ (
		.a(new_net_17),
		.b(new_net_3),
		.c(_199_)
	);

	and_bi _507_ (
		.a(new_net_4),
		.b(new_net_18),
		.c(_200_)
	);

	or_bb _508_ (
		.a(_200_),
		.b(_199_),
		.c(_201_)
	);

	and_bi _509_ (
		.a(new_net_269),
		.b(_201_),
		.c(_202_)
	);

	and_bb _510_ (
		.a(new_net_5),
		.b(new_net_283),
		.c(_203_)
	);

	and_bi _511_ (
		.a(new_net_303),
		.b(new_net_225),
		.c(_204_)
	);

	and_bi _512_ (
		.a(new_net_321),
		.b(new_net_191),
		.c(_205_)
	);

	and_bi _513_ (
		.a(new_net_168),
		.b(new_net_13),
		.c(_206_)
	);

	and_bb _514_ (
		.a(new_net_508),
		.b(new_net_336),
		.c(_207_)
	);

	and_bb _515_ (
		.a(new_net_236),
		.b(new_net_173),
		.c(_208_)
	);

	or_bb _516_ (
		.a(_208_),
		.b(new_net_509),
		.c(_209_)
	);

	or_bb _517_ (
		.a(new_net_510),
		.b(_206_),
		.c(_210_)
	);

	or_bb _518_ (
		.a(new_net_511),
		.b(_205_),
		.c(_211_)
	);

	or_bb _519_ (
		.a(new_net_512),
		.b(_204_),
		.c(_212_)
	);

	or_bb _520_ (
		.a(new_net_513),
		.b(_203_),
		.c(_213_)
	);

	or_bb _521_ (
		.a(new_net_514),
		.b(_202_),
		.c(new_net_522)
	);

	and_ii _522_ (
		.a(new_net_342),
		.b(new_net_290),
		.c(_214_)
	);

	or_bb _523_ (
		.a(_214_),
		.b(new_net_275),
		.c(new_net_566)
	);

	or_ii _524_ (
		.a(new_net_62),
		.b(new_net_50),
		.c(_215_)
	);

	and_bi _525_ (
		.a(new_net_334),
		.b(new_net_515),
		.c(new_net_550)
	);

	or_ii _526_ (
		.a(new_net_45),
		.b(new_net_65),
		.c(_216_)
	);

	or_bb _527_ (
		.a(new_net_366),
		.b(new_net_2),
		.c(new_net_554)
	);

	or_bb _528_ (
		.a(new_net_367),
		.b(new_net_396),
		.c(new_net_524)
	);

	or_bb _529_ (
		.a(new_net_28),
		.b(new_net_395),
		.c(new_net_562)
	);

	or_ii _530_ (
		.a(new_net_66),
		.b(new_net_49),
		.c(_217_)
	);

	and_bi _531_ (
		.a(new_net_206),
		.b(new_net_379),
		.c(new_net_0)
	);

	or_bb _532_ (
		.a(new_net_113),
		.b(new_net_36),
		.c(_218_)
	);

	and_bb _533_ (
		.a(new_net_114),
		.b(new_net_40),
		.c(_219_)
	);

	and_bi _534_ (
		.a(_218_),
		.b(_219_),
		.c(_220_)
	);

	and_bi _535_ (
		.a(new_net_270),
		.b(new_net_34),
		.c(_221_)
	);

	and_bi _536_ (
		.a(new_net_35),
		.b(new_net_272),
		.c(_222_)
	);

	and_ii _537_ (
		.a(_222_),
		.b(_221_),
		.c(_223_)
	);

	and_ii _538_ (
		.a(new_net_169),
		.b(new_net_152),
		.c(_224_)
	);

	and_bb _539_ (
		.a(new_net_167),
		.b(new_net_156),
		.c(_225_)
	);

	and_ii _540_ (
		.a(_225_),
		.b(_224_),
		.c(_226_)
	);

	and_bi _541_ (
		.a(new_net_216),
		.b(new_net_147),
		.c(_227_)
	);

	and_bi _542_ (
		.a(new_net_148),
		.b(new_net_217),
		.c(_228_)
	);

	or_bb _543_ (
		.a(_228_),
		.b(_227_),
		.c(_229_)
	);

	or_bi _544_ (
		.a(new_net_57),
		.b(new_net_181),
		.c(_230_)
	);

	and_bi _545_ (
		.a(new_net_58),
		.b(new_net_183),
		.c(_231_)
	);

	and_bi _546_ (
		.a(_230_),
		.b(_231_),
		.c(_232_)
	);

	and_bi _547_ (
		.a(new_net_95),
		.b(new_net_135),
		.c(_233_)
	);

	and_bi _548_ (
		.a(new_net_133),
		.b(new_net_92),
		.c(_234_)
	);

	or_bb _549_ (
		.a(_234_),
		.b(_233_),
		.c(_235_)
	);

	and_ii _550_ (
		.a(new_net_338),
		.b(new_net_277),
		.c(_236_)
	);

	and_bb _551_ (
		.a(new_net_339),
		.b(new_net_278),
		.c(_237_)
	);

	and_ii _552_ (
		.a(_237_),
		.b(_236_),
		.c(_238_)
	);

	and_ii _553_ (
		.a(new_net_387),
		.b(new_net_214),
		.c(_239_)
	);

	and_bb _554_ (
		.a(new_net_388),
		.b(new_net_215),
		.c(_240_)
	);

	and_ii _555_ (
		.a(_240_),
		.b(_239_),
		.c(_241_)
	);

	and_bi _556_ (
		.a(new_net_32),
		.b(new_net_100),
		.c(_242_)
	);

	and_bi _557_ (
		.a(new_net_101),
		.b(new_net_33),
		.c(_243_)
	);

	or_bb _558_ (
		.a(_243_),
		.b(_242_),
		.c(new_net_560)
	);

	and_ii _559_ (
		.a(new_net_273),
		.b(new_net_120),
		.c(_244_)
	);

	and_bb _560_ (
		.a(new_net_271),
		.b(new_net_122),
		.c(_245_)
	);

	or_bb _561_ (
		.a(_245_),
		.b(_244_),
		.c(_246_)
	);

	and_bi _562_ (
		.a(new_net_107),
		.b(new_net_125),
		.c(_247_)
	);

	and_bi _563_ (
		.a(new_net_126),
		.b(new_net_105),
		.c(_248_)
	);

	and_ii _564_ (
		.a(_248_),
		.b(_247_),
		.c(_249_)
	);

	and_ii _565_ (
		.a(new_net_287),
		.b(new_net_193),
		.c(_250_)
	);

	and_bb _566_ (
		.a(new_net_288),
		.b(new_net_194),
		.c(_251_)
	);

	and_ii _567_ (
		.a(_251_),
		.b(_250_),
		.c(_252_)
	);

	and_bi _568_ (
		.a(new_net_228),
		.b(new_net_244),
		.c(_253_)
	);

	and_bi _569_ (
		.a(new_net_245),
		.b(new_net_227),
		.c(_254_)
	);

	or_bb _570_ (
		.a(_254_),
		.b(_253_),
		.c(_255_)
	);

	and_bi _571_ (
		.a(new_net_130),
		.b(new_net_144),
		.c(_256_)
	);

	and_bi _572_ (
		.a(new_net_145),
		.b(new_net_129),
		.c(_257_)
	);

	and_ii _573_ (
		.a(_257_),
		.b(_256_),
		.c(_258_)
	);

	and_ii _574_ (
		.a(new_net_158),
		.b(new_net_171),
		.c(_259_)
	);

	and_bb _575_ (
		.a(new_net_159),
		.b(new_net_172),
		.c(_260_)
	);

	and_ii _576_ (
		.a(_260_),
		.b(_259_),
		.c(_261_)
	);

	and_bi _577_ (
		.a(new_net_362),
		.b(new_net_22),
		.c(_262_)
	);

	and_bi _578_ (
		.a(new_net_23),
		.b(new_net_363),
		.c(_263_)
	);

	and_ii _579_ (
		.a(_263_),
		.b(_262_),
		.c(_264_)
	);

	and_ii _580_ (
		.a(new_net_80),
		.b(new_net_304),
		.c(_265_)
	);

	and_bb _581_ (
		.a(new_net_81),
		.b(new_net_305),
		.c(_266_)
	);

	and_ii _582_ (
		.a(_266_),
		.b(_265_),
		.c(_267_)
	);

	and_bi _583_ (
		.a(new_net_136),
		.b(new_net_174),
		.c(_268_)
	);

	and_bi _584_ (
		.a(new_net_175),
		.b(new_net_137),
		.c(_269_)
	);

	or_bb _585_ (
		.a(_269_),
		.b(_268_),
		.c(new_net_520)
	);

	or_bi _586_ (
		.a(new_net_361),
		.b(new_net_516),
		.c(_270_)
	);

	and_bi _587_ (
		.a(new_net_333),
		.b(new_net_517),
		.c(new_net_534)
	);

	and_bi _588_ (
		.a(new_net_205),
		.b(new_net_15),
		.c(new_net_546)
	);

	and_bi _589_ (
		.a(new_net_213),
		.b(new_net_380),
		.c(new_net_552)
	);

	and_bb _590_ (
		.a(N86),
		.b(N85),
		.c(new_net_526)
	);

	inv _591_ (
		.din(new_net_357),
		.dout(new_net_536)
	);

	or_ii _592_ (
		.a(new_net_247),
		.b(new_net_73),
		.c(_271_)
	);

	and_ii _593_ (
		.a(new_net_208),
		.b(new_net_86),
		.c(new_net_540)
	);

	or_bb _594_ (
		.a(new_net_209),
		.b(new_net_344),
		.c(_272_)
	);

	or_bi _595_ (
		.a(new_net_237),
		.b(new_net_222),
		.c(new_net_556)
	);

	and_ii _596_ (
		.a(N88),
		.b(N87),
		.c(_273_)
	);

	and_bi _597_ (
		.a(new_net_518),
		.b(new_net_259),
		.c(new_net_558)
	);

	and_bi _598_ (
		.a(new_net_519),
		.b(new_net_260),
		.c(new_net_538)
	);

	or_bb _599_ (
		.a(new_net_238),
		.b(new_net_221),
		.c(new_net_528)
	);

	spl2 new_net_442_v_fanout (
		.a(new_net_442),
		.b(new_net_307),
		.c(new_net_306)
	);

	spl3L _109__v_fanout (
		.a(_109_),
		.b(new_net_342),
		.c(new_net_340),
		.d(new_net_341)
	);

	bfr new_net_568_bfr_before (
		.din(new_net_568),
		.dout(new_net_375)
	);

	bfr new_net_569_bfr_before (
		.din(new_net_569),
		.dout(new_net_568)
	);

	bfr new_net_570_bfr_before (
		.din(new_net_570),
		.dout(new_net_569)
	);

	spl2 new_net_437_v_fanout (
		.a(new_net_437),
		.b(new_net_570),
		.c(new_net_377)
	);

	spl3L _107__v_fanout (
		.a(_107_),
		.b(new_net_300),
		.c(new_net_299),
		.d(new_net_301)
	);

	spl2 new_net_443_v_fanout (
		.a(new_net_443),
		.b(new_net_197),
		.c(new_net_196)
	);

	bfr new_net_571_bfr_before (
		.din(new_net_571),
		.dout(new_net_437)
	);

	bfr new_net_572_bfr_before (
		.din(new_net_572),
		.dout(new_net_571)
	);

	spl2 new_net_436_v_fanout (
		.a(new_net_436),
		.b(new_net_572),
		.c(new_net_378)
	);

	spl3L _105__v_fanout (
		.a(_105_),
		.b(new_net_262),
		.c(new_net_261),
		.d(new_net_263)
	);

	spl2 new_net_444_v_fanout (
		.a(new_net_444),
		.b(new_net_79),
		.c(new_net_77)
	);

	spl3L _057__v_fanout (
		.a(_057_),
		.b(new_net_142),
		.c(new_net_140),
		.d(new_net_141)
	);

	bfr new_net_573_bfr_before (
		.din(new_net_573),
		.dout(new_net_266)
	);

	spl2 new_net_423_v_fanout (
		.a(new_net_423),
		.b(new_net_573),
		.c(new_net_265)
	);

	spl2 new_net_447_v_fanout (
		.a(new_net_447),
		.b(new_net_354),
		.c(new_net_353)
	);

	spl3L _055__v_fanout (
		.a(_055_),
		.b(new_net_89),
		.c(new_net_88),
		.d(new_net_90)
	);

	bfr new_net_574_bfr_before (
		.din(new_net_574),
		.dout(new_net_423)
	);

	bfr new_net_575_bfr_before (
		.din(new_net_575),
		.dout(new_net_574)
	);

	spl2 new_net_422_v_fanout (
		.a(new_net_422),
		.b(new_net_575),
		.c(new_net_267)
	);

	spl3L _053__v_fanout (
		.a(_053_),
		.b(new_net_55),
		.c(new_net_53),
		.d(new_net_54)
	);

	spl2 new_net_445_v_fanout (
		.a(new_net_445),
		.b(new_net_200),
		.c(new_net_199)
	);

	bfr new_net_576_bfr_before (
		.din(new_net_576),
		.dout(new_net_422)
	);

	bfr new_net_577_bfr_before (
		.din(new_net_577),
		.dout(new_net_576)
	);

	spl2 new_net_421_v_fanout (
		.a(new_net_421),
		.b(new_net_577),
		.c(new_net_269)
	);

	spl2 new_net_446_v_fanout (
		.a(new_net_446),
		.b(new_net_4),
		.c(new_net_3)
	);

	spl3L _051__v_fanout (
		.a(_051_),
		.b(new_net_18),
		.c(new_net_16),
		.d(new_net_17)
	);

	bfr new_net_578_bfr_before (
		.din(new_net_578),
		.dout(new_net_447)
	);

	bfr new_net_579_bfr_before (
		.din(new_net_579),
		.dout(new_net_578)
	);

	bfr new_net_580_bfr_before (
		.din(new_net_580),
		.dout(new_net_579)
	);

	bfr new_net_581_bfr_before (
		.din(new_net_581),
		.dout(new_net_580)
	);

	bfr new_net_582_bfr_before (
		.din(new_net_582),
		.dout(new_net_581)
	);

	spl2 _152__v_fanout (
		.a(_152_),
		.b(new_net_355),
		.c(new_net_582)
	);

	bfr new_net_583_bfr_before (
		.din(new_net_583),
		.dout(new_net_279)
	);

	bfr new_net_584_bfr_before (
		.din(new_net_584),
		.dout(new_net_583)
	);

	bfr new_net_585_bfr_before (
		.din(new_net_585),
		.dout(new_net_584)
	);

	bfr new_net_586_bfr_before (
		.din(new_net_586),
		.dout(new_net_585)
	);

	bfr new_net_587_bfr_before (
		.din(new_net_587),
		.dout(new_net_586)
	);

	bfr new_net_588_bfr_before (
		.din(new_net_588),
		.dout(new_net_587)
	);

	bfr new_net_589_bfr_before (
		.din(new_net_589),
		.dout(new_net_588)
	);

	bfr new_net_590_bfr_before (
		.din(new_net_590),
		.dout(new_net_589)
	);

	bfr new_net_591_bfr_before (
		.din(new_net_591),
		.dout(new_net_590)
	);

	bfr new_net_592_bfr_before (
		.din(new_net_592),
		.dout(new_net_591)
	);

	spl2 new_net_425_v_fanout (
		.a(new_net_425),
		.b(new_net_592),
		.c(new_net_285)
	);

	spl2 _198__v_fanout (
		.a(_198_),
		.b(new_net_5),
		.c(new_net_446)
	);

	spl4L new_net_424_v_fanout (
		.a(new_net_424),
		.b(new_net_286),
		.c(new_net_283),
		.d(new_net_425),
		.e(new_net_282)
	);

	bfr new_net_593_bfr_before (
		.din(new_net_593),
		.dout(new_net_445)
	);

	bfr new_net_594_bfr_before (
		.din(new_net_594),
		.dout(new_net_593)
	);

	bfr new_net_595_bfr_before (
		.din(new_net_595),
		.dout(new_net_594)
	);

	spl2 _166__v_fanout (
		.a(_166_),
		.b(new_net_201),
		.c(new_net_595)
	);

	spl3L _182__v_fanout (
		.a(_182_),
		.b(new_net_118),
		.c(new_net_116),
		.d(new_net_117)
	);

	bfr new_net_596_bfr_before (
		.din(new_net_596),
		.dout(new_net_384)
	);

	bfr new_net_597_bfr_before (
		.din(new_net_597),
		.dout(new_net_596)
	);

	bfr new_net_598_bfr_before (
		.din(new_net_598),
		.dout(new_net_597)
	);

	bfr new_net_599_bfr_before (
		.din(new_net_599),
		.dout(new_net_598)
	);

	bfr new_net_600_bfr_before (
		.din(new_net_600),
		.dout(new_net_599)
	);

	bfr new_net_601_bfr_before (
		.din(new_net_601),
		.dout(new_net_600)
	);

	bfr new_net_602_bfr_before (
		.din(new_net_602),
		.dout(new_net_601)
	);

	bfr new_net_603_bfr_before (
		.din(new_net_603),
		.dout(new_net_602)
	);

	bfr new_net_604_bfr_before (
		.din(new_net_604),
		.dout(new_net_603)
	);

	spl3L _028__v_fanout (
		.a(_028_),
		.b(new_net_385),
		.c(new_net_604),
		.d(new_net_386)
	);

	bfr new_net_605_bfr_before (
		.din(new_net_605),
		.dout(new_net_421)
	);

	bfr new_net_606_bfr_before (
		.din(new_net_606),
		.dout(new_net_605)
	);

	bfr new_net_607_bfr_before (
		.din(new_net_607),
		.dout(new_net_606)
	);

	spl2 new_net_420_v_fanout (
		.a(new_net_420),
		.b(new_net_607),
		.c(new_net_264)
	);

	bfr new_net_608_bfr_before (
		.din(new_net_608),
		.dout(new_net_444)
	);

	bfr new_net_609_bfr_before (
		.din(new_net_609),
		.dout(new_net_608)
	);

	bfr new_net_610_bfr_before (
		.din(new_net_610),
		.dout(new_net_609)
	);

	bfr new_net_611_bfr_before (
		.din(new_net_611),
		.dout(new_net_610)
	);

	bfr new_net_612_bfr_before (
		.din(new_net_612),
		.dout(new_net_611)
	);

	bfr new_net_613_bfr_before (
		.din(new_net_613),
		.dout(new_net_612)
	);

	bfr new_net_614_bfr_before (
		.din(new_net_614),
		.dout(new_net_613)
	);

	bfr new_net_615_bfr_before (
		.din(new_net_615),
		.dout(new_net_614)
	);

	bfr new_net_616_bfr_before (
		.din(new_net_616),
		.dout(new_net_615)
	);

	bfr new_net_617_bfr_before (
		.din(new_net_617),
		.dout(new_net_616)
	);

	bfr new_net_618_bfr_before (
		.din(new_net_618),
		.dout(new_net_617)
	);

	bfr new_net_619_bfr_before (
		.din(new_net_619),
		.dout(new_net_618)
	);

	bfr new_net_620_bfr_before (
		.din(new_net_620),
		.dout(new_net_619)
	);

	spl2 _138__v_fanout (
		.a(_138_),
		.b(new_net_78),
		.c(new_net_620)
	);

	bfr new_net_621_bfr_before (
		.din(new_net_621),
		.dout(new_net_210)
	);

	bfr new_net_622_bfr_before (
		.din(new_net_622),
		.dout(new_net_621)
	);

	bfr new_net_623_bfr_before (
		.din(new_net_623),
		.dout(new_net_622)
	);

	bfr new_net_624_bfr_before (
		.din(new_net_624),
		.dout(new_net_623)
	);

	bfr new_net_625_bfr_before (
		.din(new_net_625),
		.dout(new_net_624)
	);

	bfr new_net_626_bfr_before (
		.din(new_net_626),
		.dout(new_net_625)
	);

	bfr new_net_627_bfr_before (
		.din(new_net_627),
		.dout(new_net_626)
	);

	bfr new_net_628_bfr_before (
		.din(new_net_628),
		.dout(new_net_627)
	);

	bfr new_net_629_bfr_before (
		.din(new_net_629),
		.dout(new_net_628)
	);

	bfr new_net_630_bfr_before (
		.din(new_net_630),
		.dout(new_net_629)
	);

	bfr new_net_631_bfr_before (
		.din(new_net_631),
		.dout(new_net_630)
	);

	bfr new_net_632_bfr_before (
		.din(new_net_632),
		.dout(new_net_631)
	);

	bfr new_net_633_bfr_before (
		.din(new_net_633),
		.dout(new_net_632)
	);

	spl2 _019__v_fanout (
		.a(_019_),
		.b(new_net_211),
		.c(new_net_633)
	);

	bfr new_net_634_bfr_before (
		.din(new_net_634),
		.dout(new_net_399)
	);

	bfr new_net_635_bfr_before (
		.din(new_net_635),
		.dout(new_net_634)
	);

	bfr new_net_636_bfr_before (
		.din(new_net_636),
		.dout(new_net_635)
	);

	bfr new_net_637_bfr_before (
		.din(new_net_637),
		.dout(new_net_636)
	);

	bfr new_net_638_bfr_before (
		.din(new_net_638),
		.dout(new_net_637)
	);

	bfr new_net_639_bfr_before (
		.din(new_net_639),
		.dout(new_net_638)
	);

	bfr new_net_640_bfr_before (
		.din(new_net_640),
		.dout(new_net_639)
	);

	bfr new_net_641_bfr_before (
		.din(new_net_641),
		.dout(new_net_640)
	);

	spl2 _029__v_fanout (
		.a(_029_),
		.b(new_net_400),
		.c(new_net_641)
	);

	bfr new_net_642_bfr_before (
		.din(new_net_642),
		.dout(new_net_442)
	);

	bfr new_net_643_bfr_before (
		.din(new_net_643),
		.dout(new_net_642)
	);

	bfr new_net_644_bfr_before (
		.din(new_net_644),
		.dout(new_net_643)
	);

	bfr new_net_645_bfr_before (
		.din(new_net_645),
		.dout(new_net_644)
	);

	bfr new_net_646_bfr_before (
		.din(new_net_646),
		.dout(new_net_645)
	);

	bfr new_net_647_bfr_before (
		.din(new_net_647),
		.dout(new_net_646)
	);

	bfr new_net_648_bfr_before (
		.din(new_net_648),
		.dout(new_net_647)
	);

	bfr new_net_649_bfr_before (
		.din(new_net_649),
		.dout(new_net_648)
	);

	bfr new_net_650_bfr_before (
		.din(new_net_650),
		.dout(new_net_649)
	);

	bfr new_net_651_bfr_before (
		.din(new_net_651),
		.dout(new_net_650)
	);

	bfr new_net_652_bfr_before (
		.din(new_net_652),
		.dout(new_net_651)
	);

	bfr new_net_653_bfr_before (
		.din(new_net_653),
		.dout(new_net_652)
	);

	bfr new_net_654_bfr_before (
		.din(new_net_654),
		.dout(new_net_653)
	);

	bfr new_net_655_bfr_before (
		.din(new_net_655),
		.dout(new_net_654)
	);

	bfr new_net_656_bfr_before (
		.din(new_net_656),
		.dout(new_net_655)
	);

	bfr new_net_657_bfr_before (
		.din(new_net_657),
		.dout(new_net_656)
	);

	bfr new_net_658_bfr_before (
		.din(new_net_658),
		.dout(new_net_657)
	);

	bfr new_net_659_bfr_before (
		.din(new_net_659),
		.dout(new_net_658)
	);

	bfr new_net_660_bfr_before (
		.din(new_net_660),
		.dout(new_net_659)
	);

	spl2 _087__v_fanout (
		.a(_087_),
		.b(new_net_308),
		.c(new_net_660)
	);

	bfr new_net_661_bfr_before (
		.din(new_net_661),
		.dout(new_net_443)
	);

	bfr new_net_662_bfr_before (
		.din(new_net_662),
		.dout(new_net_661)
	);

	bfr new_net_663_bfr_before (
		.din(new_net_663),
		.dout(new_net_662)
	);

	bfr new_net_664_bfr_before (
		.din(new_net_664),
		.dout(new_net_663)
	);

	bfr new_net_665_bfr_before (
		.din(new_net_665),
		.dout(new_net_664)
	);

	bfr new_net_666_bfr_before (
		.din(new_net_666),
		.dout(new_net_665)
	);

	bfr new_net_667_bfr_before (
		.din(new_net_667),
		.dout(new_net_666)
	);

	bfr new_net_668_bfr_before (
		.din(new_net_668),
		.dout(new_net_667)
	);

	bfr new_net_669_bfr_before (
		.din(new_net_669),
		.dout(new_net_668)
	);

	bfr new_net_670_bfr_before (
		.din(new_net_670),
		.dout(new_net_669)
	);

	bfr new_net_671_bfr_before (
		.din(new_net_671),
		.dout(new_net_670)
	);

	bfr new_net_672_bfr_before (
		.din(new_net_672),
		.dout(new_net_671)
	);

	bfr new_net_673_bfr_before (
		.din(new_net_673),
		.dout(new_net_672)
	);

	bfr new_net_674_bfr_before (
		.din(new_net_674),
		.dout(new_net_673)
	);

	bfr new_net_675_bfr_before (
		.din(new_net_675),
		.dout(new_net_674)
	);

	bfr new_net_676_bfr_before (
		.din(new_net_676),
		.dout(new_net_675)
	);

	spl2 _124__v_fanout (
		.a(_124_),
		.b(new_net_198),
		.c(new_net_676)
	);

	bfr new_net_677_bfr_before (
		.din(new_net_677),
		.dout(new_net_223)
	);

	bfr new_net_678_bfr_before (
		.din(new_net_678),
		.dout(new_net_677)
	);

	bfr new_net_679_bfr_before (
		.din(new_net_679),
		.dout(new_net_678)
	);

	bfr new_net_680_bfr_before (
		.din(new_net_680),
		.dout(new_net_679)
	);

	spl3L _041__v_fanout (
		.a(_041_),
		.b(new_net_225),
		.c(new_net_680),
		.d(new_net_224)
	);

	bfr new_net_681_bfr_before (
		.din(new_net_681),
		.dout(new_net_239)
	);

	bfr new_net_682_bfr_before (
		.din(new_net_682),
		.dout(new_net_681)
	);

	bfr new_net_683_bfr_before (
		.din(new_net_683),
		.dout(new_net_682)
	);

	spl2 _042__v_fanout (
		.a(_042_),
		.b(new_net_240),
		.c(new_net_683)
	);

	bfr new_net_684_bfr_before (
		.din(new_net_684),
		.dout(new_net_351)
	);

	spl2 _047__v_fanout (
		.a(_047_),
		.b(new_net_352),
		.c(new_net_684)
	);

	bfr new_net_685_bfr_before (
		.din(new_net_685),
		.dout(new_net_102)
	);

	bfr new_net_686_bfr_before (
		.din(new_net_686),
		.dout(new_net_685)
	);

	bfr new_net_687_bfr_before (
		.din(new_net_687),
		.dout(new_net_686)
	);

	bfr new_net_688_bfr_before (
		.din(new_net_688),
		.dout(new_net_687)
	);

	bfr new_net_689_bfr_before (
		.din(new_net_689),
		.dout(new_net_688)
	);

	bfr new_net_690_bfr_before (
		.din(new_net_690),
		.dout(new_net_689)
	);

	spl2 _035__v_fanout (
		.a(_035_),
		.b(new_net_103),
		.c(new_net_690)
	);

	bfr new_net_691_bfr_before (
		.din(new_net_691),
		.dout(new_net_248)
	);

	spl3L new_net_435_v_fanout (
		.a(new_net_435),
		.b(new_net_254),
		.c(new_net_250),
		.d(new_net_691)
	);

	bfr new_net_692_bfr_before (
		.din(new_net_692),
		.dout(new_net_82)
	);

	bfr new_net_693_bfr_before (
		.din(new_net_693),
		.dout(new_net_692)
	);

	bfr new_net_694_bfr_before (
		.din(new_net_694),
		.dout(new_net_693)
	);

	bfr new_net_695_bfr_before (
		.din(new_net_695),
		.dout(new_net_694)
	);

	bfr new_net_696_bfr_before (
		.din(new_net_696),
		.dout(new_net_695)
	);

	bfr new_net_697_bfr_before (
		.din(new_net_697),
		.dout(new_net_696)
	);

	bfr new_net_698_bfr_before (
		.din(new_net_698),
		.dout(new_net_697)
	);

	spl3L _034__v_fanout (
		.a(_034_),
		.b(new_net_84),
		.c(new_net_698),
		.d(new_net_83)
	);

	spl3L _049__v_fanout (
		.a(_049_),
		.b(new_net_383),
		.c(new_net_381),
		.d(new_net_382)
	);

	bfr new_net_699_bfr_before (
		.din(new_net_699),
		.dout(new_net_275)
	);

	bfr new_net_700_bfr_before (
		.din(new_net_700),
		.dout(new_net_699)
	);

	bfr new_net_701_bfr_before (
		.din(new_net_701),
		.dout(new_net_700)
	);

	bfr new_net_702_bfr_before (
		.din(new_net_702),
		.dout(new_net_701)
	);

	bfr new_net_703_bfr_before (
		.din(new_net_703),
		.dout(new_net_702)
	);

	bfr new_net_704_bfr_before (
		.din(new_net_704),
		.dout(new_net_703)
	);

	bfr new_net_705_bfr_before (
		.din(new_net_705),
		.dout(new_net_704)
	);

	bfr new_net_706_bfr_before (
		.din(new_net_706),
		.dout(new_net_705)
	);

	bfr new_net_707_bfr_before (
		.din(new_net_707),
		.dout(new_net_706)
	);

	bfr new_net_708_bfr_before (
		.din(new_net_708),
		.dout(new_net_707)
	);

	bfr new_net_709_bfr_before (
		.din(new_net_709),
		.dout(new_net_708)
	);

	bfr new_net_710_bfr_before (
		.din(new_net_710),
		.dout(new_net_709)
	);

	bfr new_net_711_bfr_before (
		.din(new_net_711),
		.dout(new_net_710)
	);

	bfr new_net_712_bfr_before (
		.din(new_net_712),
		.dout(new_net_711)
	);

	bfr new_net_713_bfr_before (
		.din(new_net_713),
		.dout(new_net_712)
	);

	bfr new_net_714_bfr_before (
		.din(new_net_714),
		.dout(new_net_713)
	);

	bfr new_net_715_bfr_before (
		.din(new_net_715),
		.dout(new_net_714)
	);

	bfr new_net_716_bfr_before (
		.din(new_net_716),
		.dout(new_net_715)
	);

	bfr new_net_717_bfr_before (
		.din(new_net_717),
		.dout(new_net_716)
	);

	bfr new_net_718_bfr_before (
		.din(new_net_718),
		.dout(new_net_717)
	);

	bfr new_net_719_bfr_before (
		.din(new_net_719),
		.dout(new_net_718)
	);

	bfr new_net_720_bfr_before (
		.din(new_net_720),
		.dout(new_net_719)
	);

	bfr new_net_721_bfr_before (
		.din(new_net_721),
		.dout(new_net_720)
	);

	spl3L _085__v_fanout (
		.a(_085_),
		.b(new_net_276),
		.c(new_net_274),
		.d(new_net_721)
	);

	bfr new_net_722_bfr_before (
		.din(new_net_722),
		.dout(new_net_290)
	);

	bfr new_net_723_bfr_before (
		.din(new_net_723),
		.dout(new_net_722)
	);

	bfr new_net_724_bfr_before (
		.din(new_net_724),
		.dout(new_net_723)
	);

	bfr new_net_725_bfr_before (
		.din(new_net_725),
		.dout(new_net_724)
	);

	bfr new_net_726_bfr_before (
		.din(new_net_726),
		.dout(new_net_725)
	);

	bfr new_net_727_bfr_before (
		.din(new_net_727),
		.dout(new_net_726)
	);

	bfr new_net_728_bfr_before (
		.din(new_net_728),
		.dout(new_net_727)
	);

	bfr new_net_729_bfr_before (
		.din(new_net_729),
		.dout(new_net_728)
	);

	bfr new_net_730_bfr_before (
		.din(new_net_730),
		.dout(new_net_729)
	);

	bfr new_net_731_bfr_before (
		.din(new_net_731),
		.dout(new_net_730)
	);

	bfr new_net_732_bfr_before (
		.din(new_net_732),
		.dout(new_net_731)
	);

	bfr new_net_733_bfr_before (
		.din(new_net_733),
		.dout(new_net_732)
	);

	bfr new_net_734_bfr_before (
		.din(new_net_734),
		.dout(new_net_733)
	);

	bfr new_net_735_bfr_before (
		.din(new_net_735),
		.dout(new_net_734)
	);

	bfr new_net_736_bfr_before (
		.din(new_net_736),
		.dout(new_net_735)
	);

	bfr new_net_737_bfr_before (
		.din(new_net_737),
		.dout(new_net_736)
	);

	bfr new_net_738_bfr_before (
		.din(new_net_738),
		.dout(new_net_737)
	);

	bfr new_net_739_bfr_before (
		.din(new_net_739),
		.dout(new_net_738)
	);

	bfr new_net_740_bfr_before (
		.din(new_net_740),
		.dout(new_net_739)
	);

	bfr new_net_741_bfr_before (
		.din(new_net_741),
		.dout(new_net_740)
	);

	bfr new_net_742_bfr_before (
		.din(new_net_742),
		.dout(new_net_741)
	);

	bfr new_net_743_bfr_before (
		.din(new_net_743),
		.dout(new_net_742)
	);

	spl2 _086__v_fanout (
		.a(_086_),
		.b(new_net_743),
		.c(new_net_289)
	);

	spl4L new_net_434_v_fanout (
		.a(new_net_434),
		.b(new_net_251),
		.c(new_net_253),
		.d(new_net_435),
		.e(new_net_252)
	);

	bfr new_net_744_bfr_before (
		.din(new_net_744),
		.dout(new_net_218)
	);

	bfr new_net_745_bfr_before (
		.din(new_net_745),
		.dout(new_net_744)
	);

	bfr new_net_746_bfr_before (
		.din(new_net_746),
		.dout(new_net_745)
	);

	bfr new_net_747_bfr_before (
		.din(new_net_747),
		.dout(new_net_746)
	);

	bfr new_net_748_bfr_before (
		.din(new_net_748),
		.dout(new_net_747)
	);

	bfr new_net_749_bfr_before (
		.din(new_net_749),
		.dout(new_net_748)
	);

	bfr new_net_750_bfr_before (
		.din(new_net_750),
		.dout(new_net_749)
	);

	bfr new_net_751_bfr_before (
		.din(new_net_751),
		.dout(new_net_750)
	);

	bfr new_net_752_bfr_before (
		.din(new_net_752),
		.dout(new_net_751)
	);

	bfr new_net_753_bfr_before (
		.din(new_net_753),
		.dout(new_net_752)
	);

	bfr new_net_754_bfr_before (
		.din(new_net_754),
		.dout(new_net_753)
	);

	bfr new_net_755_bfr_before (
		.din(new_net_755),
		.dout(new_net_754)
	);

	bfr new_net_756_bfr_before (
		.din(new_net_756),
		.dout(new_net_755)
	);

	bfr new_net_757_bfr_before (
		.din(new_net_757),
		.dout(new_net_756)
	);

	bfr new_net_758_bfr_before (
		.din(new_net_758),
		.dout(new_net_757)
	);

	bfr new_net_759_bfr_before (
		.din(new_net_759),
		.dout(new_net_758)
	);

	spl2 _103__v_fanout (
		.a(_103_),
		.b(new_net_219),
		.c(new_net_759)
	);

	bfr new_net_760_bfr_before (
		.din(new_net_760),
		.dout(new_net_176)
	);

	bfr new_net_761_bfr_before (
		.din(new_net_761),
		.dout(new_net_760)
	);

	bfr new_net_762_bfr_before (
		.din(new_net_762),
		.dout(new_net_761)
	);

	bfr new_net_763_bfr_before (
		.din(new_net_763),
		.dout(new_net_762)
	);

	bfr new_net_764_bfr_before (
		.din(new_net_764),
		.dout(new_net_763)
	);

	bfr new_net_765_bfr_before (
		.din(new_net_765),
		.dout(new_net_764)
	);

	bfr new_net_766_bfr_before (
		.din(new_net_766),
		.dout(new_net_765)
	);

	bfr new_net_767_bfr_before (
		.din(new_net_767),
		.dout(new_net_766)
	);

	bfr new_net_768_bfr_before (
		.din(new_net_768),
		.dout(new_net_767)
	);

	bfr new_net_769_bfr_before (
		.din(new_net_769),
		.dout(new_net_768)
	);

	bfr new_net_770_bfr_before (
		.din(new_net_770),
		.dout(new_net_769)
	);

	bfr new_net_771_bfr_before (
		.din(new_net_771),
		.dout(new_net_770)
	);

	bfr new_net_772_bfr_before (
		.din(new_net_772),
		.dout(new_net_771)
	);

	bfr new_net_773_bfr_before (
		.din(new_net_773),
		.dout(new_net_772)
	);

	bfr new_net_774_bfr_before (
		.din(new_net_774),
		.dout(new_net_773)
	);

	bfr new_net_775_bfr_before (
		.din(new_net_775),
		.dout(new_net_774)
	);

	bfr new_net_776_bfr_before (
		.din(new_net_776),
		.dout(new_net_775)
	);

	spl3L _102__v_fanout (
		.a(_102_),
		.b(new_net_177),
		.c(new_net_776),
		.d(new_net_178)
	);

	spl3L _027__v_fanout (
		.a(_027_),
		.b(new_net_374),
		.c(new_net_372),
		.d(new_net_373)
	);

	bfr new_net_777_bfr_before (
		.din(new_net_777),
		.dout(new_net_63)
	);

	bfr new_net_778_bfr_before (
		.din(new_net_778),
		.dout(new_net_777)
	);

	bfr new_net_779_bfr_before (
		.din(new_net_779),
		.dout(new_net_778)
	);

	bfr new_net_780_bfr_before (
		.din(new_net_780),
		.dout(new_net_779)
	);

	bfr new_net_781_bfr_before (
		.din(new_net_781),
		.dout(new_net_780)
	);

	bfr new_net_782_bfr_before (
		.din(new_net_782),
		.dout(new_net_781)
	);

	bfr new_net_783_bfr_before (
		.din(new_net_783),
		.dout(new_net_782)
	);

	bfr new_net_784_bfr_before (
		.din(new_net_784),
		.dout(new_net_783)
	);

	bfr new_net_785_bfr_before (
		.din(new_net_785),
		.dout(new_net_784)
	);

	bfr new_net_786_bfr_before (
		.din(new_net_786),
		.dout(new_net_785)
	);

	bfr new_net_787_bfr_before (
		.din(new_net_787),
		.dout(new_net_786)
	);

	bfr new_net_788_bfr_before (
		.din(new_net_788),
		.dout(new_net_787)
	);

	bfr new_net_789_bfr_before (
		.din(new_net_789),
		.dout(new_net_788)
	);

	bfr new_net_790_bfr_before (
		.din(new_net_790),
		.dout(new_net_789)
	);

	bfr new_net_791_bfr_before (
		.din(new_net_791),
		.dout(new_net_790)
	);

	bfr new_net_792_bfr_before (
		.din(new_net_792),
		.dout(new_net_791)
	);

	bfr new_net_793_bfr_before (
		.din(new_net_793),
		.dout(new_net_792)
	);

	bfr new_net_794_bfr_before (
		.din(new_net_794),
		.dout(new_net_793)
	);

	bfr new_net_795_bfr_before (
		.din(new_net_795),
		.dout(new_net_794)
	);

	spl2 _095__v_fanout (
		.a(_095_),
		.b(new_net_64),
		.c(new_net_795)
	);

	spl2 new_net_413_v_fanout (
		.a(new_net_413),
		.b(new_net_132),
		.c(new_net_134)
	);

	bfr new_net_796_bfr_before (
		.din(new_net_796),
		.dout(new_net_41)
	);

	bfr new_net_797_bfr_before (
		.din(new_net_797),
		.dout(new_net_796)
	);

	bfr new_net_798_bfr_before (
		.din(new_net_798),
		.dout(new_net_797)
	);

	bfr new_net_799_bfr_before (
		.din(new_net_799),
		.dout(new_net_798)
	);

	bfr new_net_800_bfr_before (
		.din(new_net_800),
		.dout(new_net_799)
	);

	bfr new_net_801_bfr_before (
		.din(new_net_801),
		.dout(new_net_800)
	);

	bfr new_net_802_bfr_before (
		.din(new_net_802),
		.dout(new_net_801)
	);

	bfr new_net_803_bfr_before (
		.din(new_net_803),
		.dout(new_net_802)
	);

	bfr new_net_804_bfr_before (
		.din(new_net_804),
		.dout(new_net_803)
	);

	bfr new_net_805_bfr_before (
		.din(new_net_805),
		.dout(new_net_804)
	);

	bfr new_net_806_bfr_before (
		.din(new_net_806),
		.dout(new_net_805)
	);

	bfr new_net_807_bfr_before (
		.din(new_net_807),
		.dout(new_net_806)
	);

	bfr new_net_808_bfr_before (
		.din(new_net_808),
		.dout(new_net_807)
	);

	bfr new_net_809_bfr_before (
		.din(new_net_809),
		.dout(new_net_808)
	);

	bfr new_net_810_bfr_before (
		.din(new_net_810),
		.dout(new_net_809)
	);

	bfr new_net_811_bfr_before (
		.din(new_net_811),
		.dout(new_net_810)
	);

	bfr new_net_812_bfr_before (
		.din(new_net_812),
		.dout(new_net_811)
	);

	bfr new_net_813_bfr_before (
		.din(new_net_813),
		.dout(new_net_812)
	);

	bfr new_net_814_bfr_before (
		.din(new_net_814),
		.dout(new_net_813)
	);

	bfr new_net_815_bfr_before (
		.din(new_net_815),
		.dout(new_net_814)
	);

	spl3L _094__v_fanout (
		.a(_094_),
		.b(new_net_42),
		.c(new_net_815),
		.d(new_net_43)
	);

	bfr new_net_816_bfr_before (
		.din(new_net_816),
		.dout(new_net_185)
	);

	bfr new_net_817_bfr_before (
		.din(new_net_817),
		.dout(new_net_816)
	);

	bfr new_net_818_bfr_before (
		.din(new_net_818),
		.dout(new_net_817)
	);

	bfr new_net_819_bfr_before (
		.din(new_net_819),
		.dout(new_net_818)
	);

	bfr new_net_820_bfr_before (
		.din(new_net_820),
		.dout(new_net_819)
	);

	bfr new_net_821_bfr_before (
		.din(new_net_821),
		.dout(new_net_820)
	);

	bfr new_net_822_bfr_before (
		.din(new_net_822),
		.dout(new_net_821)
	);

	bfr new_net_823_bfr_before (
		.din(new_net_823),
		.dout(new_net_822)
	);

	bfr new_net_824_bfr_before (
		.din(new_net_824),
		.dout(new_net_823)
	);

	bfr new_net_825_bfr_before (
		.din(new_net_825),
		.dout(new_net_824)
	);

	bfr new_net_826_bfr_before (
		.din(new_net_826),
		.dout(new_net_825)
	);

	bfr new_net_827_bfr_before (
		.din(new_net_827),
		.dout(new_net_826)
	);

	bfr new_net_828_bfr_before (
		.din(new_net_828),
		.dout(new_net_827)
	);

	bfr new_net_829_bfr_before (
		.din(new_net_829),
		.dout(new_net_828)
	);

	spl3L _018__v_fanout (
		.a(_018_),
		.b(new_net_829),
		.c(new_net_184),
		.d(new_net_186)
	);

	bfr new_net_830_bfr_before (
		.din(new_net_830),
		.dout(new_net_165)
	);

	bfr new_net_831_bfr_before (
		.din(new_net_831),
		.dout(new_net_830)
	);

	bfr new_net_832_bfr_before (
		.din(new_net_832),
		.dout(new_net_831)
	);

	bfr new_net_833_bfr_before (
		.din(new_net_833),
		.dout(new_net_832)
	);

	bfr new_net_834_bfr_before (
		.din(new_net_834),
		.dout(new_net_833)
	);

	bfr new_net_835_bfr_before (
		.din(new_net_835),
		.dout(new_net_834)
	);

	bfr new_net_836_bfr_before (
		.din(new_net_836),
		.dout(new_net_835)
	);

	bfr new_net_837_bfr_before (
		.din(new_net_837),
		.dout(new_net_836)
	);

	bfr new_net_838_bfr_before (
		.din(new_net_838),
		.dout(new_net_837)
	);

	bfr new_net_839_bfr_before (
		.din(new_net_839),
		.dout(new_net_838)
	);

	bfr new_net_840_bfr_before (
		.din(new_net_840),
		.dout(new_net_839)
	);

	bfr new_net_841_bfr_before (
		.din(new_net_841),
		.dout(new_net_840)
	);

	bfr new_net_842_bfr_before (
		.din(new_net_842),
		.dout(new_net_841)
	);

	spl2 _017__v_fanout (
		.a(_017_),
		.b(new_net_842),
		.c(new_net_164)
	);

	spl3L _040__v_fanout (
		.a(_040_),
		.b(new_net_191),
		.c(new_net_189),
		.d(new_net_190)
	);

	spl2 new_net_417_v_fanout (
		.a(new_net_417),
		.b(new_net_180),
		.c(new_net_179)
	);

	spl2 new_net_415_v_fanout (
		.a(new_net_415),
		.b(new_net_153),
		.c(new_net_154)
	);

	spl3L _046__v_fanout (
		.a(_046_),
		.b(new_net_327),
		.c(new_net_325),
		.d(new_net_326)
	);

	bfr new_net_843_bfr_before (
		.din(new_net_843),
		.dout(new_net_323)
	);

	spl4L new_net_427_v_fanout (
		.a(new_net_427),
		.b(new_net_324),
		.c(new_net_320),
		.d(new_net_843),
		.e(new_net_321)
	);

	spl3L _033__v_fanout (
		.a(_033_),
		.b(new_net_68),
		.c(new_net_67),
		.d(new_net_69)
	);

	spl2 new_net_409_v_fanout (
		.a(new_net_409),
		.b(new_net_94),
		.c(new_net_91)
	);

	spl3L _101__v_fanout (
		.a(_101_),
		.b(new_net_163),
		.c(new_net_161),
		.d(new_net_162)
	);

	spl2 new_net_405_v_fanout (
		.a(new_net_405),
		.b(new_net_60),
		.c(new_net_56)
	);

	spl3L _093__v_fanout (
		.a(_093_),
		.b(new_net_21),
		.c(new_net_19),
		.d(new_net_20)
	);

	spl2 new_net_411_v_fanout (
		.a(new_net_411),
		.b(new_net_115),
		.c(new_net_111)
	);

	spl2 new_net_403_v_fanout (
		.a(new_net_403),
		.b(new_net_38),
		.c(new_net_39)
	);

	spl4L new_net_426_v_fanout (
		.a(new_net_426),
		.b(new_net_322),
		.c(new_net_318),
		.d(new_net_427),
		.e(new_net_319)
	);

	spl3L _016__v_fanout (
		.a(_016_),
		.b(new_net_151),
		.c(new_net_149),
		.d(new_net_150)
	);

	spl3L _084__v_fanout (
		.a(_084_),
		.b(new_net_242),
		.c(new_net_241),
		.d(new_net_243)
	);

	spl4L _024__v_fanout (
		.a(_024_),
		.b(new_net_315),
		.c(new_net_316),
		.d(new_net_314),
		.e(new_net_313)
	);

	spl4L new_net_440_v_fanout (
		.a(new_net_440),
		.b(new_net_292),
		.c(new_net_295),
		.d(new_net_293),
		.e(new_net_291)
	);

	spl2 _241__v_fanout (
		.a(_241_),
		.b(new_net_33),
		.c(new_net_32)
	);

	bfr new_net_844_bfr_after (
		.din(_021_),
		.dout(new_net_844)
	);

	bfr new_net_845_bfr_before (
		.din(new_net_845),
		.dout(new_net_255)
	);

	bfr new_net_846_bfr_before (
		.din(new_net_846),
		.dout(new_net_845)
	);

	spl4L _021__v_fanout (
		.a(new_net_844),
		.b(new_net_256),
		.c(new_net_257),
		.d(new_net_258),
		.e(new_net_846)
	);

	spl4L new_net_441_v_fanout (
		.a(new_net_441),
		.b(new_net_298),
		.c(new_net_297),
		.d(new_net_296),
		.e(new_net_294)
	);

	spl2 _267__v_fanout (
		.a(_267_),
		.b(new_net_137),
		.c(new_net_136)
	);

	spl4L _005__v_fanout (
		.a(_005_),
		.b(new_net_350),
		.c(new_net_348),
		.d(new_net_349),
		.e(new_net_347)
	);

	spl2 _002__v_fanout (
		.a(_002_),
		.b(new_net_441),
		.c(new_net_440)
	);

	spl4L _013__v_fanout (
		.a(_013_),
		.b(new_net_98),
		.c(new_net_99),
		.d(new_net_97),
		.e(new_net_96)
	);

	spl4L new_net_439_v_fanout (
		.a(new_net_439),
		.b(new_net_11),
		.c(new_net_12),
		.d(new_net_13),
		.e(new_net_9)
	);

	spl4L new_net_438_v_fanout (
		.a(new_net_438),
		.b(new_net_8),
		.c(new_net_10),
		.d(new_net_7),
		.e(new_net_6)
	);

	bfr new_net_847_bfr_before (
		.din(new_net_847),
		.dout(new_net_409)
	);

	bfr new_net_848_bfr_before (
		.din(new_net_848),
		.dout(new_net_847)
	);

	bfr new_net_849_bfr_before (
		.din(new_net_849),
		.dout(new_net_848)
	);

	bfr new_net_850_bfr_before (
		.din(new_net_850),
		.dout(new_net_849)
	);

	spl2 new_net_408_v_fanout (
		.a(new_net_408),
		.b(new_net_850),
		.c(new_net_93)
	);

	bfr new_net_851_bfr_before (
		.din(new_net_851),
		.dout(new_net_413)
	);

	bfr new_net_852_bfr_before (
		.din(new_net_852),
		.dout(new_net_851)
	);

	bfr new_net_853_bfr_before (
		.din(new_net_853),
		.dout(new_net_852)
	);

	bfr new_net_854_bfr_before (
		.din(new_net_854),
		.dout(new_net_853)
	);

	bfr new_net_855_bfr_before (
		.din(new_net_855),
		.dout(new_net_854)
	);

	bfr new_net_856_bfr_before (
		.din(new_net_856),
		.dout(new_net_855)
	);

	spl2 new_net_412_v_fanout (
		.a(new_net_412),
		.b(new_net_856),
		.c(new_net_131)
	);

	spl2 _072__v_fanout (
		.a(_072_),
		.b(new_net_439),
		.c(new_net_438)
	);

	spl2 _238__v_fanout (
		.a(_238_),
		.b(new_net_388),
		.c(new_net_387)
	);

	bfr new_net_857_bfr_before (
		.din(new_net_857),
		.dout(new_net_403)
	);

	bfr new_net_858_bfr_before (
		.din(new_net_858),
		.dout(new_net_857)
	);

	bfr new_net_859_bfr_before (
		.din(new_net_859),
		.dout(new_net_858)
	);

	bfr new_net_860_bfr_before (
		.din(new_net_860),
		.dout(new_net_859)
	);

	spl2 new_net_402_v_fanout (
		.a(new_net_402),
		.b(new_net_860),
		.c(new_net_37)
	);

	spl2 _011__v_fanout (
		.a(_011_),
		.b(new_net_52),
		.c(new_net_51)
	);

	spl2 _229__v_fanout (
		.a(_229_),
		.b(new_net_215),
		.c(new_net_214)
	);

	bfr new_net_861_bfr_before (
		.din(new_net_861),
		.dout(new_net_417)
	);

	bfr new_net_862_bfr_before (
		.din(new_net_862),
		.dout(new_net_861)
	);

	bfr new_net_863_bfr_before (
		.din(new_net_863),
		.dout(new_net_862)
	);

	bfr new_net_864_bfr_before (
		.din(new_net_864),
		.dout(new_net_863)
	);

	bfr new_net_865_bfr_before (
		.din(new_net_865),
		.dout(new_net_864)
	);

	spl2 new_net_416_v_fanout (
		.a(new_net_416),
		.b(new_net_865),
		.c(new_net_182)
	);

	bfr new_net_866_bfr_after (
		.din(_223_),
		.dout(new_net_866)
	);

	bfr new_net_867_bfr_after (
		.din(new_net_866),
		.dout(new_net_867)
	);

	bfr new_net_868_bfr_after (
		.din(new_net_867),
		.dout(new_net_868)
	);

	spl2 _223__v_fanout (
		.a(new_net_868),
		.b(new_net_101),
		.c(new_net_100)
	);

	bfr new_net_869_bfr_before (
		.din(new_net_869),
		.dout(new_net_415)
	);

	bfr new_net_870_bfr_before (
		.din(new_net_870),
		.dout(new_net_869)
	);

	bfr new_net_871_bfr_before (
		.din(new_net_871),
		.dout(new_net_870)
	);

	bfr new_net_872_bfr_before (
		.din(new_net_872),
		.dout(new_net_871)
	);

	bfr new_net_873_bfr_before (
		.din(new_net_873),
		.dout(new_net_872)
	);

	spl2 new_net_414_v_fanout (
		.a(new_net_414),
		.b(new_net_873),
		.c(new_net_155)
	);

	bfr new_net_874_bfr_before (
		.din(new_net_874),
		.dout(new_net_331)
	);

	spl2 _004__v_fanout (
		.a(_004_),
		.b(new_net_874),
		.c(new_net_330)
	);

	bfr new_net_875_bfr_before (
		.din(new_net_875),
		.dout(new_net_405)
	);

	bfr new_net_876_bfr_before (
		.din(new_net_876),
		.dout(new_net_875)
	);

	bfr new_net_877_bfr_before (
		.din(new_net_877),
		.dout(new_net_876)
	);

	bfr new_net_878_bfr_before (
		.din(new_net_878),
		.dout(new_net_877)
	);

	spl2 new_net_404_v_fanout (
		.a(new_net_404),
		.b(new_net_878),
		.c(new_net_59)
	);

	spl2 _255__v_fanout (
		.a(_255_),
		.b(new_net_305),
		.c(new_net_304)
	);

	bfr new_net_879_bfr_before (
		.din(new_net_879),
		.dout(new_net_411)
	);

	bfr new_net_880_bfr_before (
		.din(new_net_880),
		.dout(new_net_879)
	);

	bfr new_net_881_bfr_before (
		.din(new_net_881),
		.dout(new_net_880)
	);

	bfr new_net_882_bfr_before (
		.din(new_net_882),
		.dout(new_net_881)
	);

	spl2 new_net_410_v_fanout (
		.a(new_net_410),
		.b(new_net_882),
		.c(new_net_112)
	);

	spl2 new_net_431_v_fanout (
		.a(new_net_431),
		.b(new_net_26),
		.c(new_net_24)
	);

	spl2 _264__v_fanout (
		.a(_264_),
		.b(new_net_81),
		.c(new_net_80)
	);

	bfr new_net_883_bfr_after (
		.din(_249_),
		.dout(new_net_883)
	);

	bfr new_net_884_bfr_after (
		.din(new_net_883),
		.dout(new_net_884)
	);

	bfr new_net_885_bfr_after (
		.din(new_net_884),
		.dout(new_net_885)
	);

	spl2 _249__v_fanout (
		.a(new_net_885),
		.b(new_net_175),
		.c(new_net_174)
	);

	spl2 _272__v_fanout (
		.a(_272_),
		.b(new_net_238),
		.c(new_net_237)
	);

	spl4L _278__v_fanout (
		.a(_278_),
		.b(new_net_359),
		.c(new_net_358),
		.d(new_net_357),
		.e(new_net_356)
	);

	bfr new_net_886_bfr_after (
		.din(new_net_0),
		.dout(new_net_886)
	);

	bfr new_net_887_bfr_before (
		.din(new_net_887),
		.dout(N390)
	);

	bfr new_net_888_bfr_before (
		.din(new_net_888),
		.dout(new_net_887)
	);

	bfr new_net_889_bfr_before (
		.din(new_net_889),
		.dout(new_net_888)
	);

	bfr new_net_890_bfr_before (
		.din(new_net_890),
		.dout(new_net_889)
	);

	bfr new_net_891_bfr_before (
		.din(new_net_891),
		.dout(new_net_890)
	);

	bfr new_net_892_bfr_before (
		.din(new_net_892),
		.dout(new_net_891)
	);

	bfr new_net_893_bfr_before (
		.din(new_net_893),
		.dout(new_net_892)
	);

	bfr new_net_894_bfr_before (
		.din(new_net_894),
		.dout(new_net_893)
	);

	bfr new_net_895_bfr_before (
		.din(new_net_895),
		.dout(new_net_894)
	);

	bfr new_net_896_bfr_before (
		.din(new_net_896),
		.dout(new_net_895)
	);

	bfr new_net_897_bfr_before (
		.din(new_net_897),
		.dout(new_net_896)
	);

	bfr new_net_898_bfr_before (
		.din(new_net_898),
		.dout(new_net_897)
	);

	bfr new_net_899_bfr_before (
		.din(new_net_899),
		.dout(new_net_898)
	);

	bfr new_net_900_bfr_before (
		.din(new_net_900),
		.dout(new_net_899)
	);

	bfr new_net_901_bfr_before (
		.din(new_net_901),
		.dout(new_net_900)
	);

	bfr new_net_902_bfr_before (
		.din(new_net_902),
		.dout(new_net_901)
	);

	bfr new_net_903_bfr_before (
		.din(new_net_903),
		.dout(new_net_902)
	);

	bfr new_net_904_bfr_before (
		.din(new_net_904),
		.dout(new_net_903)
	);

	bfr new_net_905_bfr_before (
		.din(new_net_905),
		.dout(new_net_904)
	);

	bfr new_net_906_bfr_before (
		.din(new_net_906),
		.dout(new_net_905)
	);

	bfr new_net_907_bfr_before (
		.din(new_net_907),
		.dout(new_net_906)
	);

	bfr new_net_908_bfr_before (
		.din(new_net_908),
		.dout(new_net_907)
	);

	bfr new_net_909_bfr_before (
		.din(new_net_909),
		.dout(new_net_908)
	);

	bfr new_net_910_bfr_before (
		.din(new_net_910),
		.dout(new_net_909)
	);

	bfr new_net_911_bfr_before (
		.din(new_net_911),
		.dout(new_net_910)
	);

	bfr new_net_912_bfr_before (
		.din(new_net_912),
		.dout(new_net_911)
	);

	bfr new_net_913_bfr_before (
		.din(new_net_913),
		.dout(new_net_912)
	);

	bfr new_net_914_bfr_before (
		.din(new_net_914),
		.dout(new_net_913)
	);

	bfr new_net_915_bfr_before (
		.din(new_net_915),
		.dout(new_net_914)
	);

	bfr new_net_916_bfr_before (
		.din(new_net_916),
		.dout(new_net_915)
	);

	bfr new_net_917_bfr_before (
		.din(new_net_917),
		.dout(new_net_916)
	);

	bfr new_net_918_bfr_before (
		.din(new_net_918),
		.dout(new_net_917)
	);

	bfr new_net_919_bfr_before (
		.din(new_net_919),
		.dout(new_net_918)
	);

	bfr new_net_920_bfr_before (
		.din(new_net_920),
		.dout(new_net_919)
	);

	bfr new_net_921_bfr_before (
		.din(new_net_921),
		.dout(new_net_920)
	);

	spl3L new_net_0_v_fanout (
		.a(new_net_886),
		.b(new_net_221),
		.c(new_net_921),
		.d(new_net_222)
	);

	spl3L _067__v_fanout (
		.a(_067_),
		.b(new_net_333),
		.c(new_net_332),
		.d(new_net_334)
	);

	spl2 _226__v_fanout (
		.a(_226_),
		.b(new_net_148),
		.c(new_net_147)
	);

	spl2 new_net_401_v_fanout (
		.a(new_net_401),
		.b(new_net_272),
		.c(new_net_270)
	);

	spl2 _271__v_fanout (
		.a(_271_),
		.b(new_net_209),
		.c(new_net_208)
	);

	spl2 _252__v_fanout (
		.a(_252_),
		.b(new_net_245),
		.c(new_net_244)
	);

	spl2 _258__v_fanout (
		.a(_258_),
		.b(new_net_363),
		.c(new_net_362)
	);

	spl2 _235__v_fanout (
		.a(_235_),
		.b(new_net_339),
		.c(new_net_338)
	);

	spl2 _246__v_fanout (
		.a(_246_),
		.b(new_net_126),
		.c(new_net_125)
	);

	spl2 _261__v_fanout (
		.a(_261_),
		.b(new_net_23),
		.c(new_net_22)
	);

	spl2 _220__v_fanout (
		.a(_220_),
		.b(new_net_35),
		.c(new_net_34)
	);

	bfr new_net_922_bfr_before (
		.din(new_net_922),
		.dout(new_net_104)
	);

	bfr new_net_923_bfr_before (
		.din(new_net_923),
		.dout(new_net_922)
	);

	bfr new_net_924_bfr_before (
		.din(new_net_924),
		.dout(new_net_923)
	);

	bfr new_net_925_bfr_before (
		.din(new_net_925),
		.dout(new_net_924)
	);

	bfr new_net_926_bfr_before (
		.din(new_net_926),
		.dout(new_net_925)
	);

	bfr new_net_927_bfr_before (
		.din(new_net_927),
		.dout(new_net_926)
	);

	spl3L new_net_432_v_fanout (
		.a(new_net_432),
		.b(new_net_927),
		.c(new_net_105),
		.d(new_net_107)
	);

	spl2 _232__v_fanout (
		.a(_232_),
		.b(new_net_278),
		.c(new_net_277)
	);

	spl2 _216__v_fanout (
		.a(_216_),
		.b(new_net_367),
		.c(new_net_366)
	);

	bfr new_net_928_bfr_after (
		.din(_036_),
		.dout(new_net_928)
	);

	bfr new_net_929_bfr_after (
		.din(new_net_928),
		.dout(new_net_929)
	);

	bfr new_net_930_bfr_after (
		.din(new_net_929),
		.dout(new_net_930)
	);

	bfr new_net_931_bfr_after (
		.din(new_net_930),
		.dout(new_net_931)
	);

	bfr new_net_932_bfr_after (
		.din(new_net_931),
		.dout(new_net_932)
	);

	bfr new_net_933_bfr_after (
		.din(new_net_932),
		.dout(new_net_933)
	);

	bfr new_net_934_bfr_after (
		.din(new_net_933),
		.dout(new_net_934)
	);

	bfr new_net_935_bfr_after (
		.din(new_net_934),
		.dout(new_net_935)
	);

	bfr new_net_936_bfr_after (
		.din(new_net_935),
		.dout(new_net_936)
	);

	bfr new_net_937_bfr_after (
		.din(new_net_936),
		.dout(new_net_937)
	);

	bfr new_net_938_bfr_after (
		.din(new_net_937),
		.dout(new_net_938)
	);

	spl2 _036__v_fanout (
		.a(new_net_938),
		.b(new_net_124),
		.c(new_net_123)
	);

	bfr new_net_939_bfr_before (
		.din(new_net_939),
		.dout(new_net_344)
	);

	spl2 _277__v_fanout (
		.a(_277_),
		.b(new_net_939),
		.c(new_net_343)
	);

	spl2 _068__v_fanout (
		.a(_068_),
		.b(new_net_361),
		.c(new_net_360)
	);

	spl2 _283__v_fanout (
		.a(_283_),
		.b(new_net_28),
		.c(new_net_27)
	);

	bfr new_net_940_bfr_after (
		.din(_279_),
		.dout(new_net_940)
	);

	bfr new_net_941_bfr_after (
		.din(new_net_940),
		.dout(new_net_941)
	);

	spl2 _279__v_fanout (
		.a(new_net_941),
		.b(new_net_371),
		.c(new_net_370)
	);

	spl2 _009__v_fanout (
		.a(_009_),
		.b(new_net_15),
		.c(new_net_14)
	);

	spl2 _282__v_fanout (
		.a(_282_),
		.b(new_net_2),
		.c(new_net_1)
	);

	spl2 _217__v_fanout (
		.a(_217_),
		.b(new_net_380),
		.c(new_net_379)
	);

	spl2 new_net_429_v_fanout (
		.a(new_net_429),
		.b(new_net_205),
		.c(new_net_206)
	);

	spl3L _008__v_fanout (
		.a(_008_),
		.b(new_net_396),
		.c(new_net_394),
		.d(new_net_395)
	);

	bfr new_net_942_bfr_after (
		.din(_063_),
		.dout(new_net_942)
	);

	bfr new_net_943_bfr_after (
		.din(new_net_942),
		.dout(new_net_943)
	);

	bfr new_net_944_bfr_after (
		.din(new_net_943),
		.dout(new_net_944)
	);

	bfr new_net_945_bfr_after (
		.din(new_net_944),
		.dout(new_net_945)
	);

	bfr new_net_946_bfr_after (
		.din(new_net_945),
		.dout(new_net_946)
	);

	bfr new_net_947_bfr_after (
		.din(new_net_946),
		.dout(new_net_947)
	);

	bfr new_net_948_bfr_after (
		.din(new_net_947),
		.dout(new_net_948)
	);

	bfr new_net_949_bfr_after (
		.din(new_net_948),
		.dout(new_net_949)
	);

	bfr new_net_950_bfr_after (
		.din(new_net_949),
		.dout(new_net_950)
	);

	bfr new_net_951_bfr_after (
		.din(new_net_950),
		.dout(new_net_951)
	);

	bfr new_net_952_bfr_after (
		.din(new_net_951),
		.dout(new_net_952)
	);

	bfr new_net_953_bfr_before (
		.din(new_net_953),
		.dout(new_net_249)
	);

	spl2 _063__v_fanout (
		.a(new_net_952),
		.b(new_net_434),
		.c(new_net_953)
	);

	bfr new_net_954_bfr_before (
		.din(new_net_954),
		.dout(new_net_86)
	);

	spl3L _286__v_fanout (
		.a(_286_),
		.b(new_net_87),
		.c(new_net_85),
		.d(new_net_954)
	);

	bfr new_net_955_bfr_after (
		.din(_048_),
		.dout(new_net_955)
	);

	bfr new_net_956_bfr_after (
		.din(new_net_955),
		.dout(new_net_956)
	);

	bfr new_net_957_bfr_after (
		.din(new_net_956),
		.dout(new_net_957)
	);

	bfr new_net_958_bfr_after (
		.din(new_net_957),
		.dout(new_net_958)
	);

	bfr new_net_959_bfr_after (
		.din(new_net_958),
		.dout(new_net_959)
	);

	bfr new_net_960_bfr_after (
		.din(new_net_959),
		.dout(new_net_960)
	);

	bfr new_net_961_bfr_after (
		.din(new_net_960),
		.dout(new_net_961)
	);

	bfr new_net_962_bfr_after (
		.din(new_net_961),
		.dout(new_net_962)
	);

	bfr new_net_963_bfr_after (
		.din(new_net_962),
		.dout(new_net_963)
	);

	bfr new_net_964_bfr_after (
		.din(new_net_963),
		.dout(new_net_964)
	);

	bfr new_net_965_bfr_after (
		.din(new_net_964),
		.dout(new_net_965)
	);

	bfr new_net_966_bfr_after (
		.din(new_net_965),
		.dout(new_net_966)
	);

	bfr new_net_967_bfr_after (
		.din(new_net_966),
		.dout(new_net_967)
	);

	bfr new_net_968_bfr_before (
		.din(new_net_968),
		.dout(new_net_365)
	);

	bfr new_net_969_bfr_before (
		.din(new_net_969),
		.dout(new_net_968)
	);

	spl2 _048__v_fanout (
		.a(new_net_967),
		.b(new_net_969),
		.c(new_net_364)
	);

	bfr new_net_970_bfr_after (
		.din(_111_),
		.dout(new_net_970)
	);

	bfr new_net_971_bfr_after (
		.din(new_net_970),
		.dout(new_net_971)
	);

	bfr new_net_972_bfr_after (
		.din(new_net_971),
		.dout(new_net_972)
	);

	bfr new_net_973_bfr_after (
		.din(new_net_972),
		.dout(new_net_973)
	);

	bfr new_net_974_bfr_after (
		.din(new_net_973),
		.dout(new_net_974)
	);

	bfr new_net_975_bfr_after (
		.din(new_net_974),
		.dout(new_net_975)
	);

	bfr new_net_976_bfr_after (
		.din(new_net_975),
		.dout(new_net_976)
	);

	bfr new_net_977_bfr_after (
		.din(new_net_976),
		.dout(new_net_977)
	);

	bfr new_net_978_bfr_after (
		.din(new_net_977),
		.dout(new_net_978)
	);

	bfr new_net_979_bfr_after (
		.din(new_net_978),
		.dout(new_net_979)
	);

	bfr new_net_980_bfr_after (
		.din(new_net_979),
		.dout(new_net_980)
	);

	bfr new_net_981_bfr_after (
		.din(new_net_980),
		.dout(new_net_981)
	);

	bfr new_net_982_bfr_after (
		.din(new_net_981),
		.dout(new_net_982)
	);

	bfr new_net_983_bfr_after (
		.din(new_net_982),
		.dout(new_net_983)
	);

	bfr new_net_984_bfr_after (
		.din(new_net_983),
		.dout(new_net_984)
	);

	bfr new_net_985_bfr_after (
		.din(new_net_984),
		.dout(new_net_985)
	);

	bfr new_net_986_bfr_before (
		.din(new_net_986),
		.dout(new_net_436)
	);

	bfr new_net_987_bfr_before (
		.din(new_net_987),
		.dout(new_net_986)
	);

	bfr new_net_988_bfr_before (
		.din(new_net_988),
		.dout(new_net_987)
	);

	bfr new_net_989_bfr_before (
		.din(new_net_989),
		.dout(new_net_988)
	);

	bfr new_net_990_bfr_before (
		.din(new_net_990),
		.dout(new_net_989)
	);

	bfr new_net_991_bfr_before (
		.din(new_net_991),
		.dout(new_net_990)
	);

	bfr new_net_992_bfr_before (
		.din(new_net_992),
		.dout(new_net_991)
	);

	bfr new_net_993_bfr_before (
		.din(new_net_993),
		.dout(new_net_992)
	);

	bfr new_net_994_bfr_before (
		.din(new_net_994),
		.dout(new_net_993)
	);

	bfr new_net_995_bfr_before (
		.din(new_net_995),
		.dout(new_net_994)
	);

	bfr new_net_996_bfr_before (
		.din(new_net_996),
		.dout(new_net_995)
	);

	bfr new_net_997_bfr_before (
		.din(new_net_997),
		.dout(new_net_996)
	);

	spl2 _111__v_fanout (
		.a(new_net_985),
		.b(new_net_376),
		.c(new_net_997)
	);

	spl3L new_net_428_v_fanout (
		.a(new_net_428),
		.b(new_net_207),
		.c(new_net_202),
		.d(new_net_429)
	);

	spl4L new_net_418_v_fanout (
		.a(new_net_418),
		.b(new_net_232),
		.c(new_net_230),
		.d(new_net_231),
		.e(new_net_229)
	);

	bfr new_net_998_bfr_before (
		.din(new_net_998),
		.dout(new_net_119)
	);

	bfr new_net_999_bfr_before (
		.din(new_net_999),
		.dout(new_net_998)
	);

	bfr new_net_1000_bfr_before (
		.din(new_net_1000),
		.dout(new_net_999)
	);

	bfr new_net_1001_bfr_before (
		.din(new_net_1001),
		.dout(new_net_1000)
	);

	bfr new_net_1002_bfr_before (
		.din(new_net_1002),
		.dout(new_net_1001)
	);

	bfr new_net_1003_bfr_before (
		.din(new_net_1003),
		.dout(new_net_1002)
	);

	bfr new_net_1004_bfr_before (
		.din(new_net_1004),
		.dout(new_net_1003)
	);

	bfr new_net_1005_bfr_before (
		.din(new_net_1005),
		.dout(new_net_1004)
	);

	spl2 new_net_433_v_fanout (
		.a(new_net_433),
		.b(new_net_1005),
		.c(new_net_121)
	);

	bfr new_net_1006_bfr_before (
		.din(new_net_1006),
		.dout(new_net_71)
	);

	bfr new_net_1007_bfr_before (
		.din(new_net_1007),
		.dout(new_net_1006)
	);

	bfr new_net_1008_bfr_before (
		.din(new_net_1008),
		.dout(new_net_1007)
	);

	bfr new_net_1009_bfr_before (
		.din(new_net_1009),
		.dout(new_net_1008)
	);

	bfr new_net_1010_bfr_before (
		.din(new_net_1010),
		.dout(new_net_1009)
	);

	bfr new_net_1011_bfr_before (
		.din(new_net_1011),
		.dout(new_net_1010)
	);

	spl4L new_net_407_v_fanout (
		.a(new_net_407),
		.b(new_net_75),
		.c(new_net_1011),
		.d(new_net_76),
		.e(new_net_73)
	);

	spl3L new_net_406_v_fanout (
		.a(new_net_406),
		.b(new_net_72),
		.c(new_net_70),
		.d(new_net_74)
	);

	spl4L new_net_419_v_fanout (
		.a(new_net_419),
		.b(new_net_235),
		.c(new_net_234),
		.d(new_net_236),
		.e(new_net_233)
	);

	bfr new_net_1012_bfr_before (
		.din(new_net_1012),
		.dout(new_net_389)
	);

	spl2 new_net_430_v_fanout (
		.a(new_net_430),
		.b(new_net_1012),
		.c(new_net_391)
	);

	spl2 _273__v_fanout (
		.a(_273_),
		.b(new_net_260),
		.c(new_net_259)
	);

	bfr new_net_1013_bfr_before (
		.din(new_net_1013),
		.dout(new_net_401)
	);

	bfr new_net_1014_bfr_before (
		.din(new_net_1014),
		.dout(new_net_1013)
	);

	spl3L N130_v_fanout (
		.a(N130),
		.b(new_net_271),
		.c(new_net_1014),
		.d(new_net_273)
	);

	bfr new_net_1015_bfr_before (
		.din(new_net_1015),
		.dout(new_net_170)
	);

	bfr new_net_1016_bfr_before (
		.din(new_net_1016),
		.dout(new_net_1015)
	);

	bfr new_net_1017_bfr_before (
		.din(new_net_1017),
		.dout(new_net_1016)
	);

	bfr new_net_1018_bfr_before (
		.din(new_net_1018),
		.dout(new_net_1017)
	);

	bfr new_net_1019_bfr_before (
		.din(new_net_1019),
		.dout(new_net_1018)
	);

	bfr new_net_1020_bfr_before (
		.din(new_net_1020),
		.dout(new_net_1019)
	);

	bfr new_net_1021_bfr_before (
		.din(new_net_1021),
		.dout(new_net_1020)
	);

	bfr new_net_1022_bfr_before (
		.din(new_net_1022),
		.dout(new_net_1021)
	);

	bfr new_net_1023_bfr_before (
		.din(new_net_1023),
		.dout(new_net_1022)
	);

	bfr new_net_1024_bfr_before (
		.din(new_net_1024),
		.dout(new_net_173)
	);

	spl4L N116_v_fanout (
		.a(N116),
		.b(new_net_1024),
		.c(new_net_171),
		.d(new_net_172),
		.e(new_net_1023)
	);

	spl3L N96_v_fanout (
		.a(N96),
		.b(new_net_120),
		.c(new_net_433),
		.d(new_net_122)
	);

	bfr new_net_1025_bfr_before (
		.din(new_net_1025),
		.dout(new_net_414)
	);

	bfr new_net_1026_bfr_before (
		.din(new_net_1026),
		.dout(new_net_1025)
	);

	bfr new_net_1027_bfr_before (
		.din(new_net_1027),
		.dout(new_net_1026)
	);

	bfr new_net_1028_bfr_before (
		.din(new_net_1028),
		.dout(new_net_1027)
	);

	bfr new_net_1029_bfr_before (
		.din(new_net_1029),
		.dout(new_net_1028)
	);

	bfr new_net_1030_bfr_before (
		.din(new_net_1030),
		.dout(new_net_1029)
	);

	spl3L N189_v_fanout (
		.a(N189),
		.b(new_net_1030),
		.c(new_net_152),
		.d(new_net_156)
	);

	bfr new_net_1031_bfr_before (
		.din(new_net_1031),
		.dout(new_net_168)
	);

	bfr new_net_1032_bfr_before (
		.din(new_net_1032),
		.dout(new_net_1031)
	);

	bfr new_net_1033_bfr_before (
		.din(new_net_1033),
		.dout(new_net_1032)
	);

	bfr new_net_1034_bfr_before (
		.din(new_net_1034),
		.dout(new_net_1033)
	);

	bfr new_net_1035_bfr_before (
		.din(new_net_1035),
		.dout(new_net_1034)
	);

	bfr new_net_1036_bfr_before (
		.din(new_net_1036),
		.dout(new_net_1035)
	);

	bfr new_net_1037_bfr_before (
		.din(new_net_1037),
		.dout(new_net_1036)
	);

	spl4L N195_v_fanout (
		.a(N195),
		.b(new_net_1037),
		.c(new_net_169),
		.d(new_net_167),
		.e(new_net_166)
	);

	bfr new_net_1038_bfr_before (
		.din(new_net_1038),
		.dout(new_net_412)
	);

	bfr new_net_1039_bfr_before (
		.din(new_net_1039),
		.dout(new_net_1038)
	);

	bfr new_net_1040_bfr_before (
		.din(new_net_1040),
		.dout(new_net_1039)
	);

	bfr new_net_1041_bfr_before (
		.din(new_net_1041),
		.dout(new_net_1040)
	);

	bfr new_net_1042_bfr_before (
		.din(new_net_1042),
		.dout(new_net_1041)
	);

	bfr new_net_1043_bfr_before (
		.din(new_net_1043),
		.dout(new_net_1042)
	);

	spl3L N183_v_fanout (
		.a(N183),
		.b(new_net_1043),
		.c(new_net_133),
		.d(new_net_135)
	);

	bfr new_net_1044_bfr_before (
		.din(new_net_1044),
		.dout(new_net_303)
	);

	bfr new_net_1045_bfr_before (
		.din(new_net_1045),
		.dout(new_net_1044)
	);

	bfr new_net_1046_bfr_before (
		.din(new_net_1046),
		.dout(new_net_1045)
	);

	bfr new_net_1047_bfr_before (
		.din(new_net_1047),
		.dout(new_net_1046)
	);

	bfr new_net_1048_bfr_before (
		.din(new_net_1048),
		.dout(new_net_1047)
	);

	bfr new_net_1049_bfr_before (
		.din(new_net_1049),
		.dout(new_net_1048)
	);

	bfr new_net_1050_bfr_before (
		.din(new_net_1050),
		.dout(new_net_1049)
	);

	bfr new_net_1051_bfr_before (
		.din(new_net_1051),
		.dout(new_net_1050)
	);

	bfr new_net_1052_bfr_before (
		.din(new_net_1052),
		.dout(new_net_1051)
	);

	bfr new_net_1053_bfr_before (
		.din(new_net_1053),
		.dout(new_net_1052)
	);

	bfr new_net_1054_bfr_before (
		.din(new_net_1054),
		.dout(new_net_1053)
	);

	bfr new_net_1055_bfr_before (
		.din(new_net_1055),
		.dout(new_net_1054)
	);

	bfr new_net_1056_bfr_before (
		.din(new_net_1056),
		.dout(new_net_1055)
	);

	bfr new_net_1057_bfr_before (
		.din(new_net_1057),
		.dout(new_net_1056)
	);

	bfr new_net_1058_bfr_before (
		.din(new_net_1058),
		.dout(new_net_1057)
	);

	spl2 N237_v_fanout (
		.a(N237),
		.b(new_net_1058),
		.c(new_net_302)
	);

	bfr new_net_1059_bfr_before (
		.din(new_net_1059),
		.dout(new_net_402)
	);

	bfr new_net_1060_bfr_before (
		.din(new_net_1060),
		.dout(new_net_1059)
	);

	bfr new_net_1061_bfr_before (
		.din(new_net_1061),
		.dout(new_net_1060)
	);

	bfr new_net_1062_bfr_before (
		.din(new_net_1062),
		.dout(new_net_1061)
	);

	bfr new_net_1063_bfr_before (
		.din(new_net_1063),
		.dout(new_net_1062)
	);

	bfr new_net_1064_bfr_before (
		.din(new_net_1064),
		.dout(new_net_1063)
	);

	spl3L N159_v_fanout (
		.a(N159),
		.b(new_net_40),
		.c(new_net_36),
		.d(new_net_1064)
	);

	bfr new_net_1065_bfr_after (
		.din(N146),
		.dout(new_net_1065)
	);

	bfr new_net_1066_bfr_after (
		.din(new_net_1065),
		.dout(new_net_1066)
	);

	bfr new_net_1067_bfr_after (
		.din(new_net_1066),
		.dout(new_net_1067)
	);

	bfr new_net_1068_bfr_after (
		.din(new_net_1067),
		.dout(new_net_1068)
	);

	bfr new_net_1069_bfr_after (
		.din(new_net_1068),
		.dout(new_net_1069)
	);

	bfr new_net_1070_bfr_after (
		.din(new_net_1069),
		.dout(new_net_1070)
	);

	bfr new_net_1071_bfr_after (
		.din(new_net_1070),
		.dout(new_net_1071)
	);

	bfr new_net_1072_bfr_after (
		.din(new_net_1071),
		.dout(new_net_1072)
	);

	bfr new_net_1073_bfr_before (
		.din(new_net_1073),
		.dout(new_net_345)
	);

	bfr new_net_1074_bfr_before (
		.din(new_net_1074),
		.dout(new_net_1073)
	);

	spl2 N146_v_fanout (
		.a(new_net_1072),
		.b(new_net_346),
		.c(new_net_1074)
	);

	spl2 N135_v_fanout (
		.a(N135),
		.b(new_net_288),
		.c(new_net_287)
	);

	bfr new_net_1075_bfr_after (
		.din(N207),
		.dout(new_net_1075)
	);

	bfr new_net_1076_bfr_after (
		.din(new_net_1075),
		.dout(new_net_1076)
	);

	bfr new_net_1077_bfr_after (
		.din(new_net_1076),
		.dout(new_net_1077)
	);

	spl2 N207_v_fanout (
		.a(new_net_1077),
		.b(new_net_217),
		.c(new_net_216)
	);

	bfr new_net_1078_bfr_before (
		.din(new_net_1078),
		.dout(new_net_416)
	);

	bfr new_net_1079_bfr_before (
		.din(new_net_1079),
		.dout(new_net_1078)
	);

	bfr new_net_1080_bfr_before (
		.din(new_net_1080),
		.dout(new_net_1079)
	);

	bfr new_net_1081_bfr_before (
		.din(new_net_1081),
		.dout(new_net_1080)
	);

	bfr new_net_1082_bfr_before (
		.din(new_net_1082),
		.dout(new_net_1081)
	);

	bfr new_net_1083_bfr_before (
		.din(new_net_1083),
		.dout(new_net_1082)
	);

	spl3L N201_v_fanout (
		.a(N201),
		.b(new_net_181),
		.c(new_net_183),
		.d(new_net_1083)
	);

	bfr new_net_1084_bfr_after (
		.din(N91),
		.dout(new_net_1084)
	);

	bfr new_net_1085_bfr_before (
		.din(new_net_1085),
		.dout(new_net_432)
	);

	spl2 N91_v_fanout (
		.a(new_net_1084),
		.b(new_net_1085),
		.c(new_net_106)
	);

	bfr new_net_1086_bfr_before (
		.din(new_net_1086),
		.dout(new_net_110)
	);

	bfr new_net_1087_bfr_before (
		.din(new_net_1087),
		.dout(new_net_1086)
	);

	bfr new_net_1088_bfr_before (
		.din(new_net_1088),
		.dout(new_net_1087)
	);

	bfr new_net_1089_bfr_before (
		.din(new_net_1089),
		.dout(new_net_1088)
	);

	bfr new_net_1090_bfr_before (
		.din(new_net_1090),
		.dout(new_net_1089)
	);

	bfr new_net_1091_bfr_before (
		.din(new_net_1091),
		.dout(new_net_1090)
	);

	bfr new_net_1092_bfr_before (
		.din(new_net_1092),
		.dout(new_net_1091)
	);

	bfr new_net_1093_bfr_before (
		.din(new_net_1093),
		.dout(new_net_1092)
	);

	spl3L N1_v_fanout (
		.a(N1),
		.b(new_net_1093),
		.c(new_net_108),
		.d(new_net_109)
	);

	spl3L N255_v_fanout (
		.a(N255),
		.b(new_net_337),
		.c(new_net_335),
		.d(new_net_336)
	);

	bfr new_net_1094_bfr_after (
		.din(N153),
		.dout(new_net_1094)
	);

	bfr new_net_1095_bfr_after (
		.din(new_net_1094),
		.dout(new_net_1095)
	);

	bfr new_net_1096_bfr_after (
		.din(new_net_1095),
		.dout(new_net_1096)
	);

	bfr new_net_1097_bfr_after (
		.din(new_net_1096),
		.dout(new_net_1097)
	);

	bfr new_net_1098_bfr_after (
		.din(new_net_1097),
		.dout(new_net_1098)
	);

	bfr new_net_1099_bfr_after (
		.din(new_net_1098),
		.dout(new_net_1099)
	);

	bfr new_net_1100_bfr_after (
		.din(new_net_1099),
		.dout(new_net_1100)
	);

	bfr new_net_1101_bfr_after (
		.din(new_net_1100),
		.dout(new_net_1101)
	);

	bfr new_net_1102_bfr_before (
		.din(new_net_1102),
		.dout(new_net_393)
	);

	bfr new_net_1103_bfr_before (
		.din(new_net_1103),
		.dout(new_net_1102)
	);

	spl2 N153_v_fanout (
		.a(new_net_1101),
		.b(new_net_1103),
		.c(new_net_392)
	);

	bfr new_net_1104_bfr_before (
		.din(new_net_1104),
		.dout(new_net_311)
	);

	spl4L N138_v_fanout (
		.a(N138),
		.b(new_net_310),
		.c(new_net_312),
		.d(new_net_1104),
		.e(new_net_309)
	);

	bfr new_net_1105_bfr_after (
		.din(N149),
		.dout(new_net_1105)
	);

	bfr new_net_1106_bfr_after (
		.din(new_net_1105),
		.dout(new_net_1106)
	);

	bfr new_net_1107_bfr_after (
		.din(new_net_1106),
		.dout(new_net_1107)
	);

	bfr new_net_1108_bfr_after (
		.din(new_net_1107),
		.dout(new_net_1108)
	);

	bfr new_net_1109_bfr_after (
		.din(new_net_1108),
		.dout(new_net_1109)
	);

	bfr new_net_1110_bfr_after (
		.din(new_net_1109),
		.dout(new_net_1110)
	);

	bfr new_net_1111_bfr_after (
		.din(new_net_1110),
		.dout(new_net_1111)
	);

	bfr new_net_1112_bfr_after (
		.din(new_net_1111),
		.dout(new_net_1112)
	);

	bfr new_net_1113_bfr_before (
		.din(new_net_1113),
		.dout(new_net_368)
	);

	bfr new_net_1114_bfr_before (
		.din(new_net_1114),
		.dout(new_net_1113)
	);

	spl2 N149_v_fanout (
		.a(new_net_1112),
		.b(new_net_369),
		.c(new_net_1114)
	);

	spl3L N42_v_fanout (
		.a(N42),
		.b(new_net_204),
		.c(new_net_203),
		.d(new_net_428)
	);

	bfr new_net_1115_bfr_before (
		.din(new_net_1115),
		.dout(new_net_127)
	);

	bfr new_net_1116_bfr_before (
		.din(new_net_1116),
		.dout(new_net_128)
	);

	bfr new_net_1117_bfr_before (
		.din(new_net_1117),
		.dout(new_net_1116)
	);

	bfr new_net_1118_bfr_before (
		.din(new_net_1118),
		.dout(new_net_1117)
	);

	bfr new_net_1119_bfr_before (
		.din(new_net_1119),
		.dout(new_net_1118)
	);

	bfr new_net_1120_bfr_before (
		.din(new_net_1120),
		.dout(new_net_1119)
	);

	bfr new_net_1121_bfr_before (
		.din(new_net_1121),
		.dout(new_net_1120)
	);

	bfr new_net_1122_bfr_before (
		.din(new_net_1122),
		.dout(new_net_1121)
	);

	bfr new_net_1123_bfr_before (
		.din(new_net_1123),
		.dout(new_net_1122)
	);

	bfr new_net_1124_bfr_before (
		.din(new_net_1124),
		.dout(new_net_1123)
	);

	spl4L N101_v_fanout (
		.a(N101),
		.b(new_net_130),
		.c(new_net_1124),
		.d(new_net_129),
		.e(new_net_1115)
	);

	spl2 N75_v_fanout (
		.a(N75),
		.b(new_net_139),
		.c(new_net_138)
	);

	bfr new_net_1125_bfr_after (
		.din(N228),
		.dout(new_net_1125)
	);

	bfr new_net_1126_bfr_after (
		.din(new_net_1125),
		.dout(new_net_1126)
	);

	bfr new_net_1127_bfr_after (
		.din(new_net_1126),
		.dout(new_net_1127)
	);

	bfr new_net_1128_bfr_after (
		.din(new_net_1127),
		.dout(new_net_1128)
	);

	bfr new_net_1129_bfr_after (
		.din(new_net_1128),
		.dout(new_net_1129)
	);

	bfr new_net_1130_bfr_after (
		.din(new_net_1129),
		.dout(new_net_1130)
	);

	bfr new_net_1131_bfr_after (
		.din(new_net_1130),
		.dout(new_net_1131)
	);

	bfr new_net_1132_bfr_after (
		.din(new_net_1131),
		.dout(new_net_1132)
	);

	bfr new_net_1133_bfr_after (
		.din(new_net_1132),
		.dout(new_net_1133)
	);

	bfr new_net_1134_bfr_after (
		.din(new_net_1133),
		.dout(new_net_1134)
	);

	bfr new_net_1135_bfr_after (
		.din(new_net_1134),
		.dout(new_net_1135)
	);

	bfr new_net_1136_bfr_after (
		.din(new_net_1135),
		.dout(new_net_1136)
	);

	bfr new_net_1137_bfr_after (
		.din(new_net_1136),
		.dout(new_net_1137)
	);

	bfr new_net_1138_bfr_after (
		.din(new_net_1137),
		.dout(new_net_1138)
	);

	bfr new_net_1139_bfr_after (
		.din(new_net_1138),
		.dout(new_net_1139)
	);

	bfr new_net_1140_bfr_after (
		.din(new_net_1139),
		.dout(new_net_1140)
	);

	spl4L N228_v_fanout (
		.a(new_net_1140),
		.b(new_net_284),
		.c(new_net_280),
		.d(new_net_424),
		.e(new_net_281)
	);

	bfr new_net_1141_bfr_before (
		.din(new_net_1141),
		.dout(new_net_431)
	);

	bfr new_net_1142_bfr_before (
		.din(new_net_1142),
		.dout(new_net_1141)
	);

	bfr new_net_1143_bfr_before (
		.din(new_net_1143),
		.dout(new_net_1142)
	);

	bfr new_net_1144_bfr_before (
		.din(new_net_1144),
		.dout(new_net_1143)
	);

	bfr new_net_1145_bfr_before (
		.din(new_net_1145),
		.dout(new_net_1144)
	);

	spl2 N55_v_fanout (
		.a(N55),
		.b(new_net_25),
		.c(new_net_1145)
	);

	bfr new_net_1146_bfr_after (
		.din(N268),
		.dout(new_net_1146)
	);

	bfr new_net_1147_bfr_before (
		.din(new_net_1147),
		.dout(new_net_30)
	);

	bfr new_net_1148_bfr_before (
		.din(new_net_1148),
		.dout(new_net_1147)
	);

	bfr new_net_1149_bfr_before (
		.din(new_net_1149),
		.dout(new_net_1148)
	);

	bfr new_net_1150_bfr_before (
		.din(new_net_1150),
		.dout(new_net_1149)
	);

	bfr new_net_1151_bfr_before (
		.din(new_net_1151),
		.dout(new_net_1150)
	);

	bfr new_net_1152_bfr_before (
		.din(new_net_1152),
		.dout(new_net_1151)
	);

	spl3L N268_v_fanout (
		.a(new_net_1146),
		.b(new_net_31),
		.c(new_net_29),
		.d(new_net_1152)
	);

	spl4L N59_v_fanout (
		.a(N59),
		.b(new_net_47),
		.c(new_net_45),
		.d(new_net_46),
		.e(new_net_44)
	);

	spl2 N8_v_fanout (
		.a(N8),
		.b(new_net_188),
		.c(new_net_187)
	);

	spl2 N210_v_fanout (
		.a(N210),
		.b(new_net_419),
		.c(new_net_418)
	);

	spl2 N51_v_fanout (
		.a(N51),
		.b(new_net_390),
		.c(new_net_430)
	);

	bfr new_net_1153_bfr_before (
		.din(new_net_1153),
		.dout(new_net_410)
	);

	bfr new_net_1154_bfr_before (
		.din(new_net_1154),
		.dout(new_net_1153)
	);

	bfr new_net_1155_bfr_before (
		.din(new_net_1155),
		.dout(new_net_1154)
	);

	bfr new_net_1156_bfr_before (
		.din(new_net_1156),
		.dout(new_net_1155)
	);

	bfr new_net_1157_bfr_before (
		.din(new_net_1157),
		.dout(new_net_1156)
	);

	bfr new_net_1158_bfr_before (
		.din(new_net_1158),
		.dout(new_net_1157)
	);

	spl3L N177_v_fanout (
		.a(N177),
		.b(new_net_114),
		.c(new_net_1158),
		.d(new_net_113)
	);

	spl2 N17_v_fanout (
		.a(N17),
		.b(new_net_407),
		.c(new_net_406)
	);

	bfr new_net_1159_bfr_before (
		.din(new_net_1159),
		.dout(new_net_192)
	);

	bfr new_net_1160_bfr_before (
		.din(new_net_1160),
		.dout(new_net_1159)
	);

	bfr new_net_1161_bfr_before (
		.din(new_net_1161),
		.dout(new_net_1160)
	);

	bfr new_net_1162_bfr_before (
		.din(new_net_1162),
		.dout(new_net_1161)
	);

	bfr new_net_1163_bfr_before (
		.din(new_net_1163),
		.dout(new_net_1162)
	);

	bfr new_net_1164_bfr_before (
		.din(new_net_1164),
		.dout(new_net_1163)
	);

	bfr new_net_1165_bfr_before (
		.din(new_net_1165),
		.dout(new_net_1164)
	);

	bfr new_net_1166_bfr_before (
		.din(new_net_1166),
		.dout(new_net_1165)
	);

	bfr new_net_1167_bfr_before (
		.din(new_net_1167),
		.dout(new_net_1166)
	);

	bfr new_net_1168_bfr_before (
		.din(new_net_1168),
		.dout(new_net_195)
	);

	spl4L N121_v_fanout (
		.a(N121),
		.b(new_net_1168),
		.c(new_net_193),
		.d(new_net_194),
		.e(new_net_1167)
	);

	bfr new_net_1169_bfr_after (
		.din(N126),
		.dout(new_net_1169)
	);

	bfr new_net_1170_bfr_after (
		.din(new_net_1169),
		.dout(new_net_1170)
	);

	bfr new_net_1171_bfr_after (
		.din(new_net_1170),
		.dout(new_net_1171)
	);

	bfr new_net_1172_bfr_before (
		.din(new_net_1172),
		.dout(new_net_226)
	);

	bfr new_net_1173_bfr_before (
		.din(new_net_1173),
		.dout(new_net_1172)
	);

	bfr new_net_1174_bfr_before (
		.din(new_net_1174),
		.dout(new_net_1173)
	);

	bfr new_net_1175_bfr_before (
		.din(new_net_1175),
		.dout(new_net_1174)
	);

	bfr new_net_1176_bfr_before (
		.din(new_net_1176),
		.dout(new_net_1175)
	);

	bfr new_net_1177_bfr_before (
		.din(new_net_1177),
		.dout(new_net_1176)
	);

	spl3L N126_v_fanout (
		.a(new_net_1171),
		.b(new_net_228),
		.c(new_net_1177),
		.d(new_net_227)
	);

	bfr new_net_1178_bfr_after (
		.din(N246),
		.dout(new_net_1178)
	);

	bfr new_net_1179_bfr_after (
		.din(new_net_1178),
		.dout(new_net_1179)
	);

	bfr new_net_1180_bfr_after (
		.din(new_net_1179),
		.dout(new_net_1180)
	);

	bfr new_net_1181_bfr_after (
		.din(new_net_1180),
		.dout(new_net_1181)
	);

	bfr new_net_1182_bfr_after (
		.din(new_net_1181),
		.dout(new_net_1182)
	);

	bfr new_net_1183_bfr_after (
		.din(new_net_1182),
		.dout(new_net_1183)
	);

	bfr new_net_1184_bfr_after (
		.din(new_net_1183),
		.dout(new_net_1184)
	);

	bfr new_net_1185_bfr_after (
		.din(new_net_1184),
		.dout(new_net_1185)
	);

	bfr new_net_1186_bfr_after (
		.din(new_net_1185),
		.dout(new_net_1186)
	);

	bfr new_net_1187_bfr_after (
		.din(new_net_1186),
		.dout(new_net_1187)
	);

	bfr new_net_1188_bfr_after (
		.din(new_net_1187),
		.dout(new_net_1188)
	);

	bfr new_net_1189_bfr_before (
		.din(new_net_1189),
		.dout(new_net_317)
	);

	spl2 N246_v_fanout (
		.a(new_net_1188),
		.b(new_net_426),
		.c(new_net_1189)
	);

	bfr new_net_1190_bfr_before (
		.din(new_net_1190),
		.dout(new_net_213)
	);

	bfr new_net_1191_bfr_before (
		.din(new_net_1191),
		.dout(new_net_1190)
	);

	spl2 N80_v_fanout (
		.a(N80),
		.b(new_net_1191),
		.c(new_net_212)
	);

	bfr new_net_1192_bfr_before (
		.din(new_net_1192),
		.dout(new_net_404)
	);

	bfr new_net_1193_bfr_before (
		.din(new_net_1193),
		.dout(new_net_1192)
	);

	bfr new_net_1194_bfr_before (
		.din(new_net_1194),
		.dout(new_net_1193)
	);

	bfr new_net_1195_bfr_before (
		.din(new_net_1195),
		.dout(new_net_1194)
	);

	bfr new_net_1196_bfr_before (
		.din(new_net_1196),
		.dout(new_net_1195)
	);

	bfr new_net_1197_bfr_before (
		.din(new_net_1197),
		.dout(new_net_1196)
	);

	spl3L N165_v_fanout (
		.a(N165),
		.b(new_net_57),
		.c(new_net_58),
		.d(new_net_1197)
	);

	bfr new_net_1198_bfr_before (
		.din(new_net_1198),
		.dout(new_net_157)
	);

	bfr new_net_1199_bfr_before (
		.din(new_net_1199),
		.dout(new_net_1198)
	);

	bfr new_net_1200_bfr_before (
		.din(new_net_1200),
		.dout(new_net_1199)
	);

	bfr new_net_1201_bfr_before (
		.din(new_net_1201),
		.dout(new_net_1200)
	);

	bfr new_net_1202_bfr_before (
		.din(new_net_1202),
		.dout(new_net_1201)
	);

	bfr new_net_1203_bfr_before (
		.din(new_net_1203),
		.dout(new_net_1202)
	);

	bfr new_net_1204_bfr_before (
		.din(new_net_1204),
		.dout(new_net_1203)
	);

	bfr new_net_1205_bfr_before (
		.din(new_net_1205),
		.dout(new_net_1204)
	);

	bfr new_net_1206_bfr_before (
		.din(new_net_1206),
		.dout(new_net_1205)
	);

	bfr new_net_1207_bfr_before (
		.din(new_net_1207),
		.dout(new_net_160)
	);

	spl4L N111_v_fanout (
		.a(N111),
		.b(new_net_1207),
		.c(new_net_159),
		.d(new_net_158),
		.e(new_net_1206)
	);

	spl2 N68_v_fanout (
		.a(N68),
		.b(new_net_62),
		.c(new_net_61)
	);

	bfr new_net_1208_bfr_before (
		.din(new_net_1208),
		.dout(new_net_143)
	);

	bfr new_net_1209_bfr_before (
		.din(new_net_1209),
		.dout(new_net_1208)
	);

	bfr new_net_1210_bfr_before (
		.din(new_net_1210),
		.dout(new_net_1209)
	);

	bfr new_net_1211_bfr_before (
		.din(new_net_1211),
		.dout(new_net_1210)
	);

	bfr new_net_1212_bfr_before (
		.din(new_net_1212),
		.dout(new_net_1211)
	);

	bfr new_net_1213_bfr_before (
		.din(new_net_1213),
		.dout(new_net_1212)
	);

	bfr new_net_1214_bfr_before (
		.din(new_net_1214),
		.dout(new_net_1213)
	);

	bfr new_net_1215_bfr_before (
		.din(new_net_1215),
		.dout(new_net_1214)
	);

	bfr new_net_1216_bfr_before (
		.din(new_net_1216),
		.dout(new_net_1215)
	);

	bfr new_net_1217_bfr_before (
		.din(new_net_1217),
		.dout(new_net_146)
	);

	spl4L N106_v_fanout (
		.a(N106),
		.b(new_net_1217),
		.c(new_net_144),
		.d(new_net_145),
		.e(new_net_1216)
	);

	spl2 N36_v_fanout (
		.a(N36),
		.b(new_net_66),
		.c(new_net_65)
	);

	bfr new_net_1218_bfr_before (
		.din(new_net_1218),
		.dout(new_net_247)
	);

	spl2 N13_v_fanout (
		.a(N13),
		.b(new_net_1218),
		.c(new_net_246)
	);

	bfr new_net_1219_bfr_after (
		.din(N143),
		.dout(new_net_1219)
	);

	bfr new_net_1220_bfr_after (
		.din(new_net_1219),
		.dout(new_net_1220)
	);

	bfr new_net_1221_bfr_after (
		.din(new_net_1220),
		.dout(new_net_1221)
	);

	bfr new_net_1222_bfr_after (
		.din(new_net_1221),
		.dout(new_net_1222)
	);

	bfr new_net_1223_bfr_after (
		.din(new_net_1222),
		.dout(new_net_1223)
	);

	bfr new_net_1224_bfr_after (
		.din(new_net_1223),
		.dout(new_net_1224)
	);

	bfr new_net_1225_bfr_after (
		.din(new_net_1224),
		.dout(new_net_1225)
	);

	bfr new_net_1226_bfr_after (
		.din(new_net_1225),
		.dout(new_net_1226)
	);

	bfr new_net_1227_bfr_before (
		.din(new_net_1227),
		.dout(new_net_328)
	);

	bfr new_net_1228_bfr_before (
		.din(new_net_1228),
		.dout(new_net_1227)
	);

	spl2 N143_v_fanout (
		.a(new_net_1226),
		.b(new_net_329),
		.c(new_net_1228)
	);

	spl3L N29_v_fanout (
		.a(N29),
		.b(new_net_50),
		.c(new_net_48),
		.d(new_net_49)
	);

	bfr new_net_1229_bfr_before (
		.din(new_net_1229),
		.dout(new_net_420)
	);

	bfr new_net_1230_bfr_before (
		.din(new_net_1230),
		.dout(new_net_1229)
	);

	bfr new_net_1231_bfr_before (
		.din(new_net_1231),
		.dout(new_net_1230)
	);

	bfr new_net_1232_bfr_before (
		.din(new_net_1232),
		.dout(new_net_1231)
	);

	bfr new_net_1233_bfr_before (
		.din(new_net_1233),
		.dout(new_net_1232)
	);

	bfr new_net_1234_bfr_before (
		.din(new_net_1234),
		.dout(new_net_1233)
	);

	bfr new_net_1235_bfr_before (
		.din(new_net_1235),
		.dout(new_net_1234)
	);

	bfr new_net_1236_bfr_before (
		.din(new_net_1236),
		.dout(new_net_1235)
	);

	bfr new_net_1237_bfr_before (
		.din(new_net_1237),
		.dout(new_net_1236)
	);

	bfr new_net_1238_bfr_before (
		.din(new_net_1238),
		.dout(new_net_1237)
	);

	bfr new_net_1239_bfr_before (
		.din(new_net_1239),
		.dout(new_net_1238)
	);

	bfr new_net_1240_bfr_before (
		.din(new_net_1240),
		.dout(new_net_1239)
	);

	bfr new_net_1241_bfr_before (
		.din(new_net_1241),
		.dout(new_net_1240)
	);

	bfr new_net_1242_bfr_before (
		.din(new_net_1242),
		.dout(new_net_1241)
	);

	bfr new_net_1243_bfr_before (
		.din(new_net_1243),
		.dout(new_net_1242)
	);

	spl2 N219_v_fanout (
		.a(N219),
		.b(new_net_1243),
		.c(new_net_268)
	);

	bfr new_net_1244_bfr_before (
		.din(new_net_1244),
		.dout(new_net_398)
	);

	bfr new_net_1245_bfr_before (
		.din(new_net_1245),
		.dout(new_net_1244)
	);

	bfr new_net_1246_bfr_before (
		.din(new_net_1246),
		.dout(new_net_1245)
	);

	bfr new_net_1247_bfr_before (
		.din(new_net_1247),
		.dout(new_net_1246)
	);

	bfr new_net_1248_bfr_before (
		.din(new_net_1248),
		.dout(new_net_1247)
	);

	bfr new_net_1249_bfr_before (
		.din(new_net_1249),
		.dout(new_net_1248)
	);

	bfr new_net_1250_bfr_before (
		.din(new_net_1250),
		.dout(new_net_1249)
	);

	bfr new_net_1251_bfr_before (
		.din(new_net_1251),
		.dout(new_net_1250)
	);

	bfr new_net_1252_bfr_before (
		.din(new_net_1252),
		.dout(new_net_1251)
	);

	bfr new_net_1253_bfr_before (
		.din(new_net_1253),
		.dout(new_net_1252)
	);

	bfr new_net_1254_bfr_before (
		.din(new_net_1254),
		.dout(new_net_1253)
	);

	bfr new_net_1255_bfr_before (
		.din(new_net_1255),
		.dout(new_net_1254)
	);

	bfr new_net_1256_bfr_before (
		.din(new_net_1256),
		.dout(new_net_1255)
	);

	bfr new_net_1257_bfr_before (
		.din(new_net_1257),
		.dout(new_net_1256)
	);

	bfr new_net_1258_bfr_before (
		.din(new_net_1258),
		.dout(new_net_1257)
	);

	bfr new_net_1259_bfr_before (
		.din(new_net_1259),
		.dout(new_net_1258)
	);

	bfr new_net_1260_bfr_before (
		.din(new_net_1260),
		.dout(new_net_1259)
	);

	spl2 N261_v_fanout (
		.a(N261),
		.b(new_net_1260),
		.c(new_net_397)
	);

	bfr new_net_1261_bfr_before (
		.din(new_net_1261),
		.dout(new_net_408)
	);

	bfr new_net_1262_bfr_before (
		.din(new_net_1262),
		.dout(new_net_1261)
	);

	bfr new_net_1263_bfr_before (
		.din(new_net_1263),
		.dout(new_net_1262)
	);

	bfr new_net_1264_bfr_before (
		.din(new_net_1264),
		.dout(new_net_1263)
	);

	bfr new_net_1265_bfr_before (
		.din(new_net_1265),
		.dout(new_net_1264)
	);

	bfr new_net_1266_bfr_before (
		.din(new_net_1266),
		.dout(new_net_1265)
	);

	spl3L N171_v_fanout (
		.a(N171),
		.b(new_net_95),
		.c(new_net_92),
		.d(new_net_1266)
	);

	bfr new_net_479_bfr_after (
		.din(_135_),
		.dout(new_net_479)
	);

	bfr new_net_500_bfr_after (
		.din(_183_),
		.dout(new_net_500)
	);

	bfr new_net_458_bfr_after (
		.din(_066_),
		.dout(new_net_458)
	);

	bfr new_net_1267_bfr_after (
		.din(_074_),
		.dout(new_net_1267)
	);

	bfr new_net_1268_bfr_after (
		.din(new_net_1267),
		.dout(new_net_1268)
	);

	bfr new_net_1269_bfr_after (
		.din(new_net_1268),
		.dout(new_net_1269)
	);

	bfr new_net_1270_bfr_after (
		.din(new_net_1269),
		.dout(new_net_1270)
	);

	bfr new_net_1271_bfr_after (
		.din(new_net_1270),
		.dout(new_net_1271)
	);

	bfr new_net_462_bfr_after (
		.din(new_net_1271),
		.dout(new_net_462)
	);

	bfr new_net_1272_bfr_after (
		.din(_146_),
		.dout(new_net_1272)
	);

	bfr new_net_1273_bfr_after (
		.din(new_net_1272),
		.dout(new_net_1273)
	);

	bfr new_net_1274_bfr_after (
		.din(new_net_1273),
		.dout(new_net_1274)
	);

	bfr new_net_1275_bfr_after (
		.din(new_net_1274),
		.dout(new_net_1275)
	);

	bfr new_net_1276_bfr_after (
		.din(new_net_1275),
		.dout(new_net_1276)
	);

	bfr new_net_483_bfr_after (
		.din(new_net_1276),
		.dout(new_net_483)
	);

	bfr new_net_1277_bfr_after (
		.din(_194_),
		.dout(new_net_1277)
	);

	bfr new_net_1278_bfr_after (
		.din(new_net_1277),
		.dout(new_net_1278)
	);

	bfr new_net_1279_bfr_after (
		.din(new_net_1278),
		.dout(new_net_1279)
	);

	bfr new_net_1280_bfr_after (
		.din(new_net_1279),
		.dout(new_net_1280)
	);

	bfr new_net_504_bfr_after (
		.din(new_net_1280),
		.dout(new_net_504)
	);

	bfr new_net_1281_bfr_after (
		.din(_001_),
		.dout(new_net_1281)
	);

	bfr new_net_451_bfr_after (
		.din(new_net_1281),
		.dout(new_net_451)
	);

	bfr new_net_1282_bfr_after (
		.din(new_net_550),
		.dout(new_net_1282)
	);

	bfr new_net_1283_bfr_after (
		.din(new_net_1282),
		.dout(new_net_1283)
	);

	bfr new_net_1284_bfr_after (
		.din(new_net_1283),
		.dout(new_net_1284)
	);

	bfr new_net_1285_bfr_after (
		.din(new_net_1284),
		.dout(new_net_1285)
	);

	bfr new_net_1286_bfr_after (
		.din(new_net_1285),
		.dout(new_net_1286)
	);

	bfr new_net_1287_bfr_after (
		.din(new_net_1286),
		.dout(new_net_1287)
	);

	bfr new_net_1288_bfr_after (
		.din(new_net_1287),
		.dout(new_net_1288)
	);

	bfr new_net_1289_bfr_after (
		.din(new_net_1288),
		.dout(new_net_1289)
	);

	bfr new_net_1290_bfr_after (
		.din(new_net_1289),
		.dout(new_net_1290)
	);

	bfr new_net_1291_bfr_after (
		.din(new_net_1290),
		.dout(new_net_1291)
	);

	bfr new_net_1292_bfr_after (
		.din(new_net_1291),
		.dout(new_net_1292)
	);

	bfr new_net_1293_bfr_after (
		.din(new_net_1292),
		.dout(new_net_1293)
	);

	bfr new_net_1294_bfr_after (
		.din(new_net_1293),
		.dout(new_net_1294)
	);

	bfr new_net_1295_bfr_after (
		.din(new_net_1294),
		.dout(new_net_1295)
	);

	bfr new_net_1296_bfr_after (
		.din(new_net_1295),
		.dout(new_net_1296)
	);

	bfr new_net_1297_bfr_after (
		.din(new_net_1296),
		.dout(new_net_1297)
	);

	bfr new_net_1298_bfr_after (
		.din(new_net_1297),
		.dout(new_net_1298)
	);

	bfr new_net_1299_bfr_after (
		.din(new_net_1298),
		.dout(new_net_1299)
	);

	bfr new_net_1300_bfr_after (
		.din(new_net_1299),
		.dout(new_net_1300)
	);

	bfr new_net_1301_bfr_after (
		.din(new_net_1300),
		.dout(new_net_1301)
	);

	bfr new_net_1302_bfr_after (
		.din(new_net_1301),
		.dout(new_net_1302)
	);

	bfr new_net_1303_bfr_after (
		.din(new_net_1302),
		.dout(new_net_1303)
	);

	bfr new_net_1304_bfr_after (
		.din(new_net_1303),
		.dout(new_net_1304)
	);

	bfr new_net_1305_bfr_after (
		.din(new_net_1304),
		.dout(new_net_1305)
	);

	bfr new_net_1306_bfr_after (
		.din(new_net_1305),
		.dout(new_net_1306)
	);

	bfr new_net_1307_bfr_after (
		.din(new_net_1306),
		.dout(new_net_1307)
	);

	bfr new_net_1308_bfr_after (
		.din(new_net_1307),
		.dout(new_net_1308)
	);

	bfr new_net_1309_bfr_after (
		.din(new_net_1308),
		.dout(new_net_1309)
	);

	bfr new_net_1310_bfr_after (
		.din(new_net_1309),
		.dout(new_net_1310)
	);

	bfr new_net_1311_bfr_after (
		.din(new_net_1310),
		.dout(new_net_1311)
	);

	bfr new_net_1312_bfr_after (
		.din(new_net_1311),
		.dout(new_net_1312)
	);

	bfr new_net_1313_bfr_after (
		.din(new_net_1312),
		.dout(new_net_1313)
	);

	bfr new_net_1314_bfr_after (
		.din(new_net_1313),
		.dout(new_net_1314)
	);

	bfr new_net_1315_bfr_after (
		.din(new_net_1314),
		.dout(new_net_1315)
	);

	bfr N448_bfr_after (
		.din(new_net_1315),
		.dout(N448)
	);

	bfr new_net_474_bfr_after (
		.din(_122_),
		.dout(new_net_474)
	);

	bfr new_net_1316_bfr_after (
		.din(_177_),
		.dout(new_net_1316)
	);

	bfr new_net_1317_bfr_after (
		.din(new_net_1316),
		.dout(new_net_1317)
	);

	bfr new_net_1318_bfr_after (
		.din(new_net_1317),
		.dout(new_net_1318)
	);

	bfr new_net_1319_bfr_after (
		.din(new_net_1318),
		.dout(new_net_1319)
	);

	bfr new_net_495_bfr_after (
		.din(new_net_1319),
		.dout(new_net_495)
	);

	bfr new_net_1320_bfr_after (
		.din(N74),
		.dout(new_net_1320)
	);

	bfr new_net_1321_bfr_after (
		.din(new_net_1320),
		.dout(new_net_1321)
	);

	bfr new_net_516_bfr_after (
		.din(new_net_1321),
		.dout(new_net_516)
	);

	bfr new_net_1322_bfr_after (
		.din(_151_),
		.dout(new_net_1322)
	);

	bfr new_net_1323_bfr_after (
		.din(new_net_1322),
		.dout(new_net_1323)
	);

	bfr new_net_1324_bfr_after (
		.din(new_net_1323),
		.dout(new_net_1324)
	);

	bfr new_net_1325_bfr_after (
		.din(new_net_1324),
		.dout(new_net_1325)
	);

	bfr new_net_1326_bfr_after (
		.din(new_net_1325),
		.dout(new_net_1326)
	);

	bfr new_net_1327_bfr_after (
		.din(new_net_1326),
		.dout(new_net_1327)
	);

	bfr new_net_1328_bfr_after (
		.din(new_net_1327),
		.dout(new_net_1328)
	);

	bfr new_net_1329_bfr_after (
		.din(new_net_1328),
		.dout(new_net_1329)
	);

	bfr new_net_1330_bfr_after (
		.din(new_net_1329),
		.dout(new_net_1330)
	);

	bfr new_net_1331_bfr_after (
		.din(new_net_1330),
		.dout(new_net_1331)
	);

	bfr new_net_1332_bfr_after (
		.din(new_net_1331),
		.dout(new_net_1332)
	);

	bfr new_net_1333_bfr_after (
		.din(new_net_1332),
		.dout(new_net_1333)
	);

	bfr new_net_1334_bfr_after (
		.din(new_net_1333),
		.dout(new_net_1334)
	);

	bfr new_net_1335_bfr_after (
		.din(new_net_1334),
		.dout(new_net_1335)
	);

	bfr new_net_487_bfr_after (
		.din(new_net_1335),
		.dout(new_net_487)
	);

	bfr new_net_508_bfr_after (
		.din(N260),
		.dout(new_net_508)
	);

	bfr new_net_466_bfr_after (
		.din(_078_),
		.dout(new_net_466)
	);

	bfr new_net_453_bfr_after (
		.din(_010_),
		.dout(new_net_453)
	);

	bfr new_net_470_bfr_after (
		.din(_110_),
		.dout(new_net_470)
	);

	bfr new_net_491_bfr_after (
		.din(_164_),
		.dout(new_net_491)
	);

	bfr new_net_512_bfr_after (
		.din(_211_),
		.dout(new_net_512)
	);

	bfr new_net_1336_bfr_after (
		.din(new_net_522),
		.dout(new_net_1336)
	);

	bfr new_net_1337_bfr_after (
		.din(new_net_1336),
		.dout(new_net_1337)
	);

	bfr new_net_1338_bfr_after (
		.din(new_net_1337),
		.dout(new_net_1338)
	);

	bfr new_net_1339_bfr_after (
		.din(new_net_1338),
		.dout(new_net_1339)
	);

	bfr new_net_1340_bfr_after (
		.din(new_net_1339),
		.dout(new_net_1340)
	);

	bfr new_net_1341_bfr_after (
		.din(new_net_1340),
		.dout(new_net_1341)
	);

	bfr new_net_1342_bfr_after (
		.din(new_net_1341),
		.dout(new_net_1342)
	);

	bfr new_net_1343_bfr_after (
		.din(new_net_1342),
		.dout(new_net_1343)
	);

	bfr new_net_1344_bfr_after (
		.din(new_net_1343),
		.dout(new_net_1344)
	);

	bfr new_net_1345_bfr_after (
		.din(new_net_1344),
		.dout(new_net_1345)
	);

	bfr new_net_1346_bfr_after (
		.din(new_net_1345),
		.dout(new_net_1346)
	);

	bfr new_net_1347_bfr_after (
		.din(new_net_1346),
		.dout(new_net_1347)
	);

	bfr new_net_1348_bfr_after (
		.din(new_net_1347),
		.dout(new_net_1348)
	);

	bfr new_net_1349_bfr_after (
		.din(new_net_1348),
		.dout(new_net_1349)
	);

	bfr new_net_1350_bfr_after (
		.din(new_net_1349),
		.dout(new_net_1350)
	);

	bfr new_net_1351_bfr_after (
		.din(new_net_1350),
		.dout(new_net_1351)
	);

	bfr new_net_1352_bfr_after (
		.din(new_net_1351),
		.dout(new_net_1352)
	);

	bfr N865_bfr_after (
		.din(new_net_1352),
		.dout(N865)
	);

	bfr new_net_1353_bfr_after (
		.din(N90),
		.dout(new_net_1353)
	);

	bfr new_net_518_bfr_after (
		.din(new_net_1353),
		.dout(new_net_518)
	);

	bfr new_net_1354_bfr_after (
		.din(new_net_530),
		.dout(new_net_1354)
	);

	bfr new_net_1355_bfr_after (
		.din(new_net_1354),
		.dout(new_net_1355)
	);

	bfr new_net_1356_bfr_after (
		.din(new_net_1355),
		.dout(new_net_1356)
	);

	bfr new_net_1357_bfr_after (
		.din(new_net_1356),
		.dout(new_net_1357)
	);

	bfr new_net_1358_bfr_after (
		.din(new_net_1357),
		.dout(new_net_1358)
	);

	bfr new_net_1359_bfr_after (
		.din(new_net_1358),
		.dout(new_net_1359)
	);

	bfr new_net_1360_bfr_after (
		.din(new_net_1359),
		.dout(new_net_1360)
	);

	bfr new_net_1361_bfr_after (
		.din(new_net_1360),
		.dout(new_net_1361)
	);

	bfr new_net_1362_bfr_after (
		.din(new_net_1361),
		.dout(new_net_1362)
	);

	bfr new_net_1363_bfr_after (
		.din(new_net_1362),
		.dout(new_net_1363)
	);

	bfr new_net_1364_bfr_after (
		.din(new_net_1363),
		.dout(new_net_1364)
	);

	bfr new_net_1365_bfr_after (
		.din(new_net_1364),
		.dout(new_net_1365)
	);

	bfr new_net_1366_bfr_after (
		.din(new_net_1365),
		.dout(new_net_1366)
	);

	bfr new_net_1367_bfr_after (
		.din(new_net_1366),
		.dout(new_net_1367)
	);

	bfr N864_bfr_after (
		.din(new_net_1367),
		.dout(N864)
	);

	bfr new_net_1368_bfr_after (
		.din(new_net_554),
		.dout(new_net_1368)
	);

	bfr new_net_1369_bfr_after (
		.din(new_net_1368),
		.dout(new_net_1369)
	);

	bfr new_net_1370_bfr_after (
		.din(new_net_1369),
		.dout(new_net_1370)
	);

	bfr new_net_1371_bfr_after (
		.din(new_net_1370),
		.dout(new_net_1371)
	);

	bfr new_net_1372_bfr_after (
		.din(new_net_1371),
		.dout(new_net_1372)
	);

	bfr new_net_1373_bfr_after (
		.din(new_net_1372),
		.dout(new_net_1373)
	);

	bfr new_net_1374_bfr_after (
		.din(new_net_1373),
		.dout(new_net_1374)
	);

	bfr new_net_1375_bfr_after (
		.din(new_net_1374),
		.dout(new_net_1375)
	);

	bfr new_net_1376_bfr_after (
		.din(new_net_1375),
		.dout(new_net_1376)
	);

	bfr new_net_1377_bfr_after (
		.din(new_net_1376),
		.dout(new_net_1377)
	);

	bfr new_net_1378_bfr_after (
		.din(new_net_1377),
		.dout(new_net_1378)
	);

	bfr new_net_1379_bfr_after (
		.din(new_net_1378),
		.dout(new_net_1379)
	);

	bfr new_net_1380_bfr_after (
		.din(new_net_1379),
		.dout(new_net_1380)
	);

	bfr new_net_1381_bfr_after (
		.din(new_net_1380),
		.dout(new_net_1381)
	);

	bfr new_net_1382_bfr_after (
		.din(new_net_1381),
		.dout(new_net_1382)
	);

	bfr new_net_1383_bfr_after (
		.din(new_net_1382),
		.dout(new_net_1383)
	);

	bfr new_net_1384_bfr_after (
		.din(new_net_1383),
		.dout(new_net_1384)
	);

	bfr new_net_1385_bfr_after (
		.din(new_net_1384),
		.dout(new_net_1385)
	);

	bfr new_net_1386_bfr_after (
		.din(new_net_1385),
		.dout(new_net_1386)
	);

	bfr new_net_1387_bfr_after (
		.din(new_net_1386),
		.dout(new_net_1387)
	);

	bfr new_net_1388_bfr_after (
		.din(new_net_1387),
		.dout(new_net_1388)
	);

	bfr new_net_1389_bfr_after (
		.din(new_net_1388),
		.dout(new_net_1389)
	);

	bfr new_net_1390_bfr_after (
		.din(new_net_1389),
		.dout(new_net_1390)
	);

	bfr new_net_1391_bfr_after (
		.din(new_net_1390),
		.dout(new_net_1391)
	);

	bfr new_net_1392_bfr_after (
		.din(new_net_1391),
		.dout(new_net_1392)
	);

	bfr new_net_1393_bfr_after (
		.din(new_net_1392),
		.dout(new_net_1393)
	);

	bfr new_net_1394_bfr_after (
		.din(new_net_1393),
		.dout(new_net_1394)
	);

	bfr new_net_1395_bfr_after (
		.din(new_net_1394),
		.dout(new_net_1395)
	);

	bfr new_net_1396_bfr_after (
		.din(new_net_1395),
		.dout(new_net_1396)
	);

	bfr new_net_1397_bfr_after (
		.din(new_net_1396),
		.dout(new_net_1397)
	);

	bfr new_net_1398_bfr_after (
		.din(new_net_1397),
		.dout(new_net_1398)
	);

	bfr new_net_1399_bfr_after (
		.din(new_net_1398),
		.dout(new_net_1399)
	);

	bfr new_net_1400_bfr_after (
		.din(new_net_1399),
		.dout(new_net_1400)
	);

	bfr new_net_1401_bfr_after (
		.din(new_net_1400),
		.dout(new_net_1401)
	);

	bfr new_net_1402_bfr_after (
		.din(new_net_1401),
		.dout(new_net_1402)
	);

	bfr new_net_1403_bfr_after (
		.din(new_net_1402),
		.dout(new_net_1403)
	);

	bfr N422_bfr_after (
		.din(new_net_1403),
		.dout(N422)
	);

	bfr new_net_1404_bfr_after (
		.din(new_net_528),
		.dout(new_net_1404)
	);

	bfr new_net_1405_bfr_after (
		.din(new_net_1404),
		.dout(new_net_1405)
	);

	bfr new_net_1406_bfr_after (
		.din(new_net_1405),
		.dout(new_net_1406)
	);

	bfr new_net_1407_bfr_after (
		.din(new_net_1406),
		.dout(new_net_1407)
	);

	bfr new_net_1408_bfr_after (
		.din(new_net_1407),
		.dout(new_net_1408)
	);

	bfr new_net_1409_bfr_after (
		.din(new_net_1408),
		.dout(new_net_1409)
	);

	bfr new_net_1410_bfr_after (
		.din(new_net_1409),
		.dout(new_net_1410)
	);

	bfr new_net_1411_bfr_after (
		.din(new_net_1410),
		.dout(new_net_1411)
	);

	bfr new_net_1412_bfr_after (
		.din(new_net_1411),
		.dout(new_net_1412)
	);

	bfr new_net_1413_bfr_after (
		.din(new_net_1412),
		.dout(new_net_1413)
	);

	bfr new_net_1414_bfr_after (
		.din(new_net_1413),
		.dout(new_net_1414)
	);

	bfr new_net_1415_bfr_after (
		.din(new_net_1414),
		.dout(new_net_1415)
	);

	bfr new_net_1416_bfr_after (
		.din(new_net_1415),
		.dout(new_net_1416)
	);

	bfr new_net_1417_bfr_after (
		.din(new_net_1416),
		.dout(new_net_1417)
	);

	bfr new_net_1418_bfr_after (
		.din(new_net_1417),
		.dout(new_net_1418)
	);

	bfr new_net_1419_bfr_after (
		.din(new_net_1418),
		.dout(new_net_1419)
	);

	bfr new_net_1420_bfr_after (
		.din(new_net_1419),
		.dout(new_net_1420)
	);

	bfr new_net_1421_bfr_after (
		.din(new_net_1420),
		.dout(new_net_1421)
	);

	bfr new_net_1422_bfr_after (
		.din(new_net_1421),
		.dout(new_net_1422)
	);

	bfr new_net_1423_bfr_after (
		.din(new_net_1422),
		.dout(new_net_1423)
	);

	bfr new_net_1424_bfr_after (
		.din(new_net_1423),
		.dout(new_net_1424)
	);

	bfr new_net_1425_bfr_after (
		.din(new_net_1424),
		.dout(new_net_1425)
	);

	bfr new_net_1426_bfr_after (
		.din(new_net_1425),
		.dout(new_net_1426)
	);

	bfr new_net_1427_bfr_after (
		.din(new_net_1426),
		.dout(new_net_1427)
	);

	bfr new_net_1428_bfr_after (
		.din(new_net_1427),
		.dout(new_net_1428)
	);

	bfr new_net_1429_bfr_after (
		.din(new_net_1428),
		.dout(new_net_1429)
	);

	bfr new_net_1430_bfr_after (
		.din(new_net_1429),
		.dout(new_net_1430)
	);

	bfr new_net_1431_bfr_after (
		.din(new_net_1430),
		.dout(new_net_1431)
	);

	bfr new_net_1432_bfr_after (
		.din(new_net_1431),
		.dout(new_net_1432)
	);

	bfr new_net_1433_bfr_after (
		.din(new_net_1432),
		.dout(new_net_1433)
	);

	bfr new_net_1434_bfr_after (
		.din(new_net_1433),
		.dout(new_net_1434)
	);

	bfr new_net_1435_bfr_after (
		.din(new_net_1434),
		.dout(new_net_1435)
	);

	bfr new_net_1436_bfr_after (
		.din(new_net_1435),
		.dout(new_net_1436)
	);

	bfr N419_bfr_after (
		.din(new_net_1436),
		.dout(N419)
	);

	bfr new_net_1437_bfr_after (
		.din(new_net_540),
		.dout(new_net_1437)
	);

	bfr new_net_1438_bfr_after (
		.din(new_net_1437),
		.dout(new_net_1438)
	);

	bfr new_net_1439_bfr_after (
		.din(new_net_1438),
		.dout(new_net_1439)
	);

	bfr new_net_1440_bfr_after (
		.din(new_net_1439),
		.dout(new_net_1440)
	);

	bfr new_net_1441_bfr_after (
		.din(new_net_1440),
		.dout(new_net_1441)
	);

	bfr new_net_1442_bfr_after (
		.din(new_net_1441),
		.dout(new_net_1442)
	);

	bfr new_net_1443_bfr_after (
		.din(new_net_1442),
		.dout(new_net_1443)
	);

	bfr new_net_1444_bfr_after (
		.din(new_net_1443),
		.dout(new_net_1444)
	);

	bfr new_net_1445_bfr_after (
		.din(new_net_1444),
		.dout(new_net_1445)
	);

	bfr new_net_1446_bfr_after (
		.din(new_net_1445),
		.dout(new_net_1446)
	);

	bfr new_net_1447_bfr_after (
		.din(new_net_1446),
		.dout(new_net_1447)
	);

	bfr new_net_1448_bfr_after (
		.din(new_net_1447),
		.dout(new_net_1448)
	);

	bfr new_net_1449_bfr_after (
		.din(new_net_1448),
		.dout(new_net_1449)
	);

	bfr new_net_1450_bfr_after (
		.din(new_net_1449),
		.dout(new_net_1450)
	);

	bfr new_net_1451_bfr_after (
		.din(new_net_1450),
		.dout(new_net_1451)
	);

	bfr new_net_1452_bfr_after (
		.din(new_net_1451),
		.dout(new_net_1452)
	);

	bfr new_net_1453_bfr_after (
		.din(new_net_1452),
		.dout(new_net_1453)
	);

	bfr new_net_1454_bfr_after (
		.din(new_net_1453),
		.dout(new_net_1454)
	);

	bfr new_net_1455_bfr_after (
		.din(new_net_1454),
		.dout(new_net_1455)
	);

	bfr new_net_1456_bfr_after (
		.din(new_net_1455),
		.dout(new_net_1456)
	);

	bfr new_net_1457_bfr_after (
		.din(new_net_1456),
		.dout(new_net_1457)
	);

	bfr new_net_1458_bfr_after (
		.din(new_net_1457),
		.dout(new_net_1458)
	);

	bfr new_net_1459_bfr_after (
		.din(new_net_1458),
		.dout(new_net_1459)
	);

	bfr new_net_1460_bfr_after (
		.din(new_net_1459),
		.dout(new_net_1460)
	);

	bfr new_net_1461_bfr_after (
		.din(new_net_1460),
		.dout(new_net_1461)
	);

	bfr new_net_1462_bfr_after (
		.din(new_net_1461),
		.dout(new_net_1462)
	);

	bfr new_net_1463_bfr_after (
		.din(new_net_1462),
		.dout(new_net_1463)
	);

	bfr new_net_1464_bfr_after (
		.din(new_net_1463),
		.dout(new_net_1464)
	);

	bfr new_net_1465_bfr_after (
		.din(new_net_1464),
		.dout(new_net_1465)
	);

	bfr new_net_1466_bfr_after (
		.din(new_net_1465),
		.dout(new_net_1466)
	);

	bfr new_net_1467_bfr_after (
		.din(new_net_1466),
		.dout(new_net_1467)
	);

	bfr new_net_1468_bfr_after (
		.din(new_net_1467),
		.dout(new_net_1468)
	);

	bfr new_net_1469_bfr_after (
		.din(new_net_1468),
		.dout(new_net_1469)
	);

	bfr new_net_1470_bfr_after (
		.din(new_net_1469),
		.dout(new_net_1470)
	);

	bfr new_net_1471_bfr_after (
		.din(new_net_1470),
		.dout(new_net_1471)
	);

	bfr N418_bfr_after (
		.din(new_net_1471),
		.dout(N418)
	);

	bfr new_net_1472_bfr_after (
		.din(new_net_552),
		.dout(new_net_1472)
	);

	bfr new_net_1473_bfr_after (
		.din(new_net_1472),
		.dout(new_net_1473)
	);

	bfr new_net_1474_bfr_after (
		.din(new_net_1473),
		.dout(new_net_1474)
	);

	bfr new_net_1475_bfr_after (
		.din(new_net_1474),
		.dout(new_net_1475)
	);

	bfr new_net_1476_bfr_after (
		.din(new_net_1475),
		.dout(new_net_1476)
	);

	bfr new_net_1477_bfr_after (
		.din(new_net_1476),
		.dout(new_net_1477)
	);

	bfr new_net_1478_bfr_after (
		.din(new_net_1477),
		.dout(new_net_1478)
	);

	bfr new_net_1479_bfr_after (
		.din(new_net_1478),
		.dout(new_net_1479)
	);

	bfr new_net_1480_bfr_after (
		.din(new_net_1479),
		.dout(new_net_1480)
	);

	bfr new_net_1481_bfr_after (
		.din(new_net_1480),
		.dout(new_net_1481)
	);

	bfr new_net_1482_bfr_after (
		.din(new_net_1481),
		.dout(new_net_1482)
	);

	bfr new_net_1483_bfr_after (
		.din(new_net_1482),
		.dout(new_net_1483)
	);

	bfr new_net_1484_bfr_after (
		.din(new_net_1483),
		.dout(new_net_1484)
	);

	bfr new_net_1485_bfr_after (
		.din(new_net_1484),
		.dout(new_net_1485)
	);

	bfr new_net_1486_bfr_after (
		.din(new_net_1485),
		.dout(new_net_1486)
	);

	bfr new_net_1487_bfr_after (
		.din(new_net_1486),
		.dout(new_net_1487)
	);

	bfr new_net_1488_bfr_after (
		.din(new_net_1487),
		.dout(new_net_1488)
	);

	bfr new_net_1489_bfr_after (
		.din(new_net_1488),
		.dout(new_net_1489)
	);

	bfr new_net_1490_bfr_after (
		.din(new_net_1489),
		.dout(new_net_1490)
	);

	bfr new_net_1491_bfr_after (
		.din(new_net_1490),
		.dout(new_net_1491)
	);

	bfr new_net_1492_bfr_after (
		.din(new_net_1491),
		.dout(new_net_1492)
	);

	bfr new_net_1493_bfr_after (
		.din(new_net_1492),
		.dout(new_net_1493)
	);

	bfr new_net_1494_bfr_after (
		.din(new_net_1493),
		.dout(new_net_1494)
	);

	bfr new_net_1495_bfr_after (
		.din(new_net_1494),
		.dout(new_net_1495)
	);

	bfr new_net_1496_bfr_after (
		.din(new_net_1495),
		.dout(new_net_1496)
	);

	bfr new_net_1497_bfr_after (
		.din(new_net_1496),
		.dout(new_net_1497)
	);

	bfr new_net_1498_bfr_after (
		.din(new_net_1497),
		.dout(new_net_1498)
	);

	bfr new_net_1499_bfr_after (
		.din(new_net_1498),
		.dout(new_net_1499)
	);

	bfr new_net_1500_bfr_after (
		.din(new_net_1499),
		.dout(new_net_1500)
	);

	bfr new_net_1501_bfr_after (
		.din(new_net_1500),
		.dout(new_net_1501)
	);

	bfr new_net_1502_bfr_after (
		.din(new_net_1501),
		.dout(new_net_1502)
	);

	bfr new_net_1503_bfr_after (
		.din(new_net_1502),
		.dout(new_net_1503)
	);

	bfr new_net_1504_bfr_after (
		.din(new_net_1503),
		.dout(new_net_1504)
	);

	bfr new_net_1505_bfr_after (
		.din(new_net_1504),
		.dout(new_net_1505)
	);

	bfr new_net_1506_bfr_after (
		.din(new_net_1505),
		.dout(new_net_1506)
	);

	bfr new_net_1507_bfr_after (
		.din(new_net_1506),
		.dout(new_net_1507)
	);

	bfr N389_bfr_after (
		.din(new_net_1507),
		.dout(N389)
	);

	bfr new_net_1508_bfr_after (
		.din(new_net_564),
		.dout(new_net_1508)
	);

	bfr new_net_1509_bfr_after (
		.din(new_net_1508),
		.dout(new_net_1509)
	);

	bfr new_net_1510_bfr_after (
		.din(new_net_1509),
		.dout(new_net_1510)
	);

	bfr new_net_1511_bfr_after (
		.din(new_net_1510),
		.dout(new_net_1511)
	);

	bfr new_net_1512_bfr_after (
		.din(new_net_1511),
		.dout(new_net_1512)
	);

	bfr new_net_1513_bfr_after (
		.din(new_net_1512),
		.dout(new_net_1513)
	);

	bfr new_net_1514_bfr_after (
		.din(new_net_1513),
		.dout(new_net_1514)
	);

	bfr new_net_1515_bfr_after (
		.din(new_net_1514),
		.dout(new_net_1515)
	);

	bfr new_net_1516_bfr_after (
		.din(new_net_1515),
		.dout(new_net_1516)
	);

	bfr new_net_1517_bfr_after (
		.din(new_net_1516),
		.dout(new_net_1517)
	);

	bfr new_net_1518_bfr_after (
		.din(new_net_1517),
		.dout(new_net_1518)
	);

	bfr N863_bfr_after (
		.din(new_net_1518),
		.dout(N863)
	);

	bfr new_net_461_bfr_after (
		.din(_071_),
		.dout(new_net_461)
	);

	bfr new_net_1519_bfr_after (
		.din(_061_),
		.dout(new_net_1519)
	);

	bfr new_net_1520_bfr_after (
		.din(new_net_1519),
		.dout(new_net_1520)
	);

	bfr new_net_1521_bfr_after (
		.din(new_net_1520),
		.dout(new_net_1521)
	);

	bfr new_net_1522_bfr_after (
		.din(new_net_1521),
		.dout(new_net_1522)
	);

	bfr new_net_1523_bfr_after (
		.din(new_net_1522),
		.dout(new_net_1523)
	);

	bfr new_net_1524_bfr_after (
		.din(new_net_1523),
		.dout(new_net_1524)
	);

	bfr new_net_1525_bfr_after (
		.din(new_net_1524),
		.dout(new_net_1525)
	);

	bfr new_net_1526_bfr_after (
		.din(new_net_1525),
		.dout(new_net_1526)
	);

	bfr new_net_1527_bfr_after (
		.din(new_net_1526),
		.dout(new_net_1527)
	);

	bfr new_net_457_bfr_after (
		.din(new_net_1527),
		.dout(new_net_457)
	);

	bfr new_net_482_bfr_after (
		.din(_139_),
		.dout(new_net_482)
	);

	bfr new_net_1528_bfr_after (
		.din(_193_),
		.dout(new_net_1528)
	);

	bfr new_net_1529_bfr_after (
		.din(new_net_1528),
		.dout(new_net_1529)
	);

	bfr new_net_1530_bfr_after (
		.din(new_net_1529),
		.dout(new_net_1530)
	);

	bfr new_net_1531_bfr_after (
		.din(new_net_1530),
		.dout(new_net_1531)
	);

	bfr new_net_503_bfr_after (
		.din(new_net_1531),
		.dout(new_net_503)
	);

	bfr new_net_1532_bfr_after (
		.din(_134_),
		.dout(new_net_1532)
	);

	bfr new_net_1533_bfr_after (
		.din(new_net_1532),
		.dout(new_net_1533)
	);

	bfr new_net_1534_bfr_after (
		.din(new_net_1533),
		.dout(new_net_1534)
	);

	bfr new_net_478_bfr_after (
		.din(new_net_1534),
		.dout(new_net_478)
	);

	bfr new_net_1535_bfr_after (
		.din(_181_),
		.dout(new_net_1535)
	);

	bfr new_net_1536_bfr_after (
		.din(new_net_1535),
		.dout(new_net_1536)
	);

	bfr new_net_1537_bfr_after (
		.din(new_net_1536),
		.dout(new_net_1537)
	);

	bfr new_net_1538_bfr_after (
		.din(new_net_1537),
		.dout(new_net_1538)
	);

	bfr new_net_499_bfr_after (
		.din(new_net_1538),
		.dout(new_net_499)
	);

	bfr new_net_486_bfr_after (
		.din(_150_),
		.dout(new_net_486)
	);

	bfr new_net_507_bfr_after (
		.din(_197_),
		.dout(new_net_507)
	);

	bfr new_net_494_bfr_after (
		.din(_176_),
		.dout(new_net_494)
	);

	bfr new_net_490_bfr_after (
		.din(_163_),
		.dout(new_net_490)
	);

	bfr new_net_1539_bfr_after (
		.din(_210_),
		.dout(new_net_1539)
	);

	bfr new_net_1540_bfr_after (
		.din(new_net_1539),
		.dout(new_net_1540)
	);

	bfr new_net_1541_bfr_after (
		.din(new_net_1540),
		.dout(new_net_1541)
	);

	bfr new_net_1542_bfr_after (
		.din(new_net_1541),
		.dout(new_net_1542)
	);

	bfr new_net_511_bfr_after (
		.din(new_net_1542),
		.dout(new_net_511)
	);

	bfr new_net_1543_bfr_after (
		.din(_215_),
		.dout(new_net_1543)
	);

	bfr new_net_1544_bfr_after (
		.din(new_net_1543),
		.dout(new_net_1544)
	);

	bfr new_net_515_bfr_after (
		.din(new_net_1544),
		.dout(new_net_515)
	);

	bfr new_net_1545_bfr_after (
		.din(_077_),
		.dout(new_net_1545)
	);

	bfr new_net_1546_bfr_after (
		.din(new_net_1545),
		.dout(new_net_1546)
	);

	bfr new_net_1547_bfr_after (
		.din(new_net_1546),
		.dout(new_net_1547)
	);

	bfr new_net_1548_bfr_after (
		.din(new_net_1547),
		.dout(new_net_1548)
	);

	bfr new_net_1549_bfr_after (
		.din(new_net_1548),
		.dout(new_net_1549)
	);

	bfr new_net_1550_bfr_after (
		.din(new_net_1549),
		.dout(new_net_1550)
	);

	bfr new_net_1551_bfr_after (
		.din(new_net_1550),
		.dout(new_net_1551)
	);

	bfr new_net_1552_bfr_after (
		.din(new_net_1551),
		.dout(new_net_1552)
	);

	bfr new_net_1553_bfr_after (
		.din(new_net_1552),
		.dout(new_net_1553)
	);

	bfr new_net_1554_bfr_after (
		.din(new_net_1553),
		.dout(new_net_1554)
	);

	bfr new_net_1555_bfr_after (
		.din(new_net_1554),
		.dout(new_net_1555)
	);

	bfr new_net_465_bfr_after (
		.din(new_net_1555),
		.dout(new_net_465)
	);

	bfr new_net_452_bfr_after (
		.din(N152),
		.dout(new_net_452)
	);

	bfr new_net_1556_bfr_after (
		.din(_098_),
		.dout(new_net_1556)
	);

	bfr new_net_1557_bfr_after (
		.din(new_net_1556),
		.dout(new_net_1557)
	);

	bfr new_net_1558_bfr_after (
		.din(new_net_1557),
		.dout(new_net_1558)
	);

	bfr new_net_1559_bfr_after (
		.din(new_net_1558),
		.dout(new_net_1559)
	);

	bfr new_net_1560_bfr_after (
		.din(new_net_1559),
		.dout(new_net_1560)
	);

	bfr new_net_469_bfr_after (
		.din(new_net_1560),
		.dout(new_net_469)
	);

	bfr new_net_473_bfr_after (
		.din(_121_),
		.dout(new_net_473)
	);

	bfr new_net_1561_bfr_after (
		.din(new_net_534),
		.dout(new_net_1561)
	);

	bfr new_net_1562_bfr_after (
		.din(new_net_1561),
		.dout(new_net_1562)
	);

	bfr new_net_1563_bfr_after (
		.din(new_net_1562),
		.dout(new_net_1563)
	);

	bfr new_net_1564_bfr_after (
		.din(new_net_1563),
		.dout(new_net_1564)
	);

	bfr new_net_1565_bfr_after (
		.din(new_net_1564),
		.dout(new_net_1565)
	);

	bfr new_net_1566_bfr_after (
		.din(new_net_1565),
		.dout(new_net_1566)
	);

	bfr new_net_1567_bfr_after (
		.din(new_net_1566),
		.dout(new_net_1567)
	);

	bfr new_net_1568_bfr_after (
		.din(new_net_1567),
		.dout(new_net_1568)
	);

	bfr new_net_1569_bfr_after (
		.din(new_net_1568),
		.dout(new_net_1569)
	);

	bfr new_net_1570_bfr_after (
		.din(new_net_1569),
		.dout(new_net_1570)
	);

	bfr new_net_1571_bfr_after (
		.din(new_net_1570),
		.dout(new_net_1571)
	);

	bfr new_net_1572_bfr_after (
		.din(new_net_1571),
		.dout(new_net_1572)
	);

	bfr new_net_1573_bfr_after (
		.din(new_net_1572),
		.dout(new_net_1573)
	);

	bfr new_net_1574_bfr_after (
		.din(new_net_1573),
		.dout(new_net_1574)
	);

	bfr new_net_1575_bfr_after (
		.din(new_net_1574),
		.dout(new_net_1575)
	);

	bfr new_net_1576_bfr_after (
		.din(new_net_1575),
		.dout(new_net_1576)
	);

	bfr new_net_1577_bfr_after (
		.din(new_net_1576),
		.dout(new_net_1577)
	);

	bfr new_net_1578_bfr_after (
		.din(new_net_1577),
		.dout(new_net_1578)
	);

	bfr new_net_1579_bfr_after (
		.din(new_net_1578),
		.dout(new_net_1579)
	);

	bfr new_net_1580_bfr_after (
		.din(new_net_1579),
		.dout(new_net_1580)
	);

	bfr new_net_1581_bfr_after (
		.din(new_net_1580),
		.dout(new_net_1581)
	);

	bfr new_net_1582_bfr_after (
		.din(new_net_1581),
		.dout(new_net_1582)
	);

	bfr new_net_1583_bfr_after (
		.din(new_net_1582),
		.dout(new_net_1583)
	);

	bfr new_net_1584_bfr_after (
		.din(new_net_1583),
		.dout(new_net_1584)
	);

	bfr new_net_1585_bfr_after (
		.din(new_net_1584),
		.dout(new_net_1585)
	);

	bfr new_net_1586_bfr_after (
		.din(new_net_1585),
		.dout(new_net_1586)
	);

	bfr new_net_1587_bfr_after (
		.din(new_net_1586),
		.dout(new_net_1587)
	);

	bfr new_net_1588_bfr_after (
		.din(new_net_1587),
		.dout(new_net_1588)
	);

	bfr new_net_1589_bfr_after (
		.din(new_net_1588),
		.dout(new_net_1589)
	);

	bfr new_net_1590_bfr_after (
		.din(new_net_1589),
		.dout(new_net_1590)
	);

	bfr new_net_1591_bfr_after (
		.din(new_net_1590),
		.dout(new_net_1591)
	);

	bfr new_net_1592_bfr_after (
		.din(new_net_1591),
		.dout(new_net_1592)
	);

	bfr new_net_1593_bfr_after (
		.din(new_net_1592),
		.dout(new_net_1593)
	);

	bfr new_net_1594_bfr_after (
		.din(new_net_1593),
		.dout(new_net_1594)
	);

	bfr N449_bfr_after (
		.din(new_net_1594),
		.dout(N449)
	);

	bfr new_net_1595_bfr_after (
		.din(new_net_558),
		.dout(new_net_1595)
	);

	bfr new_net_1596_bfr_after (
		.din(new_net_1595),
		.dout(new_net_1596)
	);

	bfr new_net_1597_bfr_after (
		.din(new_net_1596),
		.dout(new_net_1597)
	);

	bfr new_net_1598_bfr_after (
		.din(new_net_1597),
		.dout(new_net_1598)
	);

	bfr new_net_1599_bfr_after (
		.din(new_net_1598),
		.dout(new_net_1599)
	);

	bfr new_net_1600_bfr_after (
		.din(new_net_1599),
		.dout(new_net_1600)
	);

	bfr new_net_1601_bfr_after (
		.din(new_net_1600),
		.dout(new_net_1601)
	);

	bfr new_net_1602_bfr_after (
		.din(new_net_1601),
		.dout(new_net_1602)
	);

	bfr new_net_1603_bfr_after (
		.din(new_net_1602),
		.dout(new_net_1603)
	);

	bfr new_net_1604_bfr_after (
		.din(new_net_1603),
		.dout(new_net_1604)
	);

	bfr new_net_1605_bfr_after (
		.din(new_net_1604),
		.dout(new_net_1605)
	);

	bfr new_net_1606_bfr_after (
		.din(new_net_1605),
		.dout(new_net_1606)
	);

	bfr new_net_1607_bfr_after (
		.din(new_net_1606),
		.dout(new_net_1607)
	);

	bfr new_net_1608_bfr_after (
		.din(new_net_1607),
		.dout(new_net_1608)
	);

	bfr new_net_1609_bfr_after (
		.din(new_net_1608),
		.dout(new_net_1609)
	);

	bfr new_net_1610_bfr_after (
		.din(new_net_1609),
		.dout(new_net_1610)
	);

	bfr new_net_1611_bfr_after (
		.din(new_net_1610),
		.dout(new_net_1611)
	);

	bfr new_net_1612_bfr_after (
		.din(new_net_1611),
		.dout(new_net_1612)
	);

	bfr new_net_1613_bfr_after (
		.din(new_net_1612),
		.dout(new_net_1613)
	);

	bfr new_net_1614_bfr_after (
		.din(new_net_1613),
		.dout(new_net_1614)
	);

	bfr new_net_1615_bfr_after (
		.din(new_net_1614),
		.dout(new_net_1615)
	);

	bfr new_net_1616_bfr_after (
		.din(new_net_1615),
		.dout(new_net_1616)
	);

	bfr new_net_1617_bfr_after (
		.din(new_net_1616),
		.dout(new_net_1617)
	);

	bfr new_net_1618_bfr_after (
		.din(new_net_1617),
		.dout(new_net_1618)
	);

	bfr new_net_1619_bfr_after (
		.din(new_net_1618),
		.dout(new_net_1619)
	);

	bfr new_net_1620_bfr_after (
		.din(new_net_1619),
		.dout(new_net_1620)
	);

	bfr new_net_1621_bfr_after (
		.din(new_net_1620),
		.dout(new_net_1621)
	);

	bfr new_net_1622_bfr_after (
		.din(new_net_1621),
		.dout(new_net_1622)
	);

	bfr new_net_1623_bfr_after (
		.din(new_net_1622),
		.dout(new_net_1623)
	);

	bfr new_net_1624_bfr_after (
		.din(new_net_1623),
		.dout(new_net_1624)
	);

	bfr new_net_1625_bfr_after (
		.din(new_net_1624),
		.dout(new_net_1625)
	);

	bfr new_net_1626_bfr_after (
		.din(new_net_1625),
		.dout(new_net_1626)
	);

	bfr new_net_1627_bfr_after (
		.din(new_net_1626),
		.dout(new_net_1627)
	);

	bfr new_net_1628_bfr_after (
		.din(new_net_1627),
		.dout(new_net_1628)
	);

	bfr new_net_1629_bfr_after (
		.din(new_net_1628),
		.dout(new_net_1629)
	);

	bfr new_net_1630_bfr_after (
		.din(new_net_1629),
		.dout(new_net_1630)
	);

	bfr new_net_1631_bfr_after (
		.din(new_net_1630),
		.dout(new_net_1631)
	);

	bfr N423_bfr_after (
		.din(new_net_1631),
		.dout(N423)
	);

	bfr new_net_1632_bfr_after (
		.din(new_net_524),
		.dout(new_net_1632)
	);

	bfr new_net_1633_bfr_after (
		.din(new_net_1632),
		.dout(new_net_1633)
	);

	bfr new_net_1634_bfr_after (
		.din(new_net_1633),
		.dout(new_net_1634)
	);

	bfr new_net_1635_bfr_after (
		.din(new_net_1634),
		.dout(new_net_1635)
	);

	bfr new_net_1636_bfr_after (
		.din(new_net_1635),
		.dout(new_net_1636)
	);

	bfr new_net_1637_bfr_after (
		.din(new_net_1636),
		.dout(new_net_1637)
	);

	bfr new_net_1638_bfr_after (
		.din(new_net_1637),
		.dout(new_net_1638)
	);

	bfr new_net_1639_bfr_after (
		.din(new_net_1638),
		.dout(new_net_1639)
	);

	bfr new_net_1640_bfr_after (
		.din(new_net_1639),
		.dout(new_net_1640)
	);

	bfr new_net_1641_bfr_after (
		.din(new_net_1640),
		.dout(new_net_1641)
	);

	bfr new_net_1642_bfr_after (
		.din(new_net_1641),
		.dout(new_net_1642)
	);

	bfr new_net_1643_bfr_after (
		.din(new_net_1642),
		.dout(new_net_1643)
	);

	bfr new_net_1644_bfr_after (
		.din(new_net_1643),
		.dout(new_net_1644)
	);

	bfr new_net_1645_bfr_after (
		.din(new_net_1644),
		.dout(new_net_1645)
	);

	bfr new_net_1646_bfr_after (
		.din(new_net_1645),
		.dout(new_net_1646)
	);

	bfr new_net_1647_bfr_after (
		.din(new_net_1646),
		.dout(new_net_1647)
	);

	bfr new_net_1648_bfr_after (
		.din(new_net_1647),
		.dout(new_net_1648)
	);

	bfr new_net_1649_bfr_after (
		.din(new_net_1648),
		.dout(new_net_1649)
	);

	bfr new_net_1650_bfr_after (
		.din(new_net_1649),
		.dout(new_net_1650)
	);

	bfr new_net_1651_bfr_after (
		.din(new_net_1650),
		.dout(new_net_1651)
	);

	bfr new_net_1652_bfr_after (
		.din(new_net_1651),
		.dout(new_net_1652)
	);

	bfr new_net_1653_bfr_after (
		.din(new_net_1652),
		.dout(new_net_1653)
	);

	bfr new_net_1654_bfr_after (
		.din(new_net_1653),
		.dout(new_net_1654)
	);

	bfr new_net_1655_bfr_after (
		.din(new_net_1654),
		.dout(new_net_1655)
	);

	bfr new_net_1656_bfr_after (
		.din(new_net_1655),
		.dout(new_net_1656)
	);

	bfr new_net_1657_bfr_after (
		.din(new_net_1656),
		.dout(new_net_1657)
	);

	bfr new_net_1658_bfr_after (
		.din(new_net_1657),
		.dout(new_net_1658)
	);

	bfr new_net_1659_bfr_after (
		.din(new_net_1658),
		.dout(new_net_1659)
	);

	bfr new_net_1660_bfr_after (
		.din(new_net_1659),
		.dout(new_net_1660)
	);

	bfr new_net_1661_bfr_after (
		.din(new_net_1660),
		.dout(new_net_1661)
	);

	bfr new_net_1662_bfr_after (
		.din(new_net_1661),
		.dout(new_net_1662)
	);

	bfr new_net_1663_bfr_after (
		.din(new_net_1662),
		.dout(new_net_1663)
	);

	bfr new_net_1664_bfr_after (
		.din(new_net_1663),
		.dout(new_net_1664)
	);

	bfr new_net_1665_bfr_after (
		.din(new_net_1664),
		.dout(new_net_1665)
	);

	bfr new_net_1666_bfr_after (
		.din(new_net_1665),
		.dout(new_net_1666)
	);

	bfr new_net_1667_bfr_after (
		.din(new_net_1666),
		.dout(new_net_1667)
	);

	bfr N421_bfr_after (
		.din(new_net_1667),
		.dout(N421)
	);

	bfr new_net_1668_bfr_after (
		.din(new_net_536),
		.dout(new_net_1668)
	);

	bfr new_net_1669_bfr_after (
		.din(new_net_1668),
		.dout(new_net_1669)
	);

	bfr new_net_1670_bfr_after (
		.din(new_net_1669),
		.dout(new_net_1670)
	);

	bfr new_net_1671_bfr_after (
		.din(new_net_1670),
		.dout(new_net_1671)
	);

	bfr new_net_1672_bfr_after (
		.din(new_net_1671),
		.dout(new_net_1672)
	);

	bfr new_net_1673_bfr_after (
		.din(new_net_1672),
		.dout(new_net_1673)
	);

	bfr new_net_1674_bfr_after (
		.din(new_net_1673),
		.dout(new_net_1674)
	);

	bfr new_net_1675_bfr_after (
		.din(new_net_1674),
		.dout(new_net_1675)
	);

	bfr new_net_1676_bfr_after (
		.din(new_net_1675),
		.dout(new_net_1676)
	);

	bfr new_net_1677_bfr_after (
		.din(new_net_1676),
		.dout(new_net_1677)
	);

	bfr new_net_1678_bfr_after (
		.din(new_net_1677),
		.dout(new_net_1678)
	);

	bfr new_net_1679_bfr_after (
		.din(new_net_1678),
		.dout(new_net_1679)
	);

	bfr new_net_1680_bfr_after (
		.din(new_net_1679),
		.dout(new_net_1680)
	);

	bfr new_net_1681_bfr_after (
		.din(new_net_1680),
		.dout(new_net_1681)
	);

	bfr new_net_1682_bfr_after (
		.din(new_net_1681),
		.dout(new_net_1682)
	);

	bfr new_net_1683_bfr_after (
		.din(new_net_1682),
		.dout(new_net_1683)
	);

	bfr new_net_1684_bfr_after (
		.din(new_net_1683),
		.dout(new_net_1684)
	);

	bfr new_net_1685_bfr_after (
		.din(new_net_1684),
		.dout(new_net_1685)
	);

	bfr new_net_1686_bfr_after (
		.din(new_net_1685),
		.dout(new_net_1686)
	);

	bfr new_net_1687_bfr_after (
		.din(new_net_1686),
		.dout(new_net_1687)
	);

	bfr new_net_1688_bfr_after (
		.din(new_net_1687),
		.dout(new_net_1688)
	);

	bfr new_net_1689_bfr_after (
		.din(new_net_1688),
		.dout(new_net_1689)
	);

	bfr new_net_1690_bfr_after (
		.din(new_net_1689),
		.dout(new_net_1690)
	);

	bfr new_net_1691_bfr_after (
		.din(new_net_1690),
		.dout(new_net_1691)
	);

	bfr new_net_1692_bfr_after (
		.din(new_net_1691),
		.dout(new_net_1692)
	);

	bfr new_net_1693_bfr_after (
		.din(new_net_1692),
		.dout(new_net_1693)
	);

	bfr new_net_1694_bfr_after (
		.din(new_net_1693),
		.dout(new_net_1694)
	);

	bfr new_net_1695_bfr_after (
		.din(new_net_1694),
		.dout(new_net_1695)
	);

	bfr new_net_1696_bfr_after (
		.din(new_net_1695),
		.dout(new_net_1696)
	);

	bfr new_net_1697_bfr_after (
		.din(new_net_1696),
		.dout(new_net_1697)
	);

	bfr new_net_1698_bfr_after (
		.din(new_net_1697),
		.dout(new_net_1698)
	);

	bfr new_net_1699_bfr_after (
		.din(new_net_1698),
		.dout(new_net_1699)
	);

	bfr new_net_1700_bfr_after (
		.din(new_net_1699),
		.dout(new_net_1700)
	);

	bfr new_net_1701_bfr_after (
		.din(new_net_1700),
		.dout(new_net_1701)
	);

	bfr N447_bfr_after (
		.din(new_net_1701),
		.dout(N447)
	);

	bfr new_net_1702_bfr_after (
		.din(new_net_548),
		.dout(new_net_1702)
	);

	bfr new_net_1703_bfr_after (
		.din(new_net_1702),
		.dout(new_net_1703)
	);

	bfr N879_bfr_after (
		.din(new_net_1703),
		.dout(N879)
	);

	bfr new_net_1704_bfr_after (
		.din(new_net_560),
		.dout(new_net_1704)
	);

	bfr new_net_1705_bfr_after (
		.din(new_net_1704),
		.dout(new_net_1705)
	);

	bfr new_net_1706_bfr_after (
		.din(new_net_1705),
		.dout(new_net_1706)
	);

	bfr new_net_1707_bfr_after (
		.din(new_net_1706),
		.dout(new_net_1707)
	);

	bfr new_net_1708_bfr_after (
		.din(new_net_1707),
		.dout(new_net_1708)
	);

	bfr new_net_1709_bfr_after (
		.din(new_net_1708),
		.dout(new_net_1709)
	);

	bfr new_net_1710_bfr_after (
		.din(new_net_1709),
		.dout(new_net_1710)
	);

	bfr new_net_1711_bfr_after (
		.din(new_net_1710),
		.dout(new_net_1711)
	);

	bfr new_net_1712_bfr_after (
		.din(new_net_1711),
		.dout(new_net_1712)
	);

	bfr new_net_1713_bfr_after (
		.din(new_net_1712),
		.dout(new_net_1713)
	);

	bfr new_net_1714_bfr_after (
		.din(new_net_1713),
		.dout(new_net_1714)
	);

	bfr new_net_1715_bfr_after (
		.din(new_net_1714),
		.dout(new_net_1715)
	);

	bfr new_net_1716_bfr_after (
		.din(new_net_1715),
		.dout(new_net_1716)
	);

	bfr new_net_1717_bfr_after (
		.din(new_net_1716),
		.dout(new_net_1717)
	);

	bfr new_net_1718_bfr_after (
		.din(new_net_1717),
		.dout(new_net_1718)
	);

	bfr new_net_1719_bfr_after (
		.din(new_net_1718),
		.dout(new_net_1719)
	);

	bfr new_net_1720_bfr_after (
		.din(new_net_1719),
		.dout(new_net_1720)
	);

	bfr new_net_1721_bfr_after (
		.din(new_net_1720),
		.dout(new_net_1721)
	);

	bfr new_net_1722_bfr_after (
		.din(new_net_1721),
		.dout(new_net_1722)
	);

	bfr new_net_1723_bfr_after (
		.din(new_net_1722),
		.dout(new_net_1723)
	);

	bfr new_net_1724_bfr_after (
		.din(new_net_1723),
		.dout(new_net_1724)
	);

	bfr new_net_1725_bfr_after (
		.din(new_net_1724),
		.dout(new_net_1725)
	);

	bfr new_net_1726_bfr_after (
		.din(new_net_1725),
		.dout(new_net_1726)
	);

	bfr new_net_1727_bfr_after (
		.din(new_net_1726),
		.dout(new_net_1727)
	);

	bfr new_net_1728_bfr_after (
		.din(new_net_1727),
		.dout(new_net_1728)
	);

	bfr new_net_1729_bfr_after (
		.din(new_net_1728),
		.dout(new_net_1729)
	);

	bfr new_net_1730_bfr_after (
		.din(new_net_1729),
		.dout(new_net_1730)
	);

	bfr new_net_1731_bfr_after (
		.din(new_net_1730),
		.dout(new_net_1731)
	);

	bfr N768_bfr_after (
		.din(new_net_1731),
		.dout(N768)
	);

	bfr new_net_464_bfr_after (
		.din(_076_),
		.dout(new_net_464)
	);

	bfr new_net_456_bfr_after (
		.din(_022_),
		.dout(new_net_456)
	);

	bfr new_net_1732_bfr_after (
		.din(N73),
		.dout(new_net_1732)
	);

	bfr new_net_460_bfr_after (
		.din(new_net_1732),
		.dout(new_net_460)
	);

	bfr new_net_1733_bfr_after (
		.din(_137_),
		.dout(new_net_1733)
	);

	bfr new_net_1734_bfr_after (
		.din(new_net_1733),
		.dout(new_net_1734)
	);

	bfr new_net_1735_bfr_after (
		.din(new_net_1734),
		.dout(new_net_1735)
	);

	bfr new_net_1736_bfr_after (
		.din(new_net_1735),
		.dout(new_net_1736)
	);

	bfr new_net_1737_bfr_after (
		.din(new_net_1736),
		.dout(new_net_1737)
	);

	bfr new_net_1738_bfr_after (
		.din(new_net_1737),
		.dout(new_net_1738)
	);

	bfr new_net_1739_bfr_after (
		.din(new_net_1738),
		.dout(new_net_1739)
	);

	bfr new_net_1740_bfr_after (
		.din(new_net_1739),
		.dout(new_net_1740)
	);

	bfr new_net_1741_bfr_after (
		.din(new_net_1740),
		.dout(new_net_1741)
	);

	bfr new_net_1742_bfr_after (
		.din(new_net_1741),
		.dout(new_net_1742)
	);

	bfr new_net_1743_bfr_after (
		.din(new_net_1742),
		.dout(new_net_1743)
	);

	bfr new_net_1744_bfr_after (
		.din(new_net_1743),
		.dout(new_net_1744)
	);

	bfr new_net_1745_bfr_after (
		.din(new_net_1744),
		.dout(new_net_1745)
	);

	bfr new_net_1746_bfr_after (
		.din(new_net_1745),
		.dout(new_net_1746)
	);

	bfr new_net_1747_bfr_after (
		.din(new_net_1746),
		.dout(new_net_1747)
	);

	bfr new_net_1748_bfr_after (
		.din(new_net_1747),
		.dout(new_net_1748)
	);

	bfr new_net_1749_bfr_after (
		.din(new_net_1748),
		.dout(new_net_1749)
	);

	bfr new_net_481_bfr_after (
		.din(new_net_1749),
		.dout(new_net_481)
	);

	bfr new_net_502_bfr_after (
		.din(_191_),
		.dout(new_net_502)
	);

	bfr new_net_485_bfr_after (
		.din(_149_),
		.dout(new_net_485)
	);

	bfr new_net_506_bfr_after (
		.din(_196_),
		.dout(new_net_506)
	);

	bfr new_net_1750_bfr_after (
		.din(_132_),
		.dout(new_net_1750)
	);

	bfr new_net_1751_bfr_after (
		.din(new_net_1750),
		.dout(new_net_1751)
	);

	bfr new_net_1752_bfr_after (
		.din(new_net_1751),
		.dout(new_net_1752)
	);

	bfr new_net_1753_bfr_after (
		.din(new_net_1752),
		.dout(new_net_1753)
	);

	bfr new_net_1754_bfr_after (
		.din(new_net_1753),
		.dout(new_net_1754)
	);

	bfr new_net_477_bfr_after (
		.din(new_net_1754),
		.dout(new_net_477)
	);

	bfr new_net_498_bfr_after (
		.din(_180_),
		.dout(new_net_498)
	);

	bfr new_net_1755_bfr_after (
		.din(N89),
		.dout(new_net_1755)
	);

	bfr new_net_519_bfr_after (
		.din(new_net_1755),
		.dout(new_net_519)
	);

	bfr new_net_1756_bfr_after (
		.din(new_net_538),
		.dout(new_net_1756)
	);

	bfr new_net_1757_bfr_after (
		.din(new_net_1756),
		.dout(new_net_1757)
	);

	bfr new_net_1758_bfr_after (
		.din(new_net_1757),
		.dout(new_net_1758)
	);

	bfr new_net_1759_bfr_after (
		.din(new_net_1758),
		.dout(new_net_1759)
	);

	bfr new_net_1760_bfr_after (
		.din(new_net_1759),
		.dout(new_net_1760)
	);

	bfr new_net_1761_bfr_after (
		.din(new_net_1760),
		.dout(new_net_1761)
	);

	bfr new_net_1762_bfr_after (
		.din(new_net_1761),
		.dout(new_net_1762)
	);

	bfr new_net_1763_bfr_after (
		.din(new_net_1762),
		.dout(new_net_1763)
	);

	bfr new_net_1764_bfr_after (
		.din(new_net_1763),
		.dout(new_net_1764)
	);

	bfr new_net_1765_bfr_after (
		.din(new_net_1764),
		.dout(new_net_1765)
	);

	bfr new_net_1766_bfr_after (
		.din(new_net_1765),
		.dout(new_net_1766)
	);

	bfr new_net_1767_bfr_after (
		.din(new_net_1766),
		.dout(new_net_1767)
	);

	bfr new_net_1768_bfr_after (
		.din(new_net_1767),
		.dout(new_net_1768)
	);

	bfr new_net_1769_bfr_after (
		.din(new_net_1768),
		.dout(new_net_1769)
	);

	bfr new_net_1770_bfr_after (
		.din(new_net_1769),
		.dout(new_net_1770)
	);

	bfr new_net_1771_bfr_after (
		.din(new_net_1770),
		.dout(new_net_1771)
	);

	bfr new_net_1772_bfr_after (
		.din(new_net_1771),
		.dout(new_net_1772)
	);

	bfr new_net_1773_bfr_after (
		.din(new_net_1772),
		.dout(new_net_1773)
	);

	bfr new_net_1774_bfr_after (
		.din(new_net_1773),
		.dout(new_net_1774)
	);

	bfr new_net_1775_bfr_after (
		.din(new_net_1774),
		.dout(new_net_1775)
	);

	bfr new_net_1776_bfr_after (
		.din(new_net_1775),
		.dout(new_net_1776)
	);

	bfr new_net_1777_bfr_after (
		.din(new_net_1776),
		.dout(new_net_1777)
	);

	bfr new_net_1778_bfr_after (
		.din(new_net_1777),
		.dout(new_net_1778)
	);

	bfr new_net_1779_bfr_after (
		.din(new_net_1778),
		.dout(new_net_1779)
	);

	bfr new_net_1780_bfr_after (
		.din(new_net_1779),
		.dout(new_net_1780)
	);

	bfr new_net_1781_bfr_after (
		.din(new_net_1780),
		.dout(new_net_1781)
	);

	bfr new_net_1782_bfr_after (
		.din(new_net_1781),
		.dout(new_net_1782)
	);

	bfr new_net_1783_bfr_after (
		.din(new_net_1782),
		.dout(new_net_1783)
	);

	bfr new_net_1784_bfr_after (
		.din(new_net_1783),
		.dout(new_net_1784)
	);

	bfr new_net_1785_bfr_after (
		.din(new_net_1784),
		.dout(new_net_1785)
	);

	bfr new_net_1786_bfr_after (
		.din(new_net_1785),
		.dout(new_net_1786)
	);

	bfr new_net_1787_bfr_after (
		.din(new_net_1786),
		.dout(new_net_1787)
	);

	bfr new_net_1788_bfr_after (
		.din(new_net_1787),
		.dout(new_net_1788)
	);

	bfr new_net_1789_bfr_after (
		.din(new_net_1788),
		.dout(new_net_1789)
	);

	bfr new_net_1790_bfr_after (
		.din(new_net_1789),
		.dout(new_net_1790)
	);

	bfr new_net_1791_bfr_after (
		.din(new_net_1790),
		.dout(new_net_1791)
	);

	bfr new_net_1792_bfr_after (
		.din(new_net_1791),
		.dout(new_net_1792)
	);

	bfr N450_bfr_after (
		.din(new_net_1792),
		.dout(N450)
	);

	bfr new_net_1793_bfr_after (
		.din(new_net_562),
		.dout(new_net_1793)
	);

	bfr new_net_1794_bfr_after (
		.din(new_net_1793),
		.dout(new_net_1794)
	);

	bfr new_net_1795_bfr_after (
		.din(new_net_1794),
		.dout(new_net_1795)
	);

	bfr new_net_1796_bfr_after (
		.din(new_net_1795),
		.dout(new_net_1796)
	);

	bfr new_net_1797_bfr_after (
		.din(new_net_1796),
		.dout(new_net_1797)
	);

	bfr new_net_1798_bfr_after (
		.din(new_net_1797),
		.dout(new_net_1798)
	);

	bfr new_net_1799_bfr_after (
		.din(new_net_1798),
		.dout(new_net_1799)
	);

	bfr new_net_1800_bfr_after (
		.din(new_net_1799),
		.dout(new_net_1800)
	);

	bfr new_net_1801_bfr_after (
		.din(new_net_1800),
		.dout(new_net_1801)
	);

	bfr new_net_1802_bfr_after (
		.din(new_net_1801),
		.dout(new_net_1802)
	);

	bfr new_net_1803_bfr_after (
		.din(new_net_1802),
		.dout(new_net_1803)
	);

	bfr new_net_1804_bfr_after (
		.din(new_net_1803),
		.dout(new_net_1804)
	);

	bfr new_net_1805_bfr_after (
		.din(new_net_1804),
		.dout(new_net_1805)
	);

	bfr new_net_1806_bfr_after (
		.din(new_net_1805),
		.dout(new_net_1806)
	);

	bfr new_net_1807_bfr_after (
		.din(new_net_1806),
		.dout(new_net_1807)
	);

	bfr new_net_1808_bfr_after (
		.din(new_net_1807),
		.dout(new_net_1808)
	);

	bfr new_net_1809_bfr_after (
		.din(new_net_1808),
		.dout(new_net_1809)
	);

	bfr new_net_1810_bfr_after (
		.din(new_net_1809),
		.dout(new_net_1810)
	);

	bfr new_net_1811_bfr_after (
		.din(new_net_1810),
		.dout(new_net_1811)
	);

	bfr new_net_1812_bfr_after (
		.din(new_net_1811),
		.dout(new_net_1812)
	);

	bfr new_net_1813_bfr_after (
		.din(new_net_1812),
		.dout(new_net_1813)
	);

	bfr new_net_1814_bfr_after (
		.din(new_net_1813),
		.dout(new_net_1814)
	);

	bfr new_net_1815_bfr_after (
		.din(new_net_1814),
		.dout(new_net_1815)
	);

	bfr new_net_1816_bfr_after (
		.din(new_net_1815),
		.dout(new_net_1816)
	);

	bfr new_net_1817_bfr_after (
		.din(new_net_1816),
		.dout(new_net_1817)
	);

	bfr new_net_1818_bfr_after (
		.din(new_net_1817),
		.dout(new_net_1818)
	);

	bfr new_net_1819_bfr_after (
		.din(new_net_1818),
		.dout(new_net_1819)
	);

	bfr new_net_1820_bfr_after (
		.din(new_net_1819),
		.dout(new_net_1820)
	);

	bfr new_net_1821_bfr_after (
		.din(new_net_1820),
		.dout(new_net_1821)
	);

	bfr new_net_1822_bfr_after (
		.din(new_net_1821),
		.dout(new_net_1822)
	);

	bfr new_net_1823_bfr_after (
		.din(new_net_1822),
		.dout(new_net_1823)
	);

	bfr new_net_1824_bfr_after (
		.din(new_net_1823),
		.dout(new_net_1824)
	);

	bfr new_net_1825_bfr_after (
		.din(new_net_1824),
		.dout(new_net_1825)
	);

	bfr new_net_1826_bfr_after (
		.din(new_net_1825),
		.dout(new_net_1826)
	);

	bfr new_net_1827_bfr_after (
		.din(new_net_1826),
		.dout(new_net_1827)
	);

	bfr new_net_1828_bfr_after (
		.din(new_net_1827),
		.dout(new_net_1828)
	);

	bfr N420_bfr_after (
		.din(new_net_1828),
		.dout(N420)
	);

	bfr new_net_1829_bfr_after (
		.din(_276_),
		.dout(new_net_1829)
	);

	bfr new_net_450_bfr_after (
		.din(new_net_1829),
		.dout(new_net_450)
	);

	bfr new_net_1830_bfr_after (
		.din(_162_),
		.dout(new_net_1830)
	);

	bfr new_net_1831_bfr_after (
		.din(new_net_1830),
		.dout(new_net_1831)
	);

	bfr new_net_1832_bfr_after (
		.din(new_net_1831),
		.dout(new_net_1832)
	);

	bfr new_net_1833_bfr_after (
		.din(new_net_1832),
		.dout(new_net_1833)
	);

	bfr new_net_1834_bfr_after (
		.din(new_net_1833),
		.dout(new_net_1834)
	);

	bfr new_net_489_bfr_after (
		.din(new_net_1834),
		.dout(new_net_489)
	);

	bfr new_net_1835_bfr_after (
		.din(_209_),
		.dout(new_net_1835)
	);

	bfr new_net_1836_bfr_after (
		.din(new_net_1835),
		.dout(new_net_1836)
	);

	bfr new_net_1837_bfr_after (
		.din(new_net_1836),
		.dout(new_net_1837)
	);

	bfr new_net_1838_bfr_after (
		.din(new_net_1837),
		.dout(new_net_1838)
	);

	bfr new_net_510_bfr_after (
		.din(new_net_1838),
		.dout(new_net_510)
	);

	bfr new_net_1839_bfr_after (
		.din(_090_),
		.dout(new_net_1839)
	);

	bfr new_net_1840_bfr_after (
		.din(new_net_1839),
		.dout(new_net_1840)
	);

	bfr new_net_1841_bfr_after (
		.din(new_net_1840),
		.dout(new_net_1841)
	);

	bfr new_net_1842_bfr_after (
		.din(new_net_1841),
		.dout(new_net_1842)
	);

	bfr new_net_1843_bfr_after (
		.din(new_net_1842),
		.dout(new_net_1843)
	);

	bfr new_net_1844_bfr_after (
		.din(new_net_1843),
		.dout(new_net_1844)
	);

	bfr new_net_468_bfr_after (
		.din(new_net_1844),
		.dout(new_net_468)
	);

	bfr new_net_1845_bfr_after (
		.din(_120_),
		.dout(new_net_1845)
	);

	bfr new_net_1846_bfr_after (
		.din(new_net_1845),
		.dout(new_net_1846)
	);

	bfr new_net_1847_bfr_after (
		.din(new_net_1846),
		.dout(new_net_1847)
	);

	bfr new_net_472_bfr_after (
		.din(new_net_1847),
		.dout(new_net_472)
	);

	bfr new_net_493_bfr_after (
		.din(N259),
		.dout(new_net_493)
	);

	bfr new_net_1848_bfr_after (
		.din(_213_),
		.dout(new_net_1848)
	);

	bfr new_net_514_bfr_after (
		.din(new_net_1848),
		.dout(new_net_514)
	);

	bfr new_net_1849_bfr_after (
		.din(new_net_542),
		.dout(new_net_1849)
	);

	bfr new_net_1850_bfr_after (
		.din(new_net_1849),
		.dout(new_net_1850)
	);

	bfr new_net_1851_bfr_after (
		.din(new_net_1850),
		.dout(new_net_1851)
	);

	bfr new_net_1852_bfr_after (
		.din(new_net_1851),
		.dout(new_net_1852)
	);

	bfr new_net_1853_bfr_after (
		.din(new_net_1852),
		.dout(new_net_1853)
	);

	bfr new_net_1854_bfr_after (
		.din(new_net_1853),
		.dout(new_net_1854)
	);

	bfr new_net_1855_bfr_after (
		.din(new_net_1854),
		.dout(new_net_1855)
	);

	bfr new_net_1856_bfr_after (
		.din(new_net_1855),
		.dout(new_net_1856)
	);

	bfr N874_bfr_after (
		.din(new_net_1856),
		.dout(N874)
	);

	bfr new_net_1857_bfr_after (
		.din(new_net_566),
		.dout(new_net_1857)
	);

	bfr N866_bfr_after (
		.din(new_net_1857),
		.dout(N866)
	);

	bfr new_net_448_bfr_after (
		.din(N26),
		.dout(new_net_448)
	);

	bfr new_net_480_bfr_after (
		.din(_136_),
		.dout(new_net_480)
	);

	bfr new_net_501_bfr_after (
		.din(N267),
		.dout(new_net_501)
	);

	bfr new_net_1858_bfr_after (
		.din(_007_),
		.dout(new_net_1858)
	);

	bfr new_net_1859_bfr_after (
		.din(new_net_1858),
		.dout(new_net_1859)
	);

	bfr new_net_1860_bfr_after (
		.din(new_net_1859),
		.dout(new_net_1860)
	);

	bfr new_net_1861_bfr_after (
		.din(new_net_1860),
		.dout(new_net_1861)
	);

	bfr new_net_1862_bfr_after (
		.din(new_net_1861),
		.dout(new_net_1862)
	);

	bfr new_net_1863_bfr_after (
		.din(new_net_1862),
		.dout(new_net_1863)
	);

	bfr new_net_455_bfr_after (
		.din(new_net_1863),
		.dout(new_net_455)
	);

	bfr new_net_459_bfr_after (
		.din(N72),
		.dout(new_net_459)
	);

	bfr new_net_1864_bfr_after (
		.din(_075_),
		.dout(new_net_1864)
	);

	bfr new_net_1865_bfr_after (
		.din(new_net_1864),
		.dout(new_net_1865)
	);

	bfr new_net_1866_bfr_after (
		.din(new_net_1865),
		.dout(new_net_1866)
	);

	bfr new_net_463_bfr_after (
		.din(new_net_1866),
		.dout(new_net_463)
	);

	bfr new_net_1867_bfr_after (
		.din(_148_),
		.dout(new_net_1867)
	);

	bfr new_net_1868_bfr_after (
		.din(new_net_1867),
		.dout(new_net_1868)
	);

	bfr new_net_1869_bfr_after (
		.din(new_net_1868),
		.dout(new_net_1869)
	);

	bfr new_net_484_bfr_after (
		.din(new_net_1869),
		.dout(new_net_484)
	);

	bfr new_net_505_bfr_after (
		.din(_195_),
		.dout(new_net_505)
	);

	bfr new_net_1870_bfr_after (
		.din(new_net_526),
		.dout(new_net_1870)
	);

	bfr new_net_1871_bfr_after (
		.din(new_net_1870),
		.dout(new_net_1871)
	);

	bfr new_net_1872_bfr_after (
		.din(new_net_1871),
		.dout(new_net_1872)
	);

	bfr new_net_1873_bfr_after (
		.din(new_net_1872),
		.dout(new_net_1873)
	);

	bfr new_net_1874_bfr_after (
		.din(new_net_1873),
		.dout(new_net_1874)
	);

	bfr new_net_1875_bfr_after (
		.din(new_net_1874),
		.dout(new_net_1875)
	);

	bfr new_net_1876_bfr_after (
		.din(new_net_1875),
		.dout(new_net_1876)
	);

	bfr new_net_1877_bfr_after (
		.din(new_net_1876),
		.dout(new_net_1877)
	);

	bfr new_net_1878_bfr_after (
		.din(new_net_1877),
		.dout(new_net_1878)
	);

	bfr new_net_1879_bfr_after (
		.din(new_net_1878),
		.dout(new_net_1879)
	);

	bfr new_net_1880_bfr_after (
		.din(new_net_1879),
		.dout(new_net_1880)
	);

	bfr new_net_1881_bfr_after (
		.din(new_net_1880),
		.dout(new_net_1881)
	);

	bfr new_net_1882_bfr_after (
		.din(new_net_1881),
		.dout(new_net_1882)
	);

	bfr new_net_1883_bfr_after (
		.din(new_net_1882),
		.dout(new_net_1883)
	);

	bfr new_net_1884_bfr_after (
		.din(new_net_1883),
		.dout(new_net_1884)
	);

	bfr new_net_1885_bfr_after (
		.din(new_net_1884),
		.dout(new_net_1885)
	);

	bfr new_net_1886_bfr_after (
		.din(new_net_1885),
		.dout(new_net_1886)
	);

	bfr new_net_1887_bfr_after (
		.din(new_net_1886),
		.dout(new_net_1887)
	);

	bfr new_net_1888_bfr_after (
		.din(new_net_1887),
		.dout(new_net_1888)
	);

	bfr new_net_1889_bfr_after (
		.din(new_net_1888),
		.dout(new_net_1889)
	);

	bfr new_net_1890_bfr_after (
		.din(new_net_1889),
		.dout(new_net_1890)
	);

	bfr new_net_1891_bfr_after (
		.din(new_net_1890),
		.dout(new_net_1891)
	);

	bfr new_net_1892_bfr_after (
		.din(new_net_1891),
		.dout(new_net_1892)
	);

	bfr new_net_1893_bfr_after (
		.din(new_net_1892),
		.dout(new_net_1893)
	);

	bfr new_net_1894_bfr_after (
		.din(new_net_1893),
		.dout(new_net_1894)
	);

	bfr new_net_1895_bfr_after (
		.din(new_net_1894),
		.dout(new_net_1895)
	);

	bfr new_net_1896_bfr_after (
		.din(new_net_1895),
		.dout(new_net_1896)
	);

	bfr new_net_1897_bfr_after (
		.din(new_net_1896),
		.dout(new_net_1897)
	);

	bfr new_net_1898_bfr_after (
		.din(new_net_1897),
		.dout(new_net_1898)
	);

	bfr new_net_1899_bfr_after (
		.din(new_net_1898),
		.dout(new_net_1899)
	);

	bfr new_net_1900_bfr_after (
		.din(new_net_1899),
		.dout(new_net_1900)
	);

	bfr new_net_1901_bfr_after (
		.din(new_net_1900),
		.dout(new_net_1901)
	);

	bfr new_net_1902_bfr_after (
		.din(new_net_1901),
		.dout(new_net_1902)
	);

	bfr new_net_1903_bfr_after (
		.din(new_net_1902),
		.dout(new_net_1903)
	);

	bfr new_net_1904_bfr_after (
		.din(new_net_1903),
		.dout(new_net_1904)
	);

	bfr new_net_1905_bfr_after (
		.din(new_net_1904),
		.dout(new_net_1905)
	);

	bfr new_net_1906_bfr_after (
		.din(new_net_1905),
		.dout(new_net_1906)
	);

	bfr new_net_1907_bfr_after (
		.din(new_net_1906),
		.dout(new_net_1907)
	);

	bfr new_net_1908_bfr_after (
		.din(new_net_1907),
		.dout(new_net_1908)
	);

	bfr N391_bfr_after (
		.din(new_net_1908),
		.dout(N391)
	);

	bfr new_net_476_bfr_after (
		.din(_125_),
		.dout(new_net_476)
	);

	bfr new_net_497_bfr_after (
		.din(_179_),
		.dout(new_net_497)
	);

	bfr new_net_1909_bfr_after (
		.din(new_net_520),
		.dout(new_net_1909)
	);

	bfr new_net_1910_bfr_after (
		.din(new_net_1909),
		.dout(new_net_1910)
	);

	bfr new_net_1911_bfr_after (
		.din(new_net_1910),
		.dout(new_net_1911)
	);

	bfr new_net_1912_bfr_after (
		.din(new_net_1911),
		.dout(new_net_1912)
	);

	bfr new_net_1913_bfr_after (
		.din(new_net_1912),
		.dout(new_net_1913)
	);

	bfr new_net_1914_bfr_after (
		.din(new_net_1913),
		.dout(new_net_1914)
	);

	bfr new_net_1915_bfr_after (
		.din(new_net_1914),
		.dout(new_net_1915)
	);

	bfr new_net_1916_bfr_after (
		.din(new_net_1915),
		.dout(new_net_1916)
	);

	bfr new_net_1917_bfr_after (
		.din(new_net_1916),
		.dout(new_net_1917)
	);

	bfr new_net_1918_bfr_after (
		.din(new_net_1917),
		.dout(new_net_1918)
	);

	bfr new_net_1919_bfr_after (
		.din(new_net_1918),
		.dout(new_net_1919)
	);

	bfr new_net_1920_bfr_after (
		.din(new_net_1919),
		.dout(new_net_1920)
	);

	bfr new_net_1921_bfr_after (
		.din(new_net_1920),
		.dout(new_net_1921)
	);

	bfr new_net_1922_bfr_after (
		.din(new_net_1921),
		.dout(new_net_1922)
	);

	bfr new_net_1923_bfr_after (
		.din(new_net_1922),
		.dout(new_net_1923)
	);

	bfr new_net_1924_bfr_after (
		.din(new_net_1923),
		.dout(new_net_1924)
	);

	bfr new_net_1925_bfr_after (
		.din(new_net_1924),
		.dout(new_net_1925)
	);

	bfr new_net_1926_bfr_after (
		.din(new_net_1925),
		.dout(new_net_1926)
	);

	bfr new_net_1927_bfr_after (
		.din(new_net_1926),
		.dout(new_net_1927)
	);

	bfr new_net_1928_bfr_after (
		.din(new_net_1927),
		.dout(new_net_1928)
	);

	bfr new_net_1929_bfr_after (
		.din(new_net_1928),
		.dout(new_net_1929)
	);

	bfr new_net_1930_bfr_after (
		.din(new_net_1929),
		.dout(new_net_1930)
	);

	bfr new_net_1931_bfr_after (
		.din(new_net_1930),
		.dout(new_net_1931)
	);

	bfr new_net_1932_bfr_after (
		.din(new_net_1931),
		.dout(new_net_1932)
	);

	bfr new_net_1933_bfr_after (
		.din(new_net_1932),
		.dout(new_net_1933)
	);

	bfr new_net_1934_bfr_after (
		.din(new_net_1933),
		.dout(new_net_1934)
	);

	bfr new_net_1935_bfr_after (
		.din(new_net_1934),
		.dout(new_net_1935)
	);

	bfr new_net_1936_bfr_after (
		.din(new_net_1935),
		.dout(new_net_1936)
	);

	bfr N767_bfr_after (
		.din(new_net_1936),
		.dout(N767)
	);

	bfr new_net_1937_bfr_after (
		.din(new_net_532),
		.dout(new_net_1937)
	);

	bfr new_net_1938_bfr_after (
		.din(new_net_1937),
		.dout(new_net_1938)
	);

	bfr new_net_1939_bfr_after (
		.din(new_net_1938),
		.dout(new_net_1939)
	);

	bfr new_net_1940_bfr_after (
		.din(new_net_1939),
		.dout(new_net_1940)
	);

	bfr new_net_1941_bfr_after (
		.din(new_net_1940),
		.dout(new_net_1941)
	);

	bfr N880_bfr_after (
		.din(new_net_1941),
		.dout(N880)
	);

	bfr new_net_1942_bfr_after (
		.din(new_net_544),
		.dout(new_net_1942)
	);

	bfr new_net_1943_bfr_after (
		.din(new_net_1942),
		.dout(new_net_1943)
	);

	bfr new_net_1944_bfr_after (
		.din(new_net_1943),
		.dout(new_net_1944)
	);

	bfr new_net_1945_bfr_after (
		.din(new_net_1944),
		.dout(new_net_1945)
	);

	bfr new_net_1946_bfr_after (
		.din(new_net_1945),
		.dout(new_net_1946)
	);

	bfr new_net_1947_bfr_after (
		.din(new_net_1946),
		.dout(new_net_1947)
	);

	bfr new_net_1948_bfr_after (
		.din(new_net_1947),
		.dout(new_net_1948)
	);

	bfr new_net_1949_bfr_after (
		.din(new_net_1948),
		.dout(new_net_1949)
	);

	bfr new_net_1950_bfr_after (
		.din(new_net_1949),
		.dout(new_net_1950)
	);

	bfr new_net_1951_bfr_after (
		.din(new_net_1950),
		.dout(new_net_1951)
	);

	bfr new_net_1952_bfr_after (
		.din(new_net_1951),
		.dout(new_net_1952)
	);

	bfr new_net_1953_bfr_after (
		.din(new_net_1952),
		.dout(new_net_1953)
	);

	bfr new_net_1954_bfr_after (
		.din(new_net_1953),
		.dout(new_net_1954)
	);

	bfr new_net_1955_bfr_after (
		.din(new_net_1954),
		.dout(new_net_1955)
	);

	bfr new_net_1956_bfr_after (
		.din(new_net_1955),
		.dout(new_net_1956)
	);

	bfr new_net_1957_bfr_after (
		.din(new_net_1956),
		.dout(new_net_1957)
	);

	bfr new_net_1958_bfr_after (
		.din(new_net_1957),
		.dout(new_net_1958)
	);

	bfr new_net_1959_bfr_after (
		.din(new_net_1958),
		.dout(new_net_1959)
	);

	bfr N850_bfr_after (
		.din(new_net_1959),
		.dout(N850)
	);

	bfr new_net_1960_bfr_after (
		.din(new_net_556),
		.dout(new_net_1960)
	);

	bfr new_net_1961_bfr_after (
		.din(new_net_1960),
		.dout(new_net_1961)
	);

	bfr new_net_1962_bfr_after (
		.din(new_net_1961),
		.dout(new_net_1962)
	);

	bfr new_net_1963_bfr_after (
		.din(new_net_1962),
		.dout(new_net_1963)
	);

	bfr new_net_1964_bfr_after (
		.din(new_net_1963),
		.dout(new_net_1964)
	);

	bfr new_net_1965_bfr_after (
		.din(new_net_1964),
		.dout(new_net_1965)
	);

	bfr new_net_1966_bfr_after (
		.din(new_net_1965),
		.dout(new_net_1966)
	);

	bfr new_net_1967_bfr_after (
		.din(new_net_1966),
		.dout(new_net_1967)
	);

	bfr new_net_1968_bfr_after (
		.din(new_net_1967),
		.dout(new_net_1968)
	);

	bfr new_net_1969_bfr_after (
		.din(new_net_1968),
		.dout(new_net_1969)
	);

	bfr new_net_1970_bfr_after (
		.din(new_net_1969),
		.dout(new_net_1970)
	);

	bfr new_net_1971_bfr_after (
		.din(new_net_1970),
		.dout(new_net_1971)
	);

	bfr new_net_1972_bfr_after (
		.din(new_net_1971),
		.dout(new_net_1972)
	);

	bfr new_net_1973_bfr_after (
		.din(new_net_1972),
		.dout(new_net_1973)
	);

	bfr new_net_1974_bfr_after (
		.din(new_net_1973),
		.dout(new_net_1974)
	);

	bfr new_net_1975_bfr_after (
		.din(new_net_1974),
		.dout(new_net_1975)
	);

	bfr new_net_1976_bfr_after (
		.din(new_net_1975),
		.dout(new_net_1976)
	);

	bfr new_net_1977_bfr_after (
		.din(new_net_1976),
		.dout(new_net_1977)
	);

	bfr new_net_1978_bfr_after (
		.din(new_net_1977),
		.dout(new_net_1978)
	);

	bfr new_net_1979_bfr_after (
		.din(new_net_1978),
		.dout(new_net_1979)
	);

	bfr new_net_1980_bfr_after (
		.din(new_net_1979),
		.dout(new_net_1980)
	);

	bfr new_net_1981_bfr_after (
		.din(new_net_1980),
		.dout(new_net_1981)
	);

	bfr new_net_1982_bfr_after (
		.din(new_net_1981),
		.dout(new_net_1982)
	);

	bfr new_net_1983_bfr_after (
		.din(new_net_1982),
		.dout(new_net_1983)
	);

	bfr new_net_1984_bfr_after (
		.din(new_net_1983),
		.dout(new_net_1984)
	);

	bfr new_net_1985_bfr_after (
		.din(new_net_1984),
		.dout(new_net_1985)
	);

	bfr new_net_1986_bfr_after (
		.din(new_net_1985),
		.dout(new_net_1986)
	);

	bfr new_net_1987_bfr_after (
		.din(new_net_1986),
		.dout(new_net_1987)
	);

	bfr new_net_1988_bfr_after (
		.din(new_net_1987),
		.dout(new_net_1988)
	);

	bfr new_net_1989_bfr_after (
		.din(new_net_1988),
		.dout(new_net_1989)
	);

	bfr new_net_1990_bfr_after (
		.din(new_net_1989),
		.dout(new_net_1990)
	);

	bfr new_net_1991_bfr_after (
		.din(new_net_1990),
		.dout(new_net_1991)
	);

	bfr new_net_1992_bfr_after (
		.din(new_net_1991),
		.dout(new_net_1992)
	);

	bfr N446_bfr_after (
		.din(new_net_1992),
		.dout(N446)
	);

	bfr new_net_449_bfr_after (
		.din(N156),
		.dout(new_net_449)
	);

	bfr new_net_1993_bfr_after (
		.din(_123_),
		.dout(new_net_1993)
	);

	bfr new_net_1994_bfr_after (
		.din(new_net_1993),
		.dout(new_net_1994)
	);

	bfr new_net_1995_bfr_after (
		.din(new_net_1994),
		.dout(new_net_1995)
	);

	bfr new_net_1996_bfr_after (
		.din(new_net_1995),
		.dout(new_net_1996)
	);

	bfr new_net_1997_bfr_after (
		.din(new_net_1996),
		.dout(new_net_1997)
	);

	bfr new_net_1998_bfr_after (
		.din(new_net_1997),
		.dout(new_net_1998)
	);

	bfr new_net_1999_bfr_after (
		.din(new_net_1998),
		.dout(new_net_1999)
	);

	bfr new_net_2000_bfr_after (
		.din(new_net_1999),
		.dout(new_net_2000)
	);

	bfr new_net_2001_bfr_after (
		.din(new_net_2000),
		.dout(new_net_2001)
	);

	bfr new_net_2002_bfr_after (
		.din(new_net_2001),
		.dout(new_net_2002)
	);

	bfr new_net_2003_bfr_after (
		.din(new_net_2002),
		.dout(new_net_2003)
	);

	bfr new_net_2004_bfr_after (
		.din(new_net_2003),
		.dout(new_net_2004)
	);

	bfr new_net_2005_bfr_after (
		.din(new_net_2004),
		.dout(new_net_2005)
	);

	bfr new_net_2006_bfr_after (
		.din(new_net_2005),
		.dout(new_net_2006)
	);

	bfr new_net_2007_bfr_after (
		.din(new_net_2006),
		.dout(new_net_2007)
	);

	bfr new_net_2008_bfr_after (
		.din(new_net_2007),
		.dout(new_net_2008)
	);

	bfr new_net_2009_bfr_after (
		.din(new_net_2008),
		.dout(new_net_2009)
	);

	bfr new_net_2010_bfr_after (
		.din(new_net_2009),
		.dout(new_net_2010)
	);

	bfr new_net_2011_bfr_after (
		.din(new_net_2010),
		.dout(new_net_2011)
	);

	bfr new_net_2012_bfr_after (
		.din(new_net_2011),
		.dout(new_net_2012)
	);

	bfr new_net_475_bfr_after (
		.din(new_net_2012),
		.dout(new_net_475)
	);

	bfr new_net_2013_bfr_after (
		.din(_161_),
		.dout(new_net_2013)
	);

	bfr new_net_2014_bfr_after (
		.din(new_net_2013),
		.dout(new_net_2014)
	);

	bfr new_net_2015_bfr_after (
		.din(new_net_2014),
		.dout(new_net_2015)
	);

	bfr new_net_2016_bfr_after (
		.din(new_net_2015),
		.dout(new_net_2016)
	);

	bfr new_net_2017_bfr_after (
		.din(new_net_2016),
		.dout(new_net_2017)
	);

	bfr new_net_488_bfr_after (
		.din(new_net_2017),
		.dout(new_net_488)
	);

	bfr new_net_2018_bfr_after (
		.din(_178_),
		.dout(new_net_2018)
	);

	bfr new_net_2019_bfr_after (
		.din(new_net_2018),
		.dout(new_net_2019)
	);

	bfr new_net_2020_bfr_after (
		.din(new_net_2019),
		.dout(new_net_2020)
	);

	bfr new_net_2021_bfr_after (
		.din(new_net_2020),
		.dout(new_net_2021)
	);

	bfr new_net_496_bfr_after (
		.din(new_net_2021),
		.dout(new_net_496)
	);

	bfr new_net_509_bfr_after (
		.din(_207_),
		.dout(new_net_509)
	);

	bfr new_net_517_bfr_after (
		.din(_270_),
		.dout(new_net_517)
	);

	bfr new_net_2022_bfr_after (
		.din(_012_),
		.dout(new_net_2022)
	);

	bfr new_net_2023_bfr_after (
		.din(new_net_2022),
		.dout(new_net_2023)
	);

	bfr new_net_2024_bfr_after (
		.din(new_net_2023),
		.dout(new_net_2024)
	);

	bfr new_net_454_bfr_after (
		.din(new_net_2024),
		.dout(new_net_454)
	);

	bfr new_net_2025_bfr_after (
		.din(_081_),
		.dout(new_net_2025)
	);

	bfr new_net_2026_bfr_after (
		.din(new_net_2025),
		.dout(new_net_2026)
	);

	bfr new_net_2027_bfr_after (
		.din(new_net_2026),
		.dout(new_net_2027)
	);

	bfr new_net_2028_bfr_after (
		.din(new_net_2027),
		.dout(new_net_2028)
	);

	bfr new_net_2029_bfr_after (
		.din(new_net_2028),
		.dout(new_net_2029)
	);

	bfr new_net_2030_bfr_after (
		.din(new_net_2029),
		.dout(new_net_2030)
	);

	bfr new_net_467_bfr_after (
		.din(new_net_2030),
		.dout(new_net_467)
	);

	bfr new_net_2031_bfr_after (
		.din(_119_),
		.dout(new_net_2031)
	);

	bfr new_net_2032_bfr_after (
		.din(new_net_2031),
		.dout(new_net_2032)
	);

	bfr new_net_2033_bfr_after (
		.din(new_net_2032),
		.dout(new_net_2033)
	);

	bfr new_net_2034_bfr_after (
		.din(new_net_2033),
		.dout(new_net_2034)
	);

	bfr new_net_2035_bfr_after (
		.din(new_net_2034),
		.dout(new_net_2035)
	);

	bfr new_net_471_bfr_after (
		.din(new_net_2035),
		.dout(new_net_471)
	);

	bfr new_net_2036_bfr_after (
		.din(_165_),
		.dout(new_net_2036)
	);

	bfr new_net_2037_bfr_after (
		.din(new_net_2036),
		.dout(new_net_2037)
	);

	bfr new_net_2038_bfr_after (
		.din(new_net_2037),
		.dout(new_net_2038)
	);

	bfr new_net_2039_bfr_after (
		.din(new_net_2038),
		.dout(new_net_2039)
	);

	bfr new_net_2040_bfr_after (
		.din(new_net_2039),
		.dout(new_net_2040)
	);

	bfr new_net_2041_bfr_after (
		.din(new_net_2040),
		.dout(new_net_2041)
	);

	bfr new_net_492_bfr_after (
		.din(new_net_2041),
		.dout(new_net_492)
	);

	bfr new_net_513_bfr_after (
		.din(_212_),
		.dout(new_net_513)
	);

	bfr new_net_2042_bfr_after (
		.din(new_net_546),
		.dout(new_net_2042)
	);

	bfr new_net_2043_bfr_after (
		.din(new_net_2042),
		.dout(new_net_2043)
	);

	bfr new_net_2044_bfr_after (
		.din(new_net_2043),
		.dout(new_net_2044)
	);

	bfr new_net_2045_bfr_after (
		.din(new_net_2044),
		.dout(new_net_2045)
	);

	bfr new_net_2046_bfr_after (
		.din(new_net_2045),
		.dout(new_net_2046)
	);

	bfr new_net_2047_bfr_after (
		.din(new_net_2046),
		.dout(new_net_2047)
	);

	bfr new_net_2048_bfr_after (
		.din(new_net_2047),
		.dout(new_net_2048)
	);

	bfr new_net_2049_bfr_after (
		.din(new_net_2048),
		.dout(new_net_2049)
	);

	bfr new_net_2050_bfr_after (
		.din(new_net_2049),
		.dout(new_net_2050)
	);

	bfr new_net_2051_bfr_after (
		.din(new_net_2050),
		.dout(new_net_2051)
	);

	bfr new_net_2052_bfr_after (
		.din(new_net_2051),
		.dout(new_net_2052)
	);

	bfr new_net_2053_bfr_after (
		.din(new_net_2052),
		.dout(new_net_2053)
	);

	bfr new_net_2054_bfr_after (
		.din(new_net_2053),
		.dout(new_net_2054)
	);

	bfr new_net_2055_bfr_after (
		.din(new_net_2054),
		.dout(new_net_2055)
	);

	bfr new_net_2056_bfr_after (
		.din(new_net_2055),
		.dout(new_net_2056)
	);

	bfr new_net_2057_bfr_after (
		.din(new_net_2056),
		.dout(new_net_2057)
	);

	bfr new_net_2058_bfr_after (
		.din(new_net_2057),
		.dout(new_net_2058)
	);

	bfr new_net_2059_bfr_after (
		.din(new_net_2058),
		.dout(new_net_2059)
	);

	bfr new_net_2060_bfr_after (
		.din(new_net_2059),
		.dout(new_net_2060)
	);

	bfr new_net_2061_bfr_after (
		.din(new_net_2060),
		.dout(new_net_2061)
	);

	bfr new_net_2062_bfr_after (
		.din(new_net_2061),
		.dout(new_net_2062)
	);

	bfr new_net_2063_bfr_after (
		.din(new_net_2062),
		.dout(new_net_2063)
	);

	bfr new_net_2064_bfr_after (
		.din(new_net_2063),
		.dout(new_net_2064)
	);

	bfr new_net_2065_bfr_after (
		.din(new_net_2064),
		.dout(new_net_2065)
	);

	bfr new_net_2066_bfr_after (
		.din(new_net_2065),
		.dout(new_net_2066)
	);

	bfr new_net_2067_bfr_after (
		.din(new_net_2066),
		.dout(new_net_2067)
	);

	bfr new_net_2068_bfr_after (
		.din(new_net_2067),
		.dout(new_net_2068)
	);

	bfr new_net_2069_bfr_after (
		.din(new_net_2068),
		.dout(new_net_2069)
	);

	bfr new_net_2070_bfr_after (
		.din(new_net_2069),
		.dout(new_net_2070)
	);

	bfr new_net_2071_bfr_after (
		.din(new_net_2070),
		.dout(new_net_2071)
	);

	bfr new_net_2072_bfr_after (
		.din(new_net_2071),
		.dout(new_net_2072)
	);

	bfr new_net_2073_bfr_after (
		.din(new_net_2072),
		.dout(new_net_2073)
	);

	bfr new_net_2074_bfr_after (
		.din(new_net_2073),
		.dout(new_net_2074)
	);

	bfr new_net_2075_bfr_after (
		.din(new_net_2074),
		.dout(new_net_2075)
	);

	bfr new_net_2076_bfr_after (
		.din(new_net_2075),
		.dout(new_net_2076)
	);

	bfr new_net_2077_bfr_after (
		.din(new_net_2076),
		.dout(new_net_2077)
	);

	bfr N388_bfr_after (
		.din(new_net_2077),
		.dout(N388)
	);

endmodule