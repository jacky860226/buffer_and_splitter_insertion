module c499(N97,N113,N73,N134,N57,N77,N17,N49,N93,N1,N131,N25,N109,N45,N132,N135,N61,N85,N117,N21,N33,N101,N81,N105,N41,N5,N130,N133,N89,N125,N53,N69,N29,N121,N9,N13,N137,N37,N136,N129,N65);
    wire _075_;
    wire new_Jinkela_wire_312;
    wire new_Jinkela_wire_467;
    wire new_Jinkela_wire_709;
    wire new_net_711;
    wire new_Jinkela_wire_1706;
    wire new_Jinkela_wire_690;
    wire new_Jinkela_wire_229;
    wire new_Jinkela_wire_845;
    wire _054_;
    wire new_Jinkela_wire_1464;
    wire new_Jinkela_wire_1227;
    wire new_net_697;
    wire new_Jinkela_wire_1007;
    wire new_Jinkela_wire_829;
    wire new_Jinkela_wire_629;
    wire _028_;
    wire new_Jinkela_wire_1677;
    wire new_Jinkela_wire_284;
    wire new_Jinkela_wire_1112;
    wire new_Jinkela_wire_948;
    wire _240_;
    wire new_Jinkela_wire_1122;
    wire new_Jinkela_wire_1352;
    wire _325_;
    wire new_Jinkela_wire_653;
    wire new_Jinkela_wire_273;
    wire new_Jinkela_wire_1103;
    wire new_Jinkela_wire_498;
    wire new_Jinkela_wire_1114;
    wire _337_;
    wire new_Jinkela_wire_1279;
    wire _018_;
    wire new_Jinkela_wire_1672;
    wire _174_;
    wire new_Jinkela_wire_176;
    wire _256_;
    wire _020_;
    wire new_Jinkela_wire_1014;
    wire new_Jinkela_wire_562;
    wire new_Jinkela_wire_639;
    wire new_Jinkela_wire_422;
    wire new_Jinkela_wire_432;
    wire new_Jinkela_wire_860;
    wire new_Jinkela_wire_1634;
    wire _350_;
    wire new_Jinkela_wire_678;
    wire new_Jinkela_wire_666;
    wire new_Jinkela_wire_1600;
    wire _262_;
    wire _298_;
    wire new_Jinkela_wire_324;
    wire _161_;
    wire new_Jinkela_wire_476;
    wire new_Jinkela_wire_864;
    wire _056_;
    wire new_Jinkela_wire_878;
    wire new_Jinkela_wire_1480;
    wire new_Jinkela_wire_1460;
    wire new_Jinkela_wire_1115;
    wire new_Jinkela_wire_1088;
    wire _115_;
    wire new_Jinkela_wire_395;
    wire new_Jinkela_wire_1544;
    wire _166_;
    wire new_Jinkela_wire_1427;
    wire new_Jinkela_wire_294;
    wire new_Jinkela_wire_899;
    wire new_Jinkela_wire_1218;
    wire new_Jinkela_wire_1337;
    wire new_Jinkela_wire_1246;
    wire _305_;
    wire new_Jinkela_wire_462;
    wire new_Jinkela_wire_785;
    wire new_Jinkela_wire_1639;
    wire new_Jinkela_wire_1381;
    wire new_Jinkela_wire_1553;
    wire new_Jinkela_wire_1371;
    wire new_Jinkela_wire_410;
    wire new_Jinkela_wire_1186;
    wire new_Jinkela_wire_652;
    wire new_Jinkela_wire_265;
    wire new_Jinkela_wire_1378;
    wire _040_;
    wire new_Jinkela_wire_170;
    wire new_Jinkela_wire_1468;
    wire new_Jinkela_wire_777;
    wire new_Jinkela_wire_1546;
    wire _004_;
    wire new_Jinkela_wire_798;
    wire new_Jinkela_wire_1031;
    wire _326_;
    wire new_Jinkela_wire_789;
    wire _264_;
    wire new_Jinkela_wire_1450;
    wire new_Jinkela_wire_227;
    wire new_Jinkela_wire_1043;
    wire new_Jinkela_wire_1162;
    wire new_Jinkela_wire_402;
    wire new_Jinkela_wire_287;
    wire new_Jinkela_wire_258;
    wire new_Jinkela_wire_20;
    wire new_Jinkela_wire_922;
    wire new_Jinkela_wire_212;
    wire new_Jinkela_wire_851;
    wire new_Jinkela_wire_1426;
    wire new_Jinkela_wire_48;
    wire new_Jinkela_wire_916;
    wire _250_;
    wire new_Jinkela_wire_974;
    wire new_Jinkela_wire_1080;
    wire _200_;
    wire new_Jinkela_wire_580;
    wire _108_;
    wire new_Jinkela_wire_1008;
    wire new_Jinkela_wire_438;
    wire new_Jinkela_wire_102;
    wire new_Jinkela_wire_26;
    wire new_Jinkela_wire_730;
    wire new_Jinkela_wire_1414;
    wire _210_;
    wire new_Jinkela_wire_488;
    wire new_Jinkela_wire_427;
    wire new_Jinkela_wire_1070;
    wire _137_;
    wire _345_;
    wire new_Jinkela_wire_906;
    wire new_Jinkela_wire_1135;
    wire new_Jinkela_wire_145;
    wire new_Jinkela_wire_1309;
    wire _331_;
    wire new_Jinkela_wire_753;
    wire new_Jinkela_wire_1271;
    wire new_Jinkela_wire_695;
    wire new_Jinkela_wire_523;
    wire new_Jinkela_wire_497;
    wire new_Jinkela_wire_1182;
    wire _320_;
    wire new_Jinkela_wire_1647;
    wire _280_;
    wire new_Jinkela_wire_1287;
    wire new_Jinkela_wire_1219;
    wire new_Jinkela_wire_748;
    wire new_Jinkela_wire_286;
    wire new_Jinkela_wire_778;
    wire new_Jinkela_wire_177;
    wire new_Jinkela_wire_314;
    wire new_Jinkela_wire_1291;
    wire new_Jinkela_wire_1083;
    wire new_Jinkela_wire_591;
    wire _273_;
    wire new_Jinkela_wire_53;
    wire _025_;
    wire new_Jinkela_wire_1506;
    wire _089_;
    wire new_Jinkela_wire_1689;
    wire _031_;
    wire new_Jinkela_wire_1651;
    wire new_Jinkela_wire_1377;
    wire new_Jinkela_wire_542;
    wire _184_;
    wire _236_;
    wire new_Jinkela_wire_866;
    wire new_Jinkela_wire_1534;
    wire new_Jinkela_wire_644;
    wire new_net_691;
    wire new_Jinkela_wire_1106;
    wire new_Jinkela_wire_371;
    wire new_Jinkela_wire_1382;
    wire new_Jinkela_wire_988;
    wire _204_;
    wire new_Jinkela_wire_172;
    wire new_Jinkela_wire_1342;
    wire new_Jinkela_wire_1111;
    wire new_Jinkela_wire_1074;
    wire new_Jinkela_wire_704;
    wire _042_;
    wire new_Jinkela_wire_1684;
    wire new_Jinkela_wire_801;
    wire new_Jinkela_wire_1329;
    wire new_Jinkela_wire_308;
    wire new_net_703;
    wire _100_;
    wire new_Jinkela_wire_1668;
    wire new_Jinkela_wire_931;
    wire new_Jinkela_wire_1564;
    wire _271_;
    wire new_Jinkela_wire_1095;
    wire new_Jinkela_wire_821;
    wire _101_;
    wire new_Jinkela_wire_1389;
    wire _046_;
    wire _283_;
    wire new_Jinkela_wire_862;
    wire new_Jinkela_wire_321;
    wire new_Jinkela_wire_376;
    wire new_Jinkela_wire_1277;
    wire new_Jinkela_wire_1057;
    wire new_Jinkela_wire_22;
    wire new_Jinkela_wire_854;
    wire new_Jinkela_wire_1139;
    wire new_Jinkela_wire_1631;
    wire new_Jinkela_wire_1078;
    wire new_Jinkela_wire_555;
    wire new_Jinkela_wire_157;
    wire _338_;
    wire new_Jinkela_wire_103;
    wire new_Jinkela_wire_761;
    wire new_Jinkela_wire_952;
    wire _328_;
    wire new_Jinkela_wire_1286;
    wire _022_;
    wire new_net_699;
    wire new_Jinkela_wire_1061;
    wire new_Jinkela_wire_654;
    wire new_Jinkela_wire_871;
    wire new_Jinkela_wire_769;
    wire _206_;
    wire new_Jinkela_wire_962;
    wire new_Jinkela_wire_786;
    wire new_Jinkela_wire_722;
    wire new_Jinkela_wire_260;
    wire new_Jinkela_wire_707;
    wire new_Jinkela_wire_1366;
    wire _217_;
    wire new_Jinkela_wire_784;
    wire new_Jinkela_wire_49;
    wire new_Jinkela_wire_246;
    wire new_Jinkela_wire_514;
    wire new_Jinkela_wire_734;
    wire new_Jinkela_wire_243;
    wire new_Jinkela_wire_1496;
    wire new_Jinkela_wire_736;
    wire new_Jinkela_wire_1133;
    wire new_Jinkela_wire_1116;
    wire new_Jinkela_wire_1081;
    wire new_Jinkela_wire_839;
    wire new_Jinkela_wire_224;
    wire new_Jinkela_wire_913;
    wire new_Jinkela_wire_1517;
    wire new_Jinkela_wire_708;
    wire new_Jinkela_wire_1124;
    wire new_Jinkela_wire_429;
    wire new_Jinkela_wire_558;
    wire new_Jinkela_wire_368;
    wire new_Jinkela_wire_990;
    wire _279_;
    wire new_Jinkela_wire_670;
    wire _119_;
    wire new_Jinkela_wire_1601;
    wire new_Jinkela_wire_466;
    wire new_Jinkela_wire_1033;
    wire new_Jinkela_wire_524;
    wire new_Jinkela_wire_585;
    wire new_Jinkela_wire_1569;
    wire new_Jinkela_wire_685;
    wire new_Jinkela_wire_384;
    wire new_Jinkela_wire_1385;
    wire new_Jinkela_wire_1265;
    wire new_Jinkela_wire_1536;
    wire new_Jinkela_wire_1599;
    wire _277_;
    wire _238_;
    wire new_Jinkela_wire_1422;
    wire new_Jinkela_wire_1692;
    wire new_Jinkela_wire_393;
    wire new_Jinkela_wire_927;
    wire new_Jinkela_wire_1364;
    wire _339_;
    wire new_Jinkela_wire_511;
    wire new_Jinkela_wire_627;
    wire new_Jinkela_wire_1221;
    wire new_Jinkela_wire_793;
    wire new_Jinkela_wire_1361;
    wire new_Jinkela_wire_664;
    wire new_Jinkela_wire_367;
    wire new_Jinkela_wire_835;
    wire _124_;
    wire new_Jinkela_wire_1454;
    wire new_Jinkela_wire_1363;
    wire new_Jinkela_wire_842;
    wire new_Jinkela_wire_1550;
    wire new_Jinkela_wire_1524;
    wire new_Jinkela_wire_226;
    wire new_Jinkela_wire_248;
    wire new_Jinkela_wire_655;
    wire new_Jinkela_wire_1000;
    wire new_Jinkela_wire_1025;
    wire new_Jinkela_wire_1671;
    wire new_Jinkela_wire_1065;
    wire _144_;
    wire new_Jinkela_wire_253;
    wire new_Jinkela_wire_1551;
    wire new_Jinkela_wire_756;
    wire new_Jinkela_wire_451;
    wire new_Jinkela_wire_885;
    wire _029_;
    wire new_Jinkela_wire_1359;
    wire new_Jinkela_wire_323;
    wire new_net_701;
    wire new_Jinkela_wire_135;
    wire new_Jinkela_wire_72;
    wire _288_;
    wire _340_;
    wire new_Jinkela_wire_1260;
    wire new_Jinkela_wire_755;
    wire new_Jinkela_wire_1311;
    wire new_Jinkela_wire_943;
    wire new_Jinkela_wire_1147;
    wire new_Jinkela_wire_1243;
    wire _087_;
    wire new_Jinkela_wire_547;
    wire new_Jinkela_wire_1404;
    wire _287_;
    wire new_Jinkela_wire_1241;
    wire new_Jinkela_wire_1392;
    wire new_Jinkela_wire_592;
    wire new_Jinkela_wire_1494;
    wire new_Jinkela_wire_993;
    wire new_Jinkela_wire_571;
    wire new_Jinkela_wire_40;
    wire new_Jinkela_wire_1251;
    wire new_Jinkela_wire_297;
    wire new_Jinkela_wire_1263;
    wire new_Jinkela_wire_968;
    wire new_Jinkela_wire_1053;
    wire new_Jinkela_wire_945;
    wire new_Jinkela_wire_1444;
    wire new_Jinkela_wire_77;
    wire _284_;
    wire new_Jinkela_wire_446;
    wire new_Jinkela_wire_119;
    wire _005_;
    wire new_Jinkela_wire_74;
    wire new_Jinkela_wire_183;
    wire _164_;
    wire new_Jinkela_wire_904;
    wire new_Jinkela_wire_1159;
    wire new_Jinkela_wire_1570;
    wire new_Jinkela_wire_551;
    wire new_Jinkela_wire_425;
    wire _012_;
    wire new_Jinkela_wire_32;
    wire new_Jinkela_wire_282;
    wire new_Jinkela_wire_548;
    wire new_Jinkela_wire_1375;
    wire _323_;
    wire new_Jinkela_wire_716;
    wire new_Jinkela_wire_1092;
    wire new_Jinkela_wire_0;
    wire _334_;
    wire new_Jinkela_wire_1022;
    wire new_Jinkela_wire_574;
    wire new_Jinkela_wire_8;
    wire new_Jinkela_wire_1071;
    wire new_Jinkela_wire_1435;
    wire new_Jinkela_wire_628;
    wire new_Jinkela_wire_1062;
    wire new_Jinkela_wire_667;
    wire new_Jinkela_wire_219;
    wire new_Jinkela_wire_521;
    wire new_Jinkela_wire_30;
    wire new_Jinkela_wire_517;
    wire new_Jinkela_wire_963;
    wire new_Jinkela_wire_350;
    wire new_Jinkela_wire_1049;
    wire new_Jinkela_wire_1195;
    wire new_Jinkela_wire_987;
    wire new_Jinkela_wire_471;
    wire new_Jinkela_wire_1627;
    wire new_Jinkela_wire_478;
    wire new_Jinkela_wire_951;
    wire new_Jinkela_wire_518;
    wire new_Jinkela_wire_805;
    wire _246_;
    wire new_Jinkela_wire_276;
    wire new_Jinkela_wire_1183;
    wire _041_;
    wire new_Jinkela_wire_740;
    wire new_Jinkela_wire_1121;
    wire new_Jinkela_wire_687;
    wire new_Jinkela_wire_1515;
    wire new_Jinkela_wire_1581;
    wire new_Jinkela_wire_1533;
    wire new_Jinkela_wire_1175;
    wire new_Jinkela_wire_924;
    wire new_Jinkela_wire_148;
    wire new_Jinkela_wire_831;
    wire _234_;
    wire new_Jinkela_wire_453;
    wire new_Jinkela_wire_823;
    wire new_Jinkela_wire_1586;
    wire _149_;
    wire new_Jinkela_wire_1530;
    wire new_Jinkela_wire_621;
    wire new_Jinkela_wire_1673;
    wire _021_;
    wire new_Jinkela_wire_1261;
    wire new_Jinkela_wire_1622;
    wire _195_;
    wire new_Jinkela_wire_206;
    wire new_Jinkela_wire_721;
    wire new_Jinkela_wire_163;
    wire _084_;
    wire new_net_693;
    wire new_Jinkela_wire_554;
    wire _332_;
    wire new_Jinkela_wire_433;
    wire new_Jinkela_wire_357;
    wire _008_;
    wire new_Jinkela_wire_252;
    wire new_Jinkela_wire_541;
    wire new_Jinkela_wire_1050;
    wire new_Jinkela_wire_1556;
    wire new_Jinkela_wire_283;
    wire new_Jinkela_wire_1082;
    wire new_Jinkela_wire_411;
    wire new_Jinkela_wire_1130;
    wire new_Jinkela_wire_15;
    wire new_Jinkela_wire_334;
    wire new_Jinkela_wire_280;
    wire new_Jinkela_wire_1678;
    wire new_Jinkela_wire_1502;
    wire _306_;
    wire new_Jinkela_wire_979;
    wire new_Jinkela_wire_475;
    wire new_Jinkela_wire_980;
    wire new_Jinkela_wire_1305;
    wire new_Jinkela_wire_116;
    wire new_Jinkela_wire_1003;
    wire new_Jinkela_wire_1641;
    wire _270_;
    wire new_Jinkela_wire_991;
    wire new_Jinkela_wire_443;
    wire _002_;
    wire new_Jinkela_wire_1225;
    wire new_Jinkela_wire_1244;
    wire new_Jinkela_wire_111;
    wire new_Jinkela_wire_1620;
    wire new_Jinkela_wire_776;
    wire new_Jinkela_wire_837;
    wire new_Jinkela_wire_494;
    wire new_Jinkela_wire_747;
    wire _230_;
    wire new_Jinkela_wire_174;
    wire new_Jinkela_wire_1577;
    wire new_Jinkela_wire_549;
    wire new_Jinkela_wire_474;
    wire new_Jinkela_wire_1344;
    wire new_Jinkela_wire_220;
    wire new_Jinkela_wire_787;
    wire new_Jinkela_wire_184;
    wire new_Jinkela_wire_81;
    wire _116_;
    wire new_Jinkela_wire_1500;
    wire new_Jinkela_wire_1197;
    wire new_Jinkela_wire_1486;
    wire new_Jinkela_wire_84;
    wire new_Jinkela_wire_573;
    wire new_Jinkela_wire_1273;
    wire new_Jinkela_wire_674;
    wire new_Jinkela_wire_1452;
    wire new_Jinkela_wire_503;
    wire _243_;
    wire new_Jinkela_wire_298;
    wire new_Jinkela_wire_117;
    wire new_Jinkela_wire_266;
    wire _356_;
    wire _102_;
    wire new_Jinkela_wire_659;
    wire _027_;
    wire new_Jinkela_wire_397;
    wire new_Jinkela_wire_1212;
    wire new_Jinkela_wire_836;
    wire new_Jinkela_wire_1583;
    wire _052_;
    wire new_Jinkela_wire_359;
    wire new_Jinkela_wire_442;
    wire new_Jinkela_wire_441;
    wire new_Jinkela_wire_290;
    wire _093_;
    wire new_Jinkela_wire_61;
    wire _055_;
    wire new_Jinkela_wire_242;
    wire _114_;
    wire new_Jinkela_wire_168;
    wire new_Jinkela_wire_879;
    wire new_Jinkela_wire_1403;
    wire _047_;
    wire _263_;
    wire new_Jinkela_wire_673;
    wire new_Jinkela_wire_315;
    wire new_Jinkela_wire_535;
    wire new_Jinkela_wire_955;
    wire new_Jinkela_wire_1438;
    wire new_Jinkela_wire_1370;
    wire _096_;
    wire new_Jinkela_wire_636;
    wire new_Jinkela_wire_1242;
    wire new_Jinkela_wire_256;
    wire new_Jinkela_wire_1535;
    wire new_Jinkela_wire_969;
    wire new_Jinkela_wire_1499;
    wire _252_;
    wire new_Jinkela_wire_338;
    wire _138_;
    wire new_Jinkela_wire_754;
    wire new_Jinkela_wire_167;
    wire _076_;
    wire new_Jinkela_wire_731;
    wire _312_;
    wire new_Jinkela_wire_665;
    wire new_Jinkela_wire_1128;
    wire _120_;
    wire new_Jinkela_wire_1701;
    wire new_Jinkela_wire_1594;
    wire new_Jinkela_wire_1621;
    wire _083_;
    wire new_Jinkela_wire_285;
    wire _038_;
    wire new_Jinkela_wire_13;
    wire new_Jinkela_wire_1430;
    wire new_Jinkela_wire_464;
    wire new_Jinkela_wire_1134;
    wire new_Jinkela_wire_73;
    wire new_Jinkela_wire_589;
    wire new_Jinkela_wire_470;
    wire new_Jinkela_wire_956;
    wire new_Jinkela_wire_1380;
    wire new_Jinkela_wire_643;
    wire new_Jinkela_wire_86;
    wire _024_;
    wire new_Jinkela_wire_701;
    wire new_Jinkela_wire_938;
    wire new_Jinkela_wire_108;
    wire new_Jinkela_wire_440;
    wire new_Jinkela_wire_1656;
    wire _214_;
    wire new_Jinkela_wire_1394;
    wire _173_;
    wire _346_;
    wire _167_;
    wire new_Jinkela_wire_1350;
    wire new_Jinkela_wire_43;
    wire new_Jinkela_wire_1193;
    wire new_Jinkela_wire_351;
    wire new_Jinkela_wire_647;
    wire new_Jinkela_wire_1058;
    wire new_Jinkela_wire_1048;
    wire new_Jinkela_wire_985;
    wire new_Jinkela_wire_934;
    wire new_Jinkela_wire_819;
    wire _219_;
    wire new_Jinkela_wire_391;
    wire new_Jinkela_wire_133;
    wire new_Jinkela_wire_1052;
    wire _033_;
    wire new_Jinkela_wire_407;
    wire new_Jinkela_wire_295;
    wire new_Jinkela_wire_729;
    wire new_Jinkela_wire_1343;
    wire new_Jinkela_wire_71;
    wire new_Jinkela_wire_406;
    wire new_Jinkela_wire_604;
    wire new_Jinkela_wire_949;
    wire _071_;
    wire new_Jinkela_wire_630;
    wire new_Jinkela_wire_1275;
    wire _354_;
    wire new_Jinkela_wire_1315;
    wire _245_;
    wire new_Jinkela_wire_37;
    wire new_Jinkela_wire_1449;
    wire new_Jinkela_wire_1603;
    wire new_Jinkela_wire_1376;
    wire _182_;
    wire new_Jinkela_wire_329;
    wire new_Jinkela_wire_486;
    wire _158_;
    wire new_Jinkela_wire_992;
    wire new_Jinkela_wire_1521;
    wire new_Jinkela_wire_1072;
    wire _228_;
    wire new_Jinkela_wire_143;
    wire new_Jinkela_wire_1210;
    wire new_Jinkela_wire_883;
    wire new_Jinkela_wire_7;
    wire new_Jinkela_wire_561;
    wire new_Jinkela_wire_1300;
    wire new_Jinkela_wire_677;
    wire new_Jinkela_wire_1436;
    wire _260_;
    wire new_Jinkela_wire_867;
    wire new_Jinkela_wire_1046;
    wire new_Jinkela_wire_1593;
    wire new_Jinkela_wire_1228;
    wire new_Jinkela_wire_1021;
    wire new_Jinkela_wire_1304;
    wire _133_;
    wire new_Jinkela_wire_1519;
    wire new_Jinkela_wire_512;
    wire new_Jinkela_wire_536;
    wire new_Jinkela_wire_1395;
    wire new_Jinkela_wire_1670;
    wire new_Jinkela_wire_700;
    wire new_Jinkela_wire_1044;
    wire new_Jinkela_wire_876;
    wire new_Jinkela_wire_495;
    wire new_Jinkela_wire_21;
    wire new_Jinkela_wire_1507;
    wire new_Jinkela_wire_502;
    wire new_Jinkela_wire_483;
    wire new_Jinkela_wire_702;
    wire new_Jinkela_wire_1643;
    wire new_Jinkela_wire_1419;
    wire new_Jinkela_wire_1475;
    wire new_Jinkela_wire_1029;
    wire new_Jinkela_wire_1332;
    wire new_Jinkela_wire_972;
    wire new_Jinkela_wire_1245;
    wire new_Jinkela_wire_928;
    wire new_Jinkela_wire_905;
    wire new_Jinkela_wire_765;
    wire new_Jinkela_wire_935;
    wire new_Jinkela_wire_313;
    wire new_Jinkela_wire_1509;
    wire new_Jinkela_wire_901;
    wire new_Jinkela_wire_231;
    wire new_Jinkela_wire_301;
    wire new_Jinkela_wire_1443;
    wire new_Jinkela_wire_1030;
    wire _193_;
    wire new_Jinkela_wire_1153;
    wire new_Jinkela_wire_645;
    wire new_Jinkela_wire_1520;
    wire new_Jinkela_wire_875;
    wire new_Jinkela_wire_1169;
    wire new_Jinkela_wire_59;
    wire new_Jinkela_wire_919;
    wire new_Jinkela_wire_354;
    wire new_Jinkela_wire_1471;
    wire new_Jinkela_wire_1384;
    wire new_Jinkela_wire_479;
    wire new_Jinkela_wire_539;
    wire new_Jinkela_wire_444;
    wire new_Jinkela_wire_1495;
    wire new_Jinkela_wire_1223;
    wire new_Jinkela_wire_352;
    wire new_Jinkela_wire_1649;
    wire new_Jinkela_wire_196;
    wire new_Jinkela_wire_527;
    wire new_Jinkela_wire_1158;
    wire new_Jinkela_wire_584;
    wire _289_;
    wire new_Jinkela_wire_510;
    wire new_Jinkela_wire_468;
    wire new_Jinkela_wire_1146;
    wire new_Jinkela_wire_398;
    wire new_Jinkela_wire_180;
    wire new_Jinkela_wire_613;
    wire new_Jinkela_wire_1293;
    wire new_Jinkela_wire_1064;
    wire new_Jinkela_wire_848;
    wire new_Jinkela_wire_54;
    wire _297_;
    wire new_Jinkela_wire_746;
    wire new_Jinkela_wire_619;
    wire new_Jinkela_wire_198;
    wire new_Jinkela_wire_1440;
    wire new_Jinkela_wire_162;
    wire new_Jinkela_wire_1016;
    wire new_Jinkela_wire_238;
    wire new_Jinkela_wire_487;
    wire _132_;
    wire new_Jinkela_wire_118;
    wire new_Jinkela_wire_1549;
    wire _177_;
    wire new_Jinkela_wire_1298;
    wire new_Jinkela_wire_1433;
    wire new_Jinkela_wire_83;
    wire new_Jinkela_wire_852;
    wire new_Jinkela_wire_45;
    wire new_Jinkela_wire_681;
    wire new_Jinkela_wire_953;
    wire _143_;
    wire new_Jinkela_wire_642;
    wire _053_;
    wire new_net_687;
    wire _275_;
    wire new_Jinkela_wire_1015;
    wire new_Jinkela_wire_1662;
    wire new_Jinkela_wire_1666;
    wire new_Jinkela_wire_767;
    wire new_Jinkela_wire_1568;
    wire new_Jinkela_wire_491;
    wire _282_;
    wire new_Jinkela_wire_1700;
    wire new_Jinkela_wire_1168;
    wire new_Jinkela_wire_1368;
    wire new_Jinkela_wire_1574;
    wire new_Jinkela_wire_902;
    wire new_Jinkela_wire_1131;
    wire new_Jinkela_wire_782;
    wire new_Jinkela_wire_1207;
    wire new_Jinkela_wire_1708;
    wire new_Jinkela_wire_465;
    wire new_Jinkela_wire_1323;
    wire new_Jinkela_wire_1037;
    wire new_Jinkela_wire_431;
    wire new_Jinkela_wire_872;
    wire _223_;
    wire _254_;
    wire _081_;
    wire _126_;
    wire new_Jinkela_wire_994;
    wire new_Jinkela_wire_1630;
    wire new_Jinkela_wire_1327;
    wire new_Jinkela_wire_1388;
    wire new_Jinkela_wire_1313;
    wire new_Jinkela_wire_1256;
    wire _293_;
    wire new_Jinkela_wire_1063;
    wire new_Jinkela_wire_182;
    wire new_Jinkela_wire_213;
    wire new_Jinkela_wire_1614;
    wire new_Jinkela_wire_720;
    wire new_Jinkela_wire_847;
    wire new_Jinkela_wire_1412;
    wire new_Jinkela_wire_890;
    wire new_Jinkela_wire_1379;
    wire new_Jinkela_wire_469;
    wire new_Jinkela_wire_1307;
    wire new_Jinkela_wire_565;
    wire new_Jinkela_wire_1595;
    wire new_Jinkela_wire_1628;
    wire _187_;
    wire new_Jinkela_wire_543;
    wire _127_;
    wire new_Jinkela_wire_41;
    wire new_Jinkela_wire_1602;
    wire _308_;
    wire new_Jinkela_wire_1458;
    wire new_Jinkela_wire_154;
    wire _036_;
    wire new_Jinkela_wire_1316;
    wire new_Jinkela_wire_239;
    wire new_Jinkela_wire_1638;
    wire new_Jinkela_wire_807;
    wire new_Jinkela_wire_662;
    wire new_Jinkela_wire_159;
    wire new_Jinkela_wire_82;
    wire new_Jinkela_wire_1266;
    wire _037_;
    wire new_Jinkela_wire_293;
    wire new_Jinkela_wire_1400;
    wire new_Jinkela_wire_1039;
    wire _003_;
    wire new_Jinkela_wire_937;
    wire new_Jinkela_wire_1554;
    wire new_Jinkela_wire_56;
    wire _181_;
    wire new_Jinkela_wire_546;
    wire new_Jinkela_wire_57;
    wire _048_;
    wire new_net_695;
    wire new_Jinkela_wire_932;
    wire new_Jinkela_wire_809;
    wire new_Jinkela_wire_288;
    wire new_Jinkela_wire_1170;
    wire new_Jinkela_wire_689;
    wire _202_;
    wire new_Jinkela_wire_79;
    wire _072_;
    wire new_Jinkela_wire_1118;
    wire new_Jinkela_wire_1239;
    wire new_Jinkela_wire_973;
    wire new_Jinkela_wire_343;
    wire _207_;
    wire new_Jinkela_wire_1119;
    wire new_Jinkela_wire_772;
    wire new_Jinkela_wire_214;
    wire new_Jinkela_wire_385;
    wire new_Jinkela_wire_186;
    wire _110_;
    wire new_Jinkela_wire_1633;
    wire new_Jinkela_wire_1222;
    wire _249_;
    wire new_Jinkela_wire_660;
    wire new_Jinkela_wire_1445;
    wire new_Jinkela_wire_5;
    wire new_Jinkela_wire_1616;
    wire new_Jinkela_wire_207;
    wire new_Jinkela_wire_67;
    wire _180_;
    wire new_Jinkela_wire_1085;
    wire new_Jinkela_wire_94;
    wire new_Jinkela_wire_680;
    wire new_Jinkela_wire_684;
    wire new_Jinkela_wire_232;
    wire _319_;
    wire new_Jinkela_wire_344;
    wire new_Jinkela_wire_850;
    wire new_Jinkela_wire_1528;
    wire new_Jinkela_wire_193;
    wire new_Jinkela_wire_873;
    wire new_Jinkela_wire_44;
    wire new_Jinkela_wire_737;
    wire new_Jinkela_wire_921;
    wire new_Jinkela_wire_1374;
    wire new_Jinkela_wire_1653;
    wire new_Jinkela_wire_958;
    wire new_net_707;
    wire new_Jinkela_wire_463;
    wire new_Jinkela_wire_1441;
    wire new_Jinkela_wire_85;
    wire new_Jinkela_wire_88;
    wire new_Jinkela_wire_203;
    wire new_Jinkela_wire_669;
    wire new_Jinkela_wire_550;
    wire _145_;
    wire new_Jinkela_wire_1314;
    wire new_Jinkela_wire_1232;
    wire _109_;
    wire new_Jinkela_wire_1418;
    wire new_Jinkela_wire_396;
    wire new_Jinkela_wire_893;
    wire _233_;
    wire new_Jinkela_wire_195;
    wire new_Jinkela_wire_749;
    wire new_Jinkela_wire_1181;
    wire new_Jinkela_wire_758;
    wire new_Jinkela_wire_1358;
    wire _301_;
    wire new_Jinkela_wire_1149;
    wire new_Jinkela_wire_874;
    wire new_Jinkela_wire_29;
    wire new_Jinkela_wire_1398;
    wire new_Jinkela_wire_1254;
    wire new_Jinkela_wire_1513;
    wire _302_;
    wire new_Jinkela_wire_362;
    wire new_Jinkela_wire_1386;
    wire new_Jinkela_wire_204;
    wire new_Jinkela_wire_1566;
    wire new_Jinkela_wire_9;
    wire new_Jinkela_wire_1699;
    wire _044_;
    wire new_Jinkela_wire_112;
    wire new_Jinkela_wire_326;
    wire new_Jinkela_wire_208;
    wire new_Jinkela_wire_225;
    wire new_Jinkela_wire_142;
    wire new_Jinkela_wire_719;
    wire new_Jinkela_wire_1099;
    wire new_Jinkela_wire_484;
    wire new_Jinkela_wire_1143;
    wire _039_;
    wire _136_;
    wire new_Jinkela_wire_124;
    wire _034_;
    wire new_Jinkela_wire_222;
    wire new_Jinkela_wire_461;
    wire new_Jinkela_wire_1516;
    wire new_Jinkela_wire_1320;
    wire new_Jinkela_wire_435;
    wire new_Jinkela_wire_215;
    wire new_Jinkela_wire_1479;
    wire new_Jinkela_wire_797;
    wire _131_;
    wire new_Jinkela_wire_1324;
    wire new_Jinkela_wire_1484;
    wire new_Jinkela_wire_1632;
    wire new_Jinkela_wire_1312;
    wire new_Jinkela_wire_640;
    wire new_Jinkela_wire_1538;
    wire new_Jinkela_wire_714;
    wire new_Jinkela_wire_349;
    wire new_Jinkela_wire_1476;
    wire new_Jinkela_wire_857;
    wire _152_;
    wire new_Jinkela_wire_1250;
    wire new_Jinkela_wire_480;
    wire _019_;
    wire new_Jinkela_wire_727;
    wire new_Jinkela_wire_581;
    wire new_Jinkela_wire_4;
    wire new_Jinkela_wire_1104;
    wire new_Jinkela_wire_632;
    wire new_Jinkela_wire_164;
    wire _000_;
    wire _232_;
    wire new_Jinkela_wire_369;
    wire new_Jinkela_wire_933;
    wire new_Jinkela_wire_1459;
    wire new_Jinkela_wire_1704;
    wire new_Jinkela_wire_1174;
    wire new_Jinkela_wire_46;
    wire new_Jinkela_wire_1051;
    wire new_Jinkela_wire_1695;
    wire new_Jinkela_wire_965;
    wire new_Jinkela_wire_522;
    wire new_Jinkela_wire_35;
    wire new_Jinkela_wire_525;
    wire new_Jinkela_wire_564;
    wire new_Jinkela_wire_188;
    wire new_Jinkela_wire_383;
    wire new_Jinkela_wire_599;
    wire new_Jinkela_wire_563;
    wire new_Jinkela_wire_1336;
    wire new_Jinkela_wire_880;
    wire new_Jinkela_wire_1407;
    wire _142_;
    wire new_Jinkela_wire_319;
    wire _113_;
    wire new_Jinkela_wire_50;
    wire new_Jinkela_wire_763;
    wire _329_;
    wire new_Jinkela_wire_449;
    wire new_Jinkela_wire_1596;
    wire new_Jinkela_wire_1047;
    wire new_Jinkela_wire_569;
    wire _239_;
    wire new_Jinkela_wire_966;
    wire new_Jinkela_wire_1470;
    wire new_Jinkela_wire_608;
    wire new_Jinkela_wire_903;
    wire _078_;
    wire _185_;
    wire new_Jinkela_wire_1707;
    wire new_Jinkela_wire_698;
    wire new_Jinkela_wire_688;
    wire new_Jinkela_wire_1101;
    wire new_Jinkela_wire_452;
    wire new_Jinkela_wire_618;
    wire _336_;
    wire new_Jinkela_wire_263;
    wire _104_;
    wire new_Jinkela_wire_920;
    wire new_Jinkela_wire_625;
    wire new_Jinkela_wire_310;
    wire new_Jinkela_wire_657;
    wire _255_;
    wire new_Jinkela_wire_1288;
    wire new_Jinkela_wire_360;
    wire new_Jinkela_wire_1340;
    wire new_Jinkela_wire_424;
    wire new_Jinkela_wire_614;
    wire new_Jinkela_wire_1202;
    wire new_Jinkela_wire_1076;
    wire new_Jinkela_wire_492;
    wire new_Jinkela_wire_1451;
    wire new_Jinkela_wire_23;
    wire new_Jinkela_wire_192;
    wire new_Jinkela_wire_840;
    wire new_Jinkela_wire_311;
    wire _107_;
    wire new_Jinkela_wire_1446;
    wire new_Jinkela_wire_126;
    wire new_Jinkela_wire_1648;
    wire _244_;
    wire new_Jinkela_wire_833;
    wire new_Jinkela_wire_631;
    wire _073_;
    wire new_Jinkela_wire_1335;
    wire new_Jinkela_wire_1683;
    wire new_Jinkela_wire_540;
    wire new_Jinkela_wire_1650;
    wire new_Jinkela_wire_264;
    wire new_Jinkela_wire_594;
    wire new_Jinkela_wire_1514;
    wire new_Jinkela_wire_31;
    wire new_Jinkela_wire_1204;
    wire new_Jinkela_wire_590;
    wire new_Jinkela_wire_1285;
    wire new_Jinkela_wire_671;
    wire new_Jinkela_wire_1399;
    wire new_Jinkela_wire_337;
    wire new_Jinkela_wire_448;
    wire new_Jinkela_wire_1270;
    wire new_Jinkela_wire_1086;
    wire _209_;
    wire new_Jinkela_wire_259;
    wire new_Jinkela_wire_1360;
    wire new_Jinkela_wire_1492;
    wire new_Jinkela_wire_986;
    wire _241_;
    wire _151_;
    wire new_Jinkela_wire_1491;
    wire _341_;
    wire new_Jinkela_wire_887;
    wire new_Jinkela_wire_865;
    wire new_Jinkela_wire_781;
    wire new_Jinkela_wire_1209;
    wire new_Jinkela_wire_1141;
    wire _050_;
    wire new_Jinkela_wire_1;
    wire new_Jinkela_wire_538;
    wire new_Jinkela_wire_1165;
    wire new_Jinkela_wire_137;
    wire new_Jinkela_wire_42;
    wire new_Jinkela_wire_1318;
    wire new_Jinkela_wire_1348;
    wire new_Jinkela_wire_1579;
    wire new_Jinkela_wire_1709;
    wire new_Jinkela_wire_1629;
    wire new_Jinkela_wire_1354;
    wire new_Jinkela_wire_493;
    wire new_Jinkela_wire_173;
    wire new_Jinkela_wire_926;
    wire _318_;
    wire new_Jinkela_wire_1504;
    wire _309_;
    wire new_Jinkela_wire_1349;
    wire new_Jinkela_wire_1257;
    wire new_Jinkela_wire_806;
    wire _322_;
    wire new_Jinkela_wire_703;
    wire _074_;
    wire new_Jinkela_wire_152;
    wire _068_;
    wire new_Jinkela_wire_672;
    wire new_Jinkela_wire_235;
    wire new_Jinkela_wire_881;
    wire new_Jinkela_wire_566;
    wire new_Jinkela_wire_811;
    wire new_Jinkela_wire_898;
    wire _026_;
    wire new_Jinkela_wire_447;
    wire new_Jinkela_wire_1584;
    wire new_Jinkela_wire_161;
    wire new_Jinkela_wire_1413;
    wire new_Jinkela_wire_52;
    wire new_Jinkela_wire_1532;
    wire _092_;
    wire new_Jinkela_wire_439;
    wire new_Jinkela_wire_1073;
    wire _059_;
    wire new_Jinkela_wire_1567;
    wire _065_;
    wire _333_;
    wire new_Jinkela_wire_274;
    wire new_Jinkela_wire_1322;
    wire new_Jinkela_wire_1019;
    wire new_Jinkela_wire_705;
    wire new_Jinkela_wire_964;
    wire new_Jinkela_wire_529;
    wire new_Jinkela_wire_1547;
    wire new_Jinkela_wire_779;
    wire _224_;
    wire new_Jinkela_wire_1102;
    wire new_Jinkela_wire_223;
    wire _146_;
    wire new_Jinkela_wire_1123;
    wire new_Jinkela_wire_234;
    wire new_Jinkela_wire_1040;
    wire _226_;
    wire new_Jinkela_wire_1267;
    wire _088_;
    wire new_Jinkela_wire_121;
    wire _314_;
    wire new_Jinkela_wire_774;
    wire new_Jinkela_wire_1401;
    wire new_Jinkela_wire_60;
    wire new_Jinkela_wire_1608;
    wire new_Jinkela_wire_87;
    wire new_Jinkela_wire_1696;
    wire new_Jinkela_wire_328;
    wire new_Jinkela_wire_261;
    wire new_Jinkela_wire_1234;
    wire new_Jinkela_wire_141;
    wire new_Jinkela_wire_728;
    wire new_Jinkela_wire_1226;
    wire new_net_685;
    wire _189_;
    wire new_Jinkela_wire_430;
    wire new_Jinkela_wire_317;
    wire new_Jinkela_wire_1457;
    wire new_Jinkela_wire_34;
    wire _269_;
    wire _190_;
    wire _091_;
    wire new_Jinkela_wire_1431;
    wire new_Jinkela_wire_1179;
    wire new_Jinkela_wire_458;
    wire new_Jinkela_wire_1669;
    wire new_Jinkela_wire_394;
    wire new_Jinkela_wire_1490;
    wire new_Jinkela_wire_150;
    wire _253_;
    wire new_Jinkela_wire_1467;
    wire new_Jinkela_wire_97;
    wire new_Jinkela_wire_940;
    wire new_Jinkela_wire_513;
    wire new_Jinkela_wire_1540;
    wire new_Jinkela_wire_1592;
    wire new_Jinkela_wire_1125;
    wire new_Jinkela_wire_25;
    wire new_Jinkela_wire_1606;
    wire _220_;
    wire new_Jinkela_wire_1693;
    wire new_Jinkela_wire_1117;
    wire new_Jinkela_wire_450;
    wire new_Jinkela_wire_735;
    wire new_Jinkela_wire_1654;
    wire _060_;
    wire _135_;
    wire new_Jinkela_wire_764;
    wire new_Jinkela_wire_732;
    wire new_Jinkela_wire_1006;
    wire new_Jinkela_wire_942;
    wire new_Jinkela_wire_624;
    wire new_Jinkela_wire_1663;
    wire new_Jinkela_wire_870;
    wire new_Jinkela_wire_1501;
    wire new_Jinkela_wire_76;
    wire _085_;
    wire new_Jinkela_wire_1442;
    wire new_Jinkela_wire_1269;
    wire new_Jinkela_wire_882;
    wire new_Jinkela_wire_950;
    wire new_Jinkela_wire_825;
    wire new_Jinkela_wire_827;
    wire _358_;
    wire new_Jinkela_wire_1559;
    wire new_Jinkela_wire_1575;
    wire new_Jinkela_wire_967;
    wire new_Jinkela_wire_694;
    wire new_Jinkela_wire_1562;
    wire new_Jinkela_wire_1511;
    wire new_Jinkela_wire_908;
    wire new_Jinkela_wire_66;
    wire new_Jinkela_wire_110;
    wire new_Jinkela_wire_1522;
    wire new_Jinkela_wire_296;
    wire new_Jinkela_wire_65;
    wire new_Jinkela_wire_726;
    wire new_Jinkela_wire_165;
    wire new_Jinkela_wire_75;
    wire new_Jinkela_wire_894;
    wire _118_;
    wire new_Jinkela_wire_382;
    wire _285_;
    wire _267_;
    wire _049_;
    wire new_Jinkela_wire_101;
    wire _015_;
    wire new_Jinkela_wire_1637;
    wire new_Jinkela_wire_1640;
    wire new_Jinkela_wire_348;
    wire _231_;
    wire _111_;
    wire new_Jinkela_wire_437;
    wire new_Jinkela_wire_1278;
    wire new_Jinkela_wire_386;
    wire new_Jinkela_wire_39;
    wire new_Jinkela_wire_125;
    wire new_Jinkela_wire_1113;
    wire new_Jinkela_wire_1005;
    wire new_Jinkela_wire_792;
    wire new_Jinkela_wire_1447;
    wire new_Jinkela_wire_17;
    wire new_Jinkela_wire_1034;
    wire new_Jinkela_wire_6;
    wire new_Jinkela_wire_516;
    wire _183_;
    wire new_Jinkela_wire_403;
    wire new_Jinkela_wire_27;
    wire _045_;
    wire new_Jinkela_wire_1482;
    wire new_Jinkela_wire_925;
    wire new_Jinkela_wire_683;
    wire new_Jinkela_wire_1565;
    wire new_Jinkela_wire_104;
    wire new_Jinkela_wire_999;
    wire _296_;
    wire _317_;
    wire new_Jinkela_wire_914;
    wire new_Jinkela_wire_1017;
    wire new_Jinkela_wire_1262;
    wire new_Jinkela_wire_954;
    wire _247_;
    wire new_Jinkela_wire_557;
    wire new_Jinkela_wire_318;
    wire new_Jinkela_wire_808;
    wire new_Jinkela_wire_1077;
    wire new_Jinkela_wire_582;
    wire new_Jinkela_wire_1573;
    wire new_Jinkela_wire_959;
    wire new_Jinkela_wire_1089;
    wire _153_;
    wire _169_;
    wire new_Jinkela_wire_366;
    wire new_Jinkela_wire_1408;
    wire _098_;
    wire new_Jinkela_wire_661;
    wire new_Jinkela_wire_1518;
    wire new_Jinkela_wire_1216;
    wire new_Jinkela_wire_1347;
    wire new_Jinkela_wire_810;
    wire new_Jinkela_wire_537;
    wire new_Jinkela_wire_1214;
    wire new_Jinkela_wire_374;
    wire new_Jinkela_wire_1264;
    wire new_Jinkela_wire_578;
    wire _294_;
    wire new_Jinkela_wire_1685;
    wire new_Jinkela_wire_127;
    wire new_Jinkela_wire_292;
    wire new_Jinkela_wire_1425;
    wire new_Jinkela_wire_408;
    wire new_Jinkela_wire_47;
    wire new_Jinkela_wire_526;
    wire new_Jinkela_wire_668;
    wire new_Jinkela_wire_623;
    wire new_Jinkela_wire_139;
    wire new_Jinkela_wire_711;
    wire new_Jinkela_wire_528;
    wire new_Jinkela_wire_138;
    wire new_Jinkela_wire_803;
    wire new_Jinkela_wire_1188;
    wire new_Jinkela_wire_331;
    wire new_Jinkela_wire_1020;
    wire new_Jinkela_wire_1247;
    wire new_Jinkela_wire_1252;
    wire _265_;
    wire new_Jinkela_wire_187;
    wire new_Jinkela_wire_237;
    wire new_Jinkela_wire_1527;
    wire new_Jinkela_wire_1100;
    wire new_Jinkela_wire_1107;
    wire new_Jinkela_wire_713;
    wire new_Jinkela_wire_693;
    wire new_Jinkela_wire_1461;
    wire _205_;
    wire new_Jinkela_wire_217;
    wire new_Jinkela_wire_190;
    wire new_Jinkela_wire_1372;
    wire new_Jinkela_wire_1109;
    wire new_Jinkela_wire_610;
    wire new_Jinkela_wire_679;
    wire new_Jinkela_wire_638;
    wire new_Jinkela_wire_796;
    wire new_Jinkela_wire_570;
    wire new_Jinkela_wire_1406;
    wire new_Jinkela_wire_505;
    wire new_Jinkela_wire_262;
    wire new_Jinkela_wire_1093;
    wire new_net_689;
    wire new_Jinkela_wire_1292;
    wire new_Jinkela_wire_1448;
    wire new_Jinkela_wire_822;
    wire new_Jinkela_wire_572;
    wire new_Jinkela_wire_1439;
    wire new_Jinkela_wire_1675;
    wire new_Jinkela_wire_1369;
    wire new_Jinkela_wire_1488;
    wire new_Jinkela_wire_189;
    wire new_Jinkela_wire_1390;
    wire new_Jinkela_wire_107;
    wire _197_;
    wire new_Jinkela_wire_169;
    wire new_Jinkela_wire_1558;
    wire _156_;
    wire new_Jinkela_wire_1655;
    wire _016_;
    wire new_Jinkela_wire_1383;
    wire new_Jinkela_wire_790;
    wire new_Jinkela_wire_456;
    wire new_Jinkela_wire_1280;
    wire new_Jinkela_wire_816;
    wire new_Jinkela_wire_1697;
    wire new_Jinkela_wire_340;
    wire new_net_705;
    wire new_Jinkela_wire_1018;
    wire new_net_709;
    wire new_Jinkela_wire_460;
    wire _066_;
    wire new_Jinkela_wire_1045;
    wire new_Jinkela_wire_1563;
    wire new_Jinkela_wire_92;
    wire new_Jinkela_wire_1330;
    wire new_Jinkela_wire_800;
    wire new_Jinkela_wire_506;
    wire new_Jinkela_wire_3;
    wire new_Jinkela_wire_1233;
    wire new_Jinkela_wire_576;
    wire new_Jinkela_wire_1661;
    wire new_Jinkela_wire_1284;
    wire _171_;
    wire new_Jinkela_wire_960;
    wire new_Jinkela_wire_814;
    wire new_Jinkela_wire_1075;
    wire new_Jinkela_wire_14;
    wire new_Jinkela_wire_855;
    wire new_Jinkela_wire_1658;
    wire new_Jinkela_wire_151;
    wire _352_;
    wire new_Jinkela_wire_155;
    wire new_Jinkela_wire_199;
    wire new_Jinkela_wire_1027;
    wire new_Jinkela_wire_995;
    wire new_Jinkela_wire_477;
    wire new_Jinkela_wire_197;
    wire _286_;
    wire new_Jinkela_wire_91;
    wire new_Jinkela_wire_1136;
    wire _140_;
    wire new_Jinkela_wire_109;
    wire new_Jinkela_wire_532;
    wire _194_;
    wire new_Jinkela_wire_743;
    wire new_Jinkela_wire_1642;
    wire new_Jinkela_wire_445;
    wire new_Jinkela_wire_1523;
    wire new_Jinkela_wire_345;
    wire new_Jinkela_wire_1664;
    wire new_Jinkela_wire_1151;
    wire new_Jinkela_wire_482;
    wire new_Jinkela_wire_715;
    wire new_Jinkela_wire_918;
    wire new_Jinkela_wire_1485;
    wire new_Jinkela_wire_996;
    wire new_Jinkela_wire_1597;
    wire new_Jinkela_wire_1409;
    wire _179_;
    wire new_Jinkela_wire_1087;
    wire _276_;
    wire new_Jinkela_wire_983;
    wire new_Jinkela_wire_1163;
    wire new_Jinkela_wire_1434;
    wire new_Jinkela_wire_28;
    wire new_Jinkela_wire_346;
    wire new_Jinkela_wire_724;
    wire new_Jinkela_wire_1542;
    wire new_Jinkela_wire_24;
    wire new_Jinkela_wire_1387;
    wire new_Jinkela_wire_268;
    wire _017_;
    wire new_Jinkela_wire_1580;
    wire new_Jinkela_wire_656;
    wire new_Jinkela_wire_19;
    wire new_Jinkela_wire_686;
    wire new_Jinkela_wire_1297;
    wire new_Jinkela_wire_1166;
    wire new_Jinkela_wire_1646;
    wire new_Jinkela_wire_1258;
    wire _327_;
    wire _237_;
    wire _259_;
    wire new_Jinkela_wire_105;
    wire new_Jinkela_wire_1160;
    wire _121_;
    wire new_Jinkela_wire_1126;
    wire new_Jinkela_wire_611;
    wire new_Jinkela_wire_1487;
    wire new_Jinkela_wire_1393;
    wire new_Jinkela_wire_745;
    wire new_Jinkela_wire_759;
    wire new_Jinkela_wire_175;
    wire new_Jinkela_wire_936;
    wire new_Jinkela_wire_1142;
    wire new_Jinkela_wire_160;
    wire _348_;
    wire _216_;
    wire new_Jinkela_wire_975;
    wire new_Jinkela_wire_1703;
    wire new_Jinkela_wire_1009;
    wire new_Jinkela_wire_1055;
    wire new_Jinkela_wire_335;
    wire new_Jinkela_wire_912;
    wire _112_;
    wire new_Jinkela_wire_1189;
    wire _347_;
    wire _057_;
    wire new_Jinkela_wire_915;
    wire new_Jinkela_wire_1296;
    wire new_Jinkela_wire_634;
    wire new_Jinkela_wire_271;
    wire new_Jinkela_wire_1351;
    wire new_Jinkela_wire_1154;
    wire new_Jinkela_wire_616;
    wire _014_;
    wire _023_;
    wire new_Jinkela_wire_641;
    wire new_Jinkela_wire_1489;
    wire new_Jinkela_wire_1578;
    wire new_Jinkela_wire_149;
    wire new_Jinkela_wire_744;
    wire new_Jinkela_wire_1032;
    wire new_Jinkela_wire_136;
    wire new_Jinkela_wire_818;
    wire new_Jinkela_wire_38;
    wire new_Jinkela_wire_560;
    wire new_Jinkela_wire_1035;
    wire new_Jinkela_wire_33;
    wire _304_;
    wire new_Jinkela_wire_1236;
    wire new_Jinkela_wire_891;
    wire new_Jinkela_wire_1283;
    wire _213_;
    wire new_Jinkela_wire_11;
    wire _103_;
    wire new_net_713;
    wire new_Jinkela_wire_209;
    wire new_Jinkela_wire_191;
    wire new_Jinkela_wire_583;
    wire new_Jinkela_wire_1177;
    wire new_Jinkela_wire_923;
    wire new_Jinkela_wire_1028;
    wire _198_;
    wire _125_;
    wire new_Jinkela_wire_316;
    wire new_Jinkela_wire_843;
    wire new_Jinkela_wire_322;
    wire new_Jinkela_wire_178;
    wire new_Jinkela_wire_1463;
    wire new_Jinkela_wire_909;
    wire new_Jinkela_wire_1537;
    wire new_Jinkela_wire_1274;
    wire new_Jinkela_wire_981;
    wire new_Jinkela_wire_106;
    wire new_Jinkela_wire_849;
    wire _225_;
    wire _242_;
    wire new_Jinkela_wire_1066;
    wire new_Jinkela_wire_353;
    wire new_Jinkela_wire_80;
    wire _227_;
    wire _344_;
    wire new_Jinkela_wire_236;
    wire new_Jinkela_wire_575;
    wire new_Jinkela_wire_1557;
    wire new_Jinkela_wire_113;
    wire new_Jinkela_wire_832;
    wire _117_;
    wire _128_;
    wire new_Jinkela_wire_181;
    wire new_Jinkela_wire_1609;
    wire new_Jinkela_wire_140;
    wire new_Jinkela_wire_387;
    wire new_Jinkela_wire_401;
    wire new_Jinkela_wire_637;
    wire new_Jinkela_wire_381;
    wire new_Jinkela_wire_156;
    wire new_Jinkela_wire_606;
    wire new_Jinkela_wire_1276;
    wire new_Jinkela_wire_929;
    wire new_Jinkela_wire_405;
    wire _147_;
    wire new_Jinkela_wire_499;
    wire new_Jinkela_wire_1623;
    wire new_Jinkela_wire_247;
    wire new_Jinkela_wire_1405;
    wire new_Jinkela_wire_12;
    wire new_Jinkela_wire_211;
    wire new_Jinkela_wire_409;
    wire new_Jinkela_wire_1302;
    wire new_Jinkela_wire_147;
    wire new_Jinkela_wire_1545;
    wire new_Jinkela_wire_1310;
    wire new_Jinkela_wire_597;
    wire new_Jinkela_wire_600;
    wire new_Jinkela_wire_356;
    wire new_Jinkela_wire_1456;
    wire new_Jinkela_wire_69;
    wire new_Jinkela_wire_90;
    wire new_Jinkela_wire_1067;
    wire _235_;
    wire new_Jinkela_wire_530;
    wire new_Jinkela_wire_419;
    wire new_Jinkela_wire_861;
    wire new_Jinkela_wire_1255;
    wire new_Jinkela_wire_1572;
    wire new_Jinkela_wire_1198;
    wire new_Jinkela_wire_896;
    wire _148_;
    wire new_Jinkela_wire_1493;
    wire _251_;
    wire new_Jinkela_wire_1094;
    wire new_Jinkela_wire_158;
    wire _122_;
    wire new_Jinkela_wire_249;
    wire new_Jinkela_wire_205;
    wire new_Jinkela_wire_1249;
    wire new_Jinkela_wire_1208;
    wire new_Jinkela_wire_122;
    wire _229_;
    wire new_Jinkela_wire_1319;
    wire new_Jinkela_wire_1619;
    wire new_Jinkela_wire_1024;
    wire new_Jinkela_wire_1152;
    wire new_Jinkela_wire_1635;
    wire new_Jinkela_wire_751;
    wire new_Jinkela_wire_1295;
    wire new_Jinkela_wire_826;
    wire new_Jinkela_wire_114;
    wire new_Jinkela_wire_947;
    wire new_Jinkela_wire_1679;
    wire new_Jinkela_wire_1571;
    wire new_Jinkela_wire_200;
    wire _011_;
    wire new_Jinkela_wire_976;
    wire new_Jinkela_wire_1694;
    wire new_Jinkela_wire_455;
    wire new_Jinkela_wire_473;
    wire new_Jinkela_wire_1626;
    wire _032_;
    wire new_Jinkela_wire_788;
    wire new_Jinkela_wire_1607;
    wire new_Jinkela_wire_218;
    wire new_Jinkela_wire_1164;
    wire new_Jinkela_wire_1465;
    wire _342_;
    wire _010_;
    wire new_Jinkela_wire_1155;
    wire new_Jinkela_wire_1698;
    wire new_Jinkela_wire_1145;
    wire _086_;
    wire _030_;
    wire new_Jinkela_wire_1605;
    wire new_Jinkela_wire_472;
    wire new_Jinkela_wire_1306;
    wire new_Jinkela_wire_1455;
    wire new_Jinkela_wire_228;
    wire _139_;
    wire new_Jinkela_wire_741;
    wire _272_;
    wire new_Jinkela_wire_977;
    wire new_Jinkela_wire_1478;
    wire new_Jinkela_wire_423;
    wire new_Jinkela_wire_1373;
    wire new_Jinkela_wire_598;
    wire new_Jinkela_wire_1060;
    wire new_Jinkela_wire_982;
    wire new_Jinkela_wire_1229;
    wire new_Jinkela_wire_941;
    wire _130_;
    wire new_Jinkela_wire_1589;
    wire new_Jinkela_wire_1253;
    wire new_Jinkela_wire_1054;
    wire new_Jinkela_wire_1473;
    wire new_Jinkela_wire_339;
    wire new_Jinkela_wire_459;
    wire _106_;
    wire _290_;
    wire _006_;
    wire new_Jinkela_wire_1220;
    wire _313_;
    wire new_Jinkela_wire_1328;
    wire new_Jinkela_wire_1423;
    wire new_Jinkela_wire_762;
    wire new_Jinkela_wire_533;
    wire new_Jinkela_wire_1604;
    wire new_Jinkela_wire_813;
    wire new_Jinkela_wire_1011;
    wire new_Jinkela_wire_1172;
    wire new_Jinkela_wire_567;
    wire new_Jinkela_wire_1341;
    wire new_Jinkela_wire_415;
    wire new_Jinkela_wire_1612;
    wire _335_;
    wire new_Jinkela_wire_98;
    wire new_Jinkela_wire_946;
    wire new_Jinkela_wire_1178;
    wire new_Jinkela_wire_615;
    wire new_Jinkela_wire_413;
    wire new_Jinkela_wire_303;
    wire new_Jinkela_wire_771;
    wire _082_;
    wire _316_;
    wire new_Jinkela_wire_62;
    wire new_Jinkela_wire_1415;
    wire new_Jinkela_wire_336;
    wire new_Jinkela_wire_1211;
    wire new_Jinkela_wire_1552;
    wire new_Jinkela_wire_691;
    wire new_Jinkela_wire_1235;
    wire new_Jinkela_wire_824;
    wire new_Jinkela_wire_134;
    wire new_Jinkela_wire_1068;
    wire new_Jinkela_wire_365;
    wire new_Jinkela_wire_1682;
    wire new_Jinkela_wire_696;
    wire new_Jinkela_wire_233;
    wire new_Jinkela_wire_1477;
    wire new_Jinkela_wire_1676;
    wire new_Jinkela_wire_426;
    wire new_Jinkela_wire_251;
    wire new_Jinkela_wire_341;
    wire new_Jinkela_wire_508;
    wire _191_;
    wire new_Jinkela_wire_978;
    wire new_Jinkela_wire_420;
    wire new_Jinkela_wire_1167;
    wire _097_;
    wire new_Jinkela_wire_1213;
    wire new_Jinkela_wire_692;
    wire new_Jinkela_wire_838;
    wire _162_;
    wire new_Jinkela_wire_706;
    wire new_Jinkela_wire_309;
    wire _160_;
    wire new_Jinkela_wire_507;
    wire new_Jinkela_wire_1498;
    wire new_Jinkela_wire_773;
    wire new_Jinkela_wire_327;
    wire new_Jinkela_wire_601;
    wire new_Jinkela_wire_587;
    wire new_Jinkela_wire_1097;
    wire new_Jinkela_wire_377;
    wire new_Jinkela_wire_710;
    wire _208_;
    wire new_Jinkela_wire_1108;
    wire new_Jinkela_wire_1338;
    wire new_Jinkela_wire_130;
    wire new_Jinkela_wire_306;
    wire _303_;
    wire new_Jinkela_wire_299;
    wire new_Jinkela_wire_1416;
    wire new_Jinkela_wire_255;
    wire new_Jinkela_wire_775;
    wire _013_;
    wire _266_;
    wire new_Jinkela_wire_1301;
    wire new_Jinkela_wire_485;
    wire new_Jinkela_wire_1613;
    wire new_Jinkela_wire_1617;
    wire new_Jinkela_wire_544;
    wire new_Jinkela_wire_1217;
    wire new_Jinkela_wire_129;
    wire new_Jinkela_wire_244;
    wire new_Jinkela_wire_828;
    wire new_Jinkela_wire_1105;
    wire new_Jinkela_wire_989;
    wire new_Jinkela_wire_804;
    wire _261_;
    wire new_Jinkela_wire_131;
    wire new_Jinkela_wire_1098;
    wire new_Jinkela_wire_648;
    wire new_Jinkela_wire_738;
    wire new_Jinkela_wire_1289;
    wire new_Jinkela_wire_361;
    wire _201_;
    wire new_Jinkela_wire_531;
    wire new_Jinkela_wire_302;
    wire new_Jinkela_wire_1508;
    wire new_Jinkela_wire_534;
    wire new_Jinkela_wire_1096;
    wire new_Jinkela_wire_1657;
    wire new_Jinkela_wire_612;
    wire new_Jinkela_wire_1268;
    wire new_Jinkela_wire_64;
    wire new_Jinkela_wire_392;
    wire _069_;
    wire new_Jinkela_wire_1334;
    wire _199_;
    wire new_Jinkela_wire_1013;
    wire new_Jinkela_wire_1137;
    wire _105_;
    wire new_Jinkela_wire_414;
    wire new_Jinkela_wire_399;
    wire new_Jinkela_wire_1042;
    wire _321_;
    wire new_Jinkela_wire_1303;
    wire new_Jinkela_wire_1355;
    wire _203_;
    wire new_Jinkela_wire_520;
    wire new_Jinkela_wire_1591;
    wire _062_;
    wire new_Jinkela_wire_378;
    wire new_Jinkela_wire_766;
    wire new_Jinkela_wire_500;
    wire _351_;
    wire new_Jinkela_wire_1687;
    wire _095_;
    wire new_Jinkela_wire_210;
    wire new_Jinkela_wire_1618;
    wire new_Jinkela_wire_712;
    wire new_Jinkela_wire_1317;
    wire new_Jinkela_wire_404;
    wire new_Jinkela_wire_593;
    wire new_Jinkela_wire_363;
    wire new_Jinkela_wire_1410;
    wire new_Jinkela_wire_379;
    wire new_Jinkela_wire_892;
    wire new_Jinkela_wire_1525;
    wire new_Jinkela_wire_588;
    wire new_Jinkela_wire_179;
    wire new_Jinkela_wire_418;
    wire new_Jinkela_wire_457;
    wire _360_;
    wire new_Jinkela_wire_1367;
    wire new_Jinkela_wire_1644;
    wire new_Jinkela_wire_1180;
    wire new_Jinkela_wire_1187;
    wire new_Jinkela_wire_1161;
    wire new_Jinkela_wire_1199;
    wire _218_;
    wire new_Jinkela_wire_1357;
    wire new_Jinkela_wire_146;
    wire _090_;
    wire new_Jinkela_wire_1397;
    wire new_Jinkela_wire_390;
    wire _274_;
    wire new_Jinkela_wire_279;
    wire _359_;
    wire new_Jinkela_wire_1215;
    wire new_Jinkela_wire_1362;
    wire new_Jinkela_wire_911;
    wire new_Jinkela_wire_812;
    wire new_Jinkela_wire_1110;
    wire new_Jinkela_wire_1481;
    wire new_Jinkela_wire_646;
    wire _215_;
    wire new_Jinkela_wire_144;
    wire new_Jinkela_wire_900;
    wire new_Jinkela_wire_194;
    wire new_Jinkela_wire_185;
    wire new_Jinkela_wire_1069;
    wire new_net_715;
    wire new_Jinkela_wire_1326;
    wire new_Jinkela_wire_1417;
    wire new_Jinkela_wire_1505;
    wire new_Jinkela_wire_768;
    wire _061_;
    wire new_Jinkela_wire_1171;
    wire new_Jinkela_wire_815;
    wire _009_;
    wire _212_;
    wire new_Jinkela_wire_417;
    wire new_Jinkela_wire_651;
    wire new_Jinkela_wire_1483;
    wire new_Jinkela_wire_63;
    wire _141_;
    wire new_Jinkela_wire_649;
    wire new_Jinkela_wire_586;
    wire new_Jinkela_wire_1294;
    wire _063_;
    wire new_Jinkela_wire_1702;
    wire _188_;
    wire new_Jinkela_wire_1200;
    wire _170_;
    wire new_Jinkela_wire_1038;
    wire new_Jinkela_wire_305;
    wire new_Jinkela_wire_1462;
    wire new_Jinkela_wire_364;
    wire new_Jinkela_wire_1224;
    wire _292_;
    wire new_Jinkela_wire_1353;
    wire new_Jinkela_wire_1345;
    wire new_Jinkela_wire_1191;
    wire new_Jinkela_wire_676;
    wire new_Jinkela_wire_658;
    wire new_Jinkela_wire_1588;
    wire new_Jinkela_wire_1056;
    wire new_Jinkela_wire_1576;
    wire _099_;
    wire new_Jinkela_wire_1036;
    wire _258_;
    wire new_Jinkela_wire_1652;
    wire new_Jinkela_wire_347;
    wire new_Jinkela_wire_1615;
    wire new_Jinkela_wire_1420;
    wire new_Jinkela_wire_16;
    wire new_Jinkela_wire_55;
    wire new_Jinkela_wire_633;
    wire new_Jinkela_wire_416;
    wire _353_;
    wire new_Jinkela_wire_1282;
    wire new_Jinkela_wire_332;
    wire new_Jinkela_wire_1705;
    wire new_Jinkela_wire_254;
    wire new_Jinkela_wire_552;
    wire new_Jinkela_wire_780;
    wire new_Jinkela_wire_1526;
    wire new_Jinkela_wire_650;
    wire new_Jinkela_wire_275;
    wire new_Jinkela_wire_723;
    wire _058_;
    wire new_Jinkela_wire_957;
    wire new_Jinkela_wire_895;
    wire _299_;
    wire new_Jinkela_wire_68;
    wire new_Jinkela_wire_997;
    wire new_Jinkela_wire_216;
    wire new_Jinkela_wire_699;
    wire new_Jinkela_wire_752;
    wire new_Jinkela_wire_10;
    wire _172_;
    wire _192_;
    wire new_Jinkela_wire_78;
    wire new_Jinkela_wire_939;
    wire new_Jinkela_wire_1645;
    wire new_Jinkela_wire_100;
    wire new_Jinkela_wire_307;
    wire new_Jinkela_wire_1259;
    wire new_Jinkela_wire_820;
    wire new_Jinkela_wire_750;
    wire new_Jinkela_wire_1432;
    wire new_Jinkela_wire_388;
    wire new_Jinkela_wire_504;
    wire new_Jinkela_wire_733;
    wire _159_;
    wire _094_;
    wire new_Jinkela_wire_519;
    wire new_Jinkela_wire_626;
    wire new_Jinkela_wire_545;
    wire new_Jinkela_wire_602;
    wire new_Jinkela_wire_1004;
    wire new_Jinkela_wire_1120;
    wire new_Jinkela_wire_897;
    wire new_Jinkela_wire_342;
    wire new_Jinkela_wire_434;
    wire _070_;
    wire new_Jinkela_wire_257;
    wire new_Jinkela_wire_95;
    wire new_Jinkela_wire_509;
    wire _067_;
    wire new_Jinkela_wire_496;
    wire new_Jinkela_wire_725;
    wire new_Jinkela_wire_1132;
    wire new_Jinkela_wire_1681;
    wire new_Jinkela_wire_1660;
    wire new_Jinkela_wire_888;
    wire new_Jinkela_wire_605;
    wire new_Jinkela_wire_1691;
    wire _248_;
    wire new_Jinkela_wire_304;
    wire new_Jinkela_wire_1561;
    wire new_Jinkela_wire_1272;
    wire new_Jinkela_wire_355;
    wire new_Jinkela_wire_907;
    wire _291_;
    wire new_Jinkela_wire_559;
    wire new_Jinkela_wire_230;
    wire new_Jinkela_wire_1503;
    wire _324_;
    wire new_Jinkela_wire_1402;
    wire new_Jinkela_wire_269;
    wire _361_;
    wire new_Jinkela_wire_1299;
    wire new_Jinkela_wire_984;
    wire new_Jinkela_wire_830;
    wire new_Jinkela_wire_1428;
    wire new_Jinkela_wire_166;
    wire new_Jinkela_wire_853;
    wire new_Jinkela_wire_278;
    wire new_Jinkela_wire_1453;
    wire new_Jinkela_wire_375;
    wire new_Jinkela_wire_1173;
    wire new_Jinkela_wire_171;
    wire new_Jinkela_wire_412;
    wire new_Jinkela_wire_454;
    wire new_Jinkela_wire_1548;
    wire _307_;
    wire new_Jinkela_wire_791;
    wire new_Jinkela_wire_300;
    wire new_Jinkela_wire_325;
    wire new_Jinkela_wire_1411;
    wire _168_;
    wire new_Jinkela_wire_370;
    wire new_Jinkela_wire_123;
    wire new_Jinkela_wire_609;
    wire _079_;
    wire _257_;
    wire new_Jinkela_wire_1365;
    wire new_Jinkela_wire_1001;
    wire new_Jinkela_wire_272;
    wire new_Jinkela_wire_603;
    wire _315_;
    wire new_Jinkela_wire_635;
    wire new_Jinkela_wire_1346;
    wire new_Jinkela_wire_400;
    wire new_Jinkela_wire_1585;
    wire new_Jinkela_wire_1205;
    wire new_Jinkela_wire_884;
    wire new_Jinkela_wire_595;
    wire new_Jinkela_wire_910;
    wire new_Jinkela_wire_241;
    wire _134_;
    wire new_Jinkela_wire_1667;
    wire new_Jinkela_wire_1190;
    wire new_Jinkela_wire_1091;
    wire _077_;
    wire new_Jinkela_wire_93;
    wire new_Jinkela_wire_281;
    wire new_Jinkela_wire_930;
    wire _300_;
    wire new_Jinkela_wire_51;
    wire _196_;
    wire new_Jinkela_wire_568;
    wire new_Jinkela_wire_1680;
    wire new_Jinkela_wire_501;
    wire _343_;
    wire new_Jinkela_wire_917;
    wire new_Jinkela_wire_2;
    wire new_Jinkela_wire_675;
    wire new_Jinkela_wire_1512;
    wire new_Jinkela_wire_1555;
    wire new_Jinkela_wire_1339;
    wire new_Jinkela_wire_1148;
    wire _155_;
    wire _268_;
    wire new_Jinkela_wire_579;
    wire new_Jinkela_wire_1203;
    wire new_Jinkela_wire_1079;
    wire new_Jinkela_wire_1129;
    wire new_Jinkela_wire_58;
    wire new_Jinkela_wire_1659;
    wire new_Jinkela_wire_1321;
    wire new_Jinkela_wire_1686;
    wire new_Jinkela_wire_1590;
    wire new_Jinkela_wire_620;
    wire new_Jinkela_wire_817;
    wire new_Jinkela_wire_1238;
    wire new_Jinkela_wire_320;
    wire new_Jinkela_wire_858;
    wire new_Jinkela_wire_1529;
    wire _357_;
    wire new_Jinkela_wire_863;
    wire new_Jinkela_wire_1041;
    wire new_Jinkela_wire_841;
    wire new_Jinkela_wire_380;
    wire _157_;
    wire new_Jinkela_wire_1510;
    wire new_Jinkela_wire_1437;
    wire new_Jinkela_wire_1472;
    wire new_Jinkela_wire_844;
    wire _080_;
    wire new_Jinkela_wire_998;
    wire new_Jinkela_wire_436;
    wire new_Jinkela_wire_877;
    wire new_Jinkela_wire_944;
    wire new_Jinkela_wire_1185;
    wire new_Jinkela_wire_490;
    wire new_Jinkela_wire_128;
    wire new_Jinkela_wire_889;
    wire new_Jinkela_wire_1582;
    wire new_Jinkela_wire_718;
    wire new_Jinkela_wire_267;
    wire new_Jinkela_wire_1541;
    wire new_Jinkela_wire_1391;
    wire _175_;
    wire new_Jinkela_wire_481;
    wire new_Jinkela_wire_1240;
    wire new_Jinkela_wire_277;
    wire new_Jinkela_wire_697;
    wire new_Jinkela_wire_1688;
    wire new_Jinkela_wire_1230;
    wire new_Jinkela_wire_1201;
    wire new_Jinkela_wire_783;
    wire new_Jinkela_wire_856;
    wire new_Jinkela_wire_1084;
    wire new_Jinkela_wire_1429;
    wire new_Jinkela_wire_89;
    wire new_Jinkela_wire_373;
    wire _043_;
    wire new_Jinkela_wire_1625;
    wire new_Jinkela_wire_245;
    wire new_Jinkela_wire_868;
    wire new_Jinkela_wire_153;
    wire new_Jinkela_wire_1598;
    wire new_Jinkela_wire_794;
    wire new_Jinkela_wire_1140;
    wire new_Jinkela_wire_358;
    wire _163_;
    wire new_Jinkela_wire_115;
    wire _311_;
    wire new_Jinkela_wire_1497;
    wire new_Jinkela_wire_1690;
    wire new_Jinkela_wire_240;
    wire _186_;
    wire new_Jinkela_wire_1176;
    wire new_Jinkela_wire_859;
    wire new_Jinkela_wire_489;
    wire new_Jinkela_wire_1587;
    wire new_Jinkela_wire_202;
    wire new_Jinkela_wire_70;
    wire new_Jinkela_wire_739;
    wire _064_;
    wire new_Jinkela_wire_1194;
    wire new_Jinkela_wire_1474;
    wire new_Jinkela_wire_971;
    wire new_Jinkela_wire_556;
    wire _150_;
    wire new_Jinkela_wire_1010;
    wire new_Jinkela_wire_886;
    wire _001_;
    wire new_Jinkela_wire_1023;
    wire new_Jinkela_wire_421;
    wire new_Jinkela_wire_795;
    wire _154_;
    wire new_Jinkela_wire_577;
    wire new_Jinkela_wire_1308;
    wire new_Jinkela_wire_250;
    wire new_Jinkela_wire_1539;
    wire _349_;
    wire new_Jinkela_wire_970;
    wire new_Jinkela_wire_1424;
    wire new_Jinkela_wire_663;
    wire _123_;
    wire new_Jinkela_wire_961;
    wire new_Jinkela_wire_682;
    wire _278_;
    wire new_Jinkela_wire_1026;
    wire new_Jinkela_wire_1674;
    wire new_Jinkela_wire_1184;
    wire new_Jinkela_wire_596;
    wire _051_;
    wire new_Jinkela_wire_1157;
    wire new_Jinkela_wire_428;
    wire new_Jinkela_wire_515;
    wire new_Jinkela_wire_1127;
    wire new_Jinkela_wire_799;
    wire new_Jinkela_wire_1466;
    wire new_Jinkela_wire_553;
    wire new_Jinkela_wire_1290;
    wire new_Jinkela_wire_1281;
    wire new_Jinkela_wire_1248;
    wire new_Jinkela_wire_289;
    wire new_Jinkela_wire_770;
    wire new_Jinkela_wire_802;
    wire new_Jinkela_wire_389;
    wire new_Jinkela_wire_1090;
    wire _295_;
    wire new_Jinkela_wire_18;
    wire new_Jinkela_wire_1206;
    wire new_Jinkela_wire_1237;
    wire new_Jinkela_wire_717;
    wire new_Jinkela_wire_1012;
    wire new_Jinkela_wire_834;
    wire new_Jinkela_wire_1144;
    wire new_Jinkela_wire_1636;
    wire new_Jinkela_wire_201;
    wire new_Jinkela_wire_1356;
    wire new_Jinkela_wire_221;
    wire new_Jinkela_wire_1156;
    wire _129_;
    wire new_Jinkela_wire_1059;
    wire new_Jinkela_wire_1325;
    wire new_Jinkela_wire_1196;
    wire new_Jinkela_wire_1665;
    wire new_Jinkela_wire_1150;
    wire new_Jinkela_wire_1560;
    wire _281_;
    wire new_Jinkela_wire_622;
    wire new_Jinkela_wire_1710;
    wire new_Jinkela_wire_270;
    wire new_Jinkela_wire_869;
    wire _330_;
    wire new_Jinkela_wire_333;
    wire new_Jinkela_wire_1192;
    wire new_Jinkela_wire_760;
    wire new_Jinkela_wire_1624;
    wire new_Jinkela_wire_846;
    wire new_Jinkela_wire_330;
    wire new_Jinkela_wire_742;
    wire _221_;
    wire _178_;
    wire new_Jinkela_wire_96;
    wire new_Jinkela_wire_291;
    wire new_Jinkela_wire_1331;
    wire new_Jinkela_wire_1002;
    wire new_Jinkela_wire_1610;
    wire new_Jinkela_wire_1396;
    wire new_Jinkela_wire_1231;
    wire _211_;
    wire new_Jinkela_wire_607;
    wire new_Jinkela_wire_1543;
    wire new_Jinkela_wire_132;
    wire _035_;
    wire new_Jinkela_wire_99;
    wire _165_;
    wire new_Jinkela_wire_1531;
    wire new_Jinkela_wire_1421;
    wire _176_;
    wire new_Jinkela_wire_36;
    wire _222_;
    wire _007_;
    wire new_Jinkela_wire_1469;
    wire new_Jinkela_wire_120;
    wire new_Jinkela_wire_617;
    wire new_Jinkela_wire_1138;
    wire new_Jinkela_wire_1611;
    wire new_Jinkela_wire_372;
    wire _355_;
    wire new_Jinkela_wire_757;
    wire new_Jinkela_wire_1333;
    wire _310_;
    input N97;
    input N113;
    input N73;
    input N134;
    input N57;
    input N77;
    input N17;
    input N49;
    input N93;
    input N1;
    input N131;
    input N25;
    input N109;
    input N45;
    input N132;
    input N135;
    input N61;
    input N85;
    input N117;
    input N21;
    input N33;
    input N101;
    input N81;
    input N105;
    input N41;
    input N5;
    input N130;
    input N133;
    input N89;
    input N125;
    input N53;
    input N69;
    input N29;
    input N121;
    input N9;
    input N13;
    input N137;
    input N37;
    input N136;
    input N129;
    input N65;
    output N750;
    output N738;
    output N755;
    output N736;
    output N754;
    output N731;
    output N726;
    output N740;
    output N728;
    output N752;
    output N745;
    output N733;
    output N753;
    output N739;
    output N747;
    output N724;
    output N743;
    output N737;
    output N735;
    output N727;
    output N742;
    output N741;
    output N749;
    output N734;
    output N751;
    output N725;
    output N729;
    output N748;
    output N744;
    output N732;
    output N746;
    output N730;

    or_bb _559_ (
        .a(new_Jinkela_wire_1475),
        .b(new_Jinkela_wire_1594),
        .c(_171_)
    );

    or_ii _560_ (
        .a(new_Jinkela_wire_1474),
        .b(new_Jinkela_wire_1593),
        .c(_172_)
    );

    or_ii _561_ (
        .a(new_Jinkela_wire_1660),
        .b(new_Jinkela_wire_1503),
        .c(_173_)
    );

    or_bb _562_ (
        .a(new_Jinkela_wire_1347),
        .b(new_Jinkela_wire_1236),
        .c(_174_)
    );

    and_bi _563_ (
        .a(_173_),
        .b(new_Jinkela_wire_1138),
        .c(_175_)
    );

    and_bi _564_ (
        .a(_170_),
        .b(new_Jinkela_wire_1682),
        .c(_176_)
    );

    and_bi _565_ (
        .a(new_Jinkela_wire_1),
        .b(new_Jinkela_wire_39),
        .c(_177_)
    );

    and_bi _566_ (
        .a(new_Jinkela_wire_38),
        .b(new_Jinkela_wire_4),
        .c(_178_)
    );

    or_bb _567_ (
        .a(_178_),
        .b(_177_),
        .c(_179_)
    );

    or_ii _568_ (
        .a(new_Jinkela_wire_770),
        .b(new_Jinkela_wire_1048),
        .c(_180_)
    );

    or_bi _569_ (
        .a(new_Jinkela_wire_630),
        .b(new_Jinkela_wire_1101),
        .c(_181_)
    );

    and_bi _570_ (
        .a(new_Jinkela_wire_634),
        .b(new_Jinkela_wire_1097),
        .c(_182_)
    );

    and_bi _571_ (
        .a(_181_),
        .b(_182_),
        .c(_183_)
    );

    and_bi _572_ (
        .a(new_Jinkela_wire_1471),
        .b(new_Jinkela_wire_1344),
        .c(_184_)
    );

    and_bi _573_ (
        .a(new_Jinkela_wire_1343),
        .b(new_Jinkela_wire_1470),
        .c(_185_)
    );

    or_bb _574_ (
        .a(_185_),
        .b(_184_),
        .c(_186_)
    );

    or_bb _575_ (
        .a(new_Jinkela_wire_1687),
        .b(new_Jinkela_wire_1518),
        .c(_187_)
    );

    and_bb _576_ (
        .a(new_Jinkela_wire_1686),
        .b(new_Jinkela_wire_1517),
        .c(_188_)
    );

    and_bi _577_ (
        .a(_187_),
        .b(_188_),
        .c(_189_)
    );

    or_bb _578_ (
        .a(new_Jinkela_wire_1627),
        .b(new_Jinkela_wire_1589),
        .c(_190_)
    );

    and_bb _579_ (
        .a(new_Jinkela_wire_1626),
        .b(new_Jinkela_wire_1588),
        .c(_191_)
    );

    and_bi _580_ (
        .a(_190_),
        .b(_191_),
        .c(_192_)
    );

    or_bi _581_ (
        .a(new_Jinkela_wire_1433),
        .b(new_Jinkela_wire_1662),
        .c(_193_)
    );

    and_bi _582_ (
        .a(new_Jinkela_wire_1432),
        .b(new_Jinkela_wire_1661),
        .c(_194_)
    );

    and_bi _583_ (
        .a(new_Jinkela_wire_1298),
        .b(new_Jinkela_wire_1513),
        .c(_195_)
    );

    and_bi _584_ (
        .a(new_Jinkela_wire_596),
        .b(new_Jinkela_wire_496),
        .c(_196_)
    );

    and_bi _585_ (
        .a(new_Jinkela_wire_492),
        .b(new_Jinkela_wire_598),
        .c(_197_)
    );

    or_bb _586_ (
        .a(_197_),
        .b(_196_),
        .c(_198_)
    );

    or_ii _587_ (
        .a(new_Jinkela_wire_103),
        .b(new_Jinkela_wire_1055),
        .c(_199_)
    );

    or_bi _588_ (
        .a(new_Jinkela_wire_462),
        .b(new_Jinkela_wire_875),
        .c(_200_)
    );

    and_bi _589_ (
        .a(new_Jinkela_wire_461),
        .b(new_Jinkela_wire_877),
        .c(_201_)
    );

    and_bi _590_ (
        .a(_200_),
        .b(_201_),
        .c(_202_)
    );

    and_bi _591_ (
        .a(new_Jinkela_wire_1330),
        .b(new_Jinkela_wire_1633),
        .c(_203_)
    );

    and_bi _592_ (
        .a(new_Jinkela_wire_1632),
        .b(new_Jinkela_wire_1329),
        .c(_204_)
    );

    or_bb _593_ (
        .a(_204_),
        .b(_203_),
        .c(_205_)
    );

    or_bb _594_ (
        .a(new_Jinkela_wire_1497),
        .b(new_Jinkela_wire_1545),
        .c(_206_)
    );

    and_bb _595_ (
        .a(new_Jinkela_wire_1496),
        .b(new_Jinkela_wire_1544),
        .c(_207_)
    );

    and_bi _596_ (
        .a(_206_),
        .b(_207_),
        .c(_208_)
    );

    or_bb _597_ (
        .a(new_Jinkela_wire_1378),
        .b(new_Jinkela_wire_1191),
        .c(_209_)
    );

    and_bi _598_ (
        .a(new_Jinkela_wire_1190),
        .b(new_Jinkela_wire_1679),
        .c(_210_)
    );

    and_bi _599_ (
        .a(_209_),
        .b(_210_),
        .c(_211_)
    );

    or_bi _600_ (
        .a(new_Jinkela_wire_1623),
        .b(new_Jinkela_wire_1704),
        .c(_212_)
    );

    bfr new_Jinkela_buffer_288 (
        .din(new_Jinkela_wire_373),
        .dout(new_Jinkela_wire_374)
    );

    bfr new_Jinkela_buffer_699 (
        .din(new_Jinkela_wire_904),
        .dout(new_Jinkela_wire_905)
    );

    and_bi _388_ (
        .a(new_Jinkela_wire_600),
        .b(new_Jinkela_wire_5),
        .c(_000_)
    );

    or_bi _389_ (
        .a(_000_),
        .b(_361_),
        .c(_001_)
    );

    bfr new_Jinkela_buffer_353 (
        .din(new_Jinkela_wire_457),
        .dout(new_Jinkela_wire_458)
    );

    bfr new_Jinkela_buffer_780 (
        .din(new_Jinkela_wire_1012),
        .dout(new_Jinkela_wire_1013)
    );

    bfr new_Jinkela_buffer_289 (
        .din(new_Jinkela_wire_374),
        .dout(new_Jinkela_wire_375)
    );

    spl2 new_Jinkela_splitter_77 (
        .a(new_Jinkela_wire_905),
        .b(new_Jinkela_wire_906),
        .c(new_Jinkela_wire_907)
    );

    or_bi _390_ (
        .a(new_Jinkela_wire_1641),
        .b(new_Jinkela_wire_1689),
        .c(_002_)
    );

    bfr new_Jinkela_buffer_304 (
        .din(new_Jinkela_wire_397),
        .dout(new_Jinkela_wire_398)
    );

    bfr new_Jinkela_buffer_732 (
        .din(new_Jinkela_wire_953),
        .dout(new_Jinkela_wire_954)
    );

    and_bi _391_ (
        .a(new_Jinkela_wire_1640),
        .b(new_Jinkela_wire_1688),
        .c(_003_)
    );

    bfr new_Jinkela_buffer_290 (
        .din(new_Jinkela_wire_375),
        .dout(new_Jinkela_wire_376)
    );

    bfr new_Jinkela_buffer_712 (
        .din(new_Jinkela_wire_925),
        .dout(new_Jinkela_wire_926)
    );

    and_bi _392_ (
        .a(_002_),
        .b(_003_),
        .c(_004_)
    );

    spl2 new_Jinkela_splitter_45 (
        .a(N21),
        .b(new_Jinkela_wire_525),
        .c(new_Jinkela_wire_527)
    );

    bfr new_Jinkela_buffer_713 (
        .din(new_Jinkela_wire_926),
        .dout(new_Jinkela_wire_927)
    );

    or_bb _393_ (
        .a(new_Jinkela_wire_1146),
        .b(new_Jinkela_wire_1676),
        .c(_005_)
    );

    bfr new_Jinkela_buffer_354 (
        .din(new_Jinkela_wire_463),
        .dout(new_Jinkela_wire_464)
    );

    bfr new_Jinkela_buffer_291 (
        .din(new_Jinkela_wire_376),
        .dout(new_Jinkela_wire_377)
    );

    and_bb _394_ (
        .a(new_Jinkela_wire_1145),
        .b(new_Jinkela_wire_1674),
        .c(_006_)
    );

    bfr new_Jinkela_buffer_781 (
        .din(new_Jinkela_wire_1018),
        .dout(new_Jinkela_wire_1019)
    );

    bfr new_Jinkela_buffer_305 (
        .din(new_Jinkela_wire_398),
        .dout(new_Jinkela_wire_399)
    );

    bfr new_Jinkela_buffer_714 (
        .din(new_Jinkela_wire_927),
        .dout(new_Jinkela_wire_928)
    );

    and_bi _395_ (
        .a(_005_),
        .b(_006_),
        .c(_007_)
    );

    bfr new_Jinkela_buffer_292 (
        .din(new_Jinkela_wire_377),
        .dout(new_Jinkela_wire_378)
    );

    bfr new_Jinkela_buffer_733 (
        .din(new_Jinkela_wire_954),
        .dout(new_Jinkela_wire_955)
    );

    or_bi _396_ (
        .a(new_Jinkela_wire_1529),
        .b(new_Jinkela_wire_1710),
        .c(_008_)
    );

    bfr new_Jinkela_buffer_328 (
        .din(new_Jinkela_wire_429),
        .dout(new_Jinkela_wire_430)
    );

    bfr new_Jinkela_buffer_715 (
        .din(new_Jinkela_wire_928),
        .dout(new_Jinkela_wire_929)
    );

    and_bi _397_ (
        .a(new_Jinkela_wire_1528),
        .b(new_Jinkela_wire_1709),
        .c(_009_)
    );

    bfr new_Jinkela_buffer_293 (
        .din(new_Jinkela_wire_378),
        .dout(new_Jinkela_wire_379)
    );

    bfr new_Jinkela_buffer_755 (
        .din(new_Jinkela_wire_984),
        .dout(new_Jinkela_wire_985)
    );

    and_bi _398_ (
        .a(new_Jinkela_wire_1232),
        .b(new_Jinkela_wire_1653),
        .c(_010_)
    );

    bfr new_Jinkela_buffer_306 (
        .din(new_Jinkela_wire_399),
        .dout(new_Jinkela_wire_400)
    );

    bfr new_Jinkela_buffer_716 (
        .din(new_Jinkela_wire_929),
        .dout(new_Jinkela_wire_930)
    );

    or_ii _399_ (
        .a(new_Jinkela_wire_421),
        .b(new_Jinkela_wire_1054),
        .c(_011_)
    );

    bfr new_Jinkela_buffer_294 (
        .din(new_Jinkela_wire_379),
        .dout(new_Jinkela_wire_380)
    );

    bfr new_Jinkela_buffer_734 (
        .din(new_Jinkela_wire_955),
        .dout(new_Jinkela_wire_956)
    );

    or_bi _400_ (
        .a(new_Jinkela_wire_944),
        .b(new_Jinkela_wire_664),
        .c(_012_)
    );

    bfr new_Jinkela_buffer_717 (
        .din(new_Jinkela_wire_930),
        .dout(new_Jinkela_wire_931)
    );

    and_bi _401_ (
        .a(new_Jinkela_wire_946),
        .b(new_Jinkela_wire_666),
        .c(_013_)
    );

    spl2 new_Jinkela_splitter_32 (
        .a(new_Jinkela_wire_380),
        .b(new_Jinkela_wire_381),
        .c(new_Jinkela_wire_382)
    );

    or_bi _402_ (
        .a(_013_),
        .b(_012_),
        .c(_014_)
    );

    bfr new_Jinkela_buffer_329 (
        .din(new_Jinkela_wire_430),
        .dout(new_Jinkela_wire_431)
    );

    bfr new_Jinkela_buffer_718 (
        .din(new_Jinkela_wire_931),
        .dout(new_Jinkela_wire_932)
    );

    or_bi _403_ (
        .a(new_Jinkela_wire_772),
        .b(new_Jinkela_wire_69),
        .c(_015_)
    );

    bfr new_Jinkela_buffer_307 (
        .din(new_Jinkela_wire_400),
        .dout(new_Jinkela_wire_401)
    );

    bfr new_Jinkela_buffer_735 (
        .din(new_Jinkela_wire_956),
        .dout(new_Jinkela_wire_957)
    );

    and_bi _404_ (
        .a(new_Jinkela_wire_774),
        .b(new_Jinkela_wire_73),
        .c(_016_)
    );

    bfr new_Jinkela_buffer_308 (
        .din(new_Jinkela_wire_401),
        .dout(new_Jinkela_wire_402)
    );

    bfr new_Jinkela_buffer_719 (
        .din(new_Jinkela_wire_932),
        .dout(new_Jinkela_wire_933)
    );

    or_bi _405_ (
        .a(_016_),
        .b(_015_),
        .c(_017_)
    );

    bfr new_Jinkela_buffer_756 (
        .din(new_Jinkela_wire_985),
        .dout(new_Jinkela_wire_986)
    );

    or_bi _406_ (
        .a(new_Jinkela_wire_1535),
        .b(new_Jinkela_wire_1522),
        .c(_018_)
    );

    bfr new_Jinkela_buffer_309 (
        .din(new_Jinkela_wire_402),
        .dout(new_Jinkela_wire_403)
    );

    bfr new_Jinkela_buffer_720 (
        .din(new_Jinkela_wire_933),
        .dout(new_Jinkela_wire_934)
    );

    and_bi _407_ (
        .a(new_Jinkela_wire_1534),
        .b(new_Jinkela_wire_1521),
        .c(_019_)
    );

    bfr new_Jinkela_buffer_330 (
        .din(new_Jinkela_wire_431),
        .dout(new_Jinkela_wire_432)
    );

    bfr new_Jinkela_buffer_736 (
        .din(new_Jinkela_wire_957),
        .dout(new_Jinkela_wire_958)
    );

    and_bi _411_ (
        .a(_021_),
        .b(_022_),
        .c(_023_)
    );

    bfr new_Jinkela_buffer_310 (
        .din(new_Jinkela_wire_403),
        .dout(new_Jinkela_wire_404)
    );

    bfr new_Jinkela_buffer_721 (
        .din(new_Jinkela_wire_934),
        .dout(new_Jinkela_wire_935)
    );

    or_bb _412_ (
        .a(new_Jinkela_wire_1015),
        .b(new_Jinkela_wire_980),
        .c(_024_)
    );

    spl4L new_Jinkela_splitter_43 (
        .a(new_Jinkela_wire_493),
        .d(new_Jinkela_wire_494),
        .e(new_Jinkela_wire_495),
        .b(new_Jinkela_wire_496),
        .c(new_Jinkela_wire_497)
    );

    and_bb _413_ (
        .a(new_Jinkela_wire_1013),
        .b(new_Jinkela_wire_978),
        .c(_025_)
    );

    spl2 new_Jinkela_splitter_93 (
        .a(N37),
        .b(new_Jinkela_wire_1057),
        .c(new_Jinkela_wire_1059)
    );

    bfr new_Jinkela_buffer_311 (
        .din(new_Jinkela_wire_404),
        .dout(new_Jinkela_wire_405)
    );

    bfr new_Jinkela_buffer_722 (
        .din(new_Jinkela_wire_935),
        .dout(new_Jinkela_wire_936)
    );

    and_bi _414_ (
        .a(_024_),
        .b(_025_),
        .c(_026_)
    );

    bfr new_Jinkela_buffer_331 (
        .din(new_Jinkela_wire_432),
        .dout(new_Jinkela_wire_433)
    );

    bfr new_Jinkela_buffer_737 (
        .din(new_Jinkela_wire_958),
        .dout(new_Jinkela_wire_959)
    );

    or_bi _415_ (
        .a(new_Jinkela_wire_737),
        .b(new_Jinkela_wire_282),
        .c(_027_)
    );

    bfr new_Jinkela_buffer_312 (
        .din(new_Jinkela_wire_405),
        .dout(new_Jinkela_wire_406)
    );

    bfr new_Jinkela_buffer_723 (
        .din(new_Jinkela_wire_936),
        .dout(new_Jinkela_wire_937)
    );

    and_bi _416_ (
        .a(new_Jinkela_wire_733),
        .b(new_Jinkela_wire_280),
        .c(_028_)
    );

    bfr new_Jinkela_buffer_757 (
        .din(new_Jinkela_wire_986),
        .dout(new_Jinkela_wire_987)
    );

    or_bi _417_ (
        .a(_028_),
        .b(_027_),
        .c(_029_)
    );

    bfr new_Jinkela_buffer_379 (
        .din(new_Jinkela_wire_491),
        .dout(new_Jinkela_wire_492)
    );

    bfr new_Jinkela_buffer_313 (
        .din(new_Jinkela_wire_406),
        .dout(new_Jinkela_wire_407)
    );

    bfr new_Jinkela_buffer_724 (
        .din(new_Jinkela_wire_937),
        .dout(new_Jinkela_wire_938)
    );

    or_bi _418_ (
        .a(new_Jinkela_wire_1406),
        .b(new_Jinkela_wire_1175),
        .c(_030_)
    );

    bfr new_Jinkela_buffer_332 (
        .din(new_Jinkela_wire_433),
        .dout(new_Jinkela_wire_434)
    );

    bfr new_Jinkela_buffer_738 (
        .din(new_Jinkela_wire_959),
        .dout(new_Jinkela_wire_960)
    );

    and_bi _419_ (
        .a(new_Jinkela_wire_1405),
        .b(new_Jinkela_wire_1174),
        .c(_031_)
    );

    bfr new_Jinkela_buffer_314 (
        .din(new_Jinkela_wire_407),
        .dout(new_Jinkela_wire_408)
    );

    bfr new_Jinkela_buffer_725 (
        .din(new_Jinkela_wire_938),
        .dout(new_Jinkela_wire_939)
    );

    and_bi _420_ (
        .a(_030_),
        .b(_031_),
        .c(_032_)
    );

    bfr new_Jinkela_buffer_355 (
        .din(new_Jinkela_wire_464),
        .dout(new_Jinkela_wire_465)
    );

    spl4L new_Jinkela_splitter_92 (
        .a(new_Jinkela_wire_1052),
        .d(new_Jinkela_wire_1053),
        .e(new_Jinkela_wire_1054),
        .b(new_Jinkela_wire_1055),
        .c(new_Jinkela_wire_1056)
    );

    or_bb _421_ (
        .a(new_Jinkela_wire_386),
        .b(new_Jinkela_wire_700),
        .c(_033_)
    );

    bfr new_Jinkela_buffer_315 (
        .din(new_Jinkela_wire_408),
        .dout(new_Jinkela_wire_409)
    );

    bfr new_Jinkela_buffer_726 (
        .din(new_Jinkela_wire_939),
        .dout(new_Jinkela_wire_940)
    );

    and_bb _422_ (
        .a(new_Jinkela_wire_387),
        .b(new_Jinkela_wire_701),
        .c(_034_)
    );

    bfr new_Jinkela_buffer_333 (
        .din(new_Jinkela_wire_434),
        .dout(new_Jinkela_wire_435)
    );

    bfr new_Jinkela_buffer_739 (
        .din(new_Jinkela_wire_960),
        .dout(new_Jinkela_wire_961)
    );

    and_bi _423_ (
        .a(_033_),
        .b(_034_),
        .c(_035_)
    );

    bfr new_Jinkela_buffer_316 (
        .din(new_Jinkela_wire_409),
        .dout(new_Jinkela_wire_410)
    );

    spl2 new_Jinkela_splitter_80 (
        .a(new_Jinkela_wire_940),
        .b(new_Jinkela_wire_941),
        .c(new_Jinkela_wire_942)
    );

    or_bi _424_ (
        .a(new_Jinkela_wire_1061),
        .b(new_Jinkela_wire_563),
        .c(_036_)
    );

    spl4L new_Jinkela_splitter_46 (
        .a(new_Jinkela_wire_527),
        .d(new_Jinkela_wire_528),
        .e(new_Jinkela_wire_529),
        .b(new_Jinkela_wire_530),
        .c(new_Jinkela_wire_531)
    );

    bfr new_Jinkela_buffer_740 (
        .din(new_Jinkela_wire_961),
        .dout(new_Jinkela_wire_962)
    );

    and_bi _425_ (
        .a(new_Jinkela_wire_1060),
        .b(new_Jinkela_wire_561),
        .c(_037_)
    );

    spl2 new_Jinkela_splitter_48 (
        .a(N33),
        .b(new_Jinkela_wire_560),
        .c(new_Jinkela_wire_562)
    );

    bfr new_Jinkela_buffer_317 (
        .din(new_Jinkela_wire_410),
        .dout(new_Jinkela_wire_411)
    );

    bfr new_Jinkela_buffer_758 (
        .din(new_Jinkela_wire_987),
        .dout(new_Jinkela_wire_988)
    );

    or_bi _426_ (
        .a(_037_),
        .b(_036_),
        .c(_038_)
    );

    bfr new_Jinkela_buffer_334 (
        .din(new_Jinkela_wire_435),
        .dout(new_Jinkela_wire_436)
    );

    spl4L new_Jinkela_splitter_94 (
        .a(new_Jinkela_wire_1059),
        .d(new_Jinkela_wire_1060),
        .e(new_Jinkela_wire_1061),
        .b(new_Jinkela_wire_1062),
        .c(new_Jinkela_wire_1063)
    );

    or_bi _427_ (
        .a(new_Jinkela_wire_1706),
        .b(new_Jinkela_wire_1288),
        .c(_039_)
    );

    spl4L new_Jinkela_splitter_91 (
        .a(new_Jinkela_wire_1047),
        .d(new_Jinkela_wire_1048),
        .e(new_Jinkela_wire_1049),
        .b(new_Jinkela_wire_1050),
        .c(new_Jinkela_wire_1051)
    );

    bfr new_Jinkela_buffer_318 (
        .din(new_Jinkela_wire_411),
        .dout(new_Jinkela_wire_412)
    );

    bfr new_Jinkela_buffer_741 (
        .din(new_Jinkela_wire_962),
        .dout(new_Jinkela_wire_963)
    );

    and_bi _428_ (
        .a(new_Jinkela_wire_1705),
        .b(new_Jinkela_wire_1287),
        .c(_040_)
    );

    bfr new_Jinkela_buffer_356 (
        .din(new_Jinkela_wire_465),
        .dout(new_Jinkela_wire_466)
    );

    bfr new_Jinkela_buffer_759 (
        .din(new_Jinkela_wire_988),
        .dout(new_Jinkela_wire_989)
    );

    and_bi _429_ (
        .a(_039_),
        .b(_040_),
        .c(_041_)
    );

    bfr new_Jinkela_buffer_319 (
        .din(new_Jinkela_wire_412),
        .dout(new_Jinkela_wire_413)
    );

    bfr new_Jinkela_buffer_742 (
        .din(new_Jinkela_wire_963),
        .dout(new_Jinkela_wire_964)
    );

    or_bb _430_ (
        .a(new_Jinkela_wire_1188),
        .b(new_Jinkela_wire_1590),
        .c(_042_)
    );

    bfr new_Jinkela_buffer_335 (
        .din(new_Jinkela_wire_436),
        .dout(new_Jinkela_wire_437)
    );

    bfr new_Jinkela_buffer_782 (
        .din(new_Jinkela_wire_1019),
        .dout(new_Jinkela_wire_1020)
    );

    and_bb _431_ (
        .a(new_Jinkela_wire_1187),
        .b(new_Jinkela_wire_1587),
        .c(_043_)
    );

    bfr new_Jinkela_buffer_320 (
        .din(new_Jinkela_wire_413),
        .dout(new_Jinkela_wire_414)
    );

    bfr new_Jinkela_buffer_743 (
        .din(new_Jinkela_wire_964),
        .dout(new_Jinkela_wire_965)
    );

    and_bi _432_ (
        .a(_042_),
        .b(_043_),
        .c(_044_)
    );

    bfr new_Jinkela_buffer_0 (
        .din(new_Jinkela_wire_0),
        .dout(new_Jinkela_wire_1)
    );

    spl2 new_Jinkela_splitter_0 (
        .a(N97),
        .b(new_Jinkela_wire_0),
        .c(new_Jinkela_wire_2)
    );

    spl2 new_Jinkela_splitter_6 (
        .a(N73),
        .b(new_Jinkela_wire_68),
        .c(new_Jinkela_wire_70)
    );

    spl2 new_Jinkela_splitter_3 (
        .a(N113),
        .b(new_Jinkela_wire_34),
        .c(new_Jinkela_wire_36)
    );

    spl4L new_Jinkela_splitter_1 (
        .a(new_Jinkela_wire_2),
        .d(new_Jinkela_wire_3),
        .e(new_Jinkela_wire_4),
        .b(new_Jinkela_wire_5),
        .c(new_Jinkela_wire_6)
    );

    spl4L new_Jinkela_splitter_4 (
        .a(new_Jinkela_wire_36),
        .d(new_Jinkela_wire_37),
        .e(new_Jinkela_wire_38),
        .b(new_Jinkela_wire_39),
        .c(new_Jinkela_wire_40)
    );

    bfr new_Jinkela_buffer_893 (
        .din(new_Jinkela_wire_1210),
        .dout(new_Jinkela_wire_1211)
    );

    bfr new_Jinkela_buffer_510 (
        .din(new_Jinkela_wire_659),
        .dout(new_Jinkela_wire_660)
    );

    bfr new_Jinkela_buffer_887 (
        .din(new_Jinkela_wire_1198),
        .dout(new_Jinkela_wire_1199)
    );

    or_bi _409_ (
        .a(new_Jinkela_wire_1586),
        .b(new_Jinkela_wire_1140),
        .c(_021_)
    );

    spl2 new_Jinkela_splitter_66 (
        .a(N89),
        .b(new_Jinkela_wire_771),
        .c(new_Jinkela_wire_773)
    );

    spl2 new_Jinkela_splitter_56 (
        .a(new_Jinkela_wire_660),
        .b(new_Jinkela_wire_661),
        .c(new_Jinkela_wire_662)
    );

    bfr new_Jinkela_buffer_888 (
        .din(new_Jinkela_wire_1199),
        .dout(new_Jinkela_wire_1200)
    );

    bfr new_Jinkela_buffer_542 (
        .din(new_Jinkela_wire_707),
        .dout(new_Jinkela_wire_708)
    );

    bfr new_Jinkela_buffer_897 (
        .din(new_Jinkela_wire_1216),
        .dout(new_Jinkela_wire_1217)
    );

    bfr new_Jinkela_buffer_894 (
        .din(new_Jinkela_wire_1211),
        .dout(new_Jinkela_wire_1212)
    );

    bfr new_Jinkela_buffer_523 (
        .din(new_Jinkela_wire_680),
        .dout(new_Jinkela_wire_681)
    );

    bfr new_Jinkela_buffer_889 (
        .din(new_Jinkela_wire_1200),
        .dout(new_Jinkela_wire_1201)
    );

    bfr new_Jinkela_buffer_524 (
        .din(new_Jinkela_wire_681),
        .dout(new_Jinkela_wire_682)
    );

    spl2 new_Jinkela_splitter_69 (
        .a(N125),
        .b(new_Jinkela_wire_805),
        .c(new_Jinkela_wire_807)
    );

    bfr new_Jinkela_buffer_594 (
        .din(new_Jinkela_wire_769),
        .dout(new_Jinkela_wire_770)
    );

    bfr new_Jinkela_buffer_890 (
        .din(new_Jinkela_wire_1201),
        .dout(new_Jinkela_wire_1202)
    );

    bfr new_Jinkela_buffer_525 (
        .din(new_Jinkela_wire_682),
        .dout(new_Jinkela_wire_683)
    );

    bfr new_Jinkela_buffer_895 (
        .din(new_Jinkela_wire_1212),
        .dout(new_Jinkela_wire_1213)
    );

    bfr new_Jinkela_buffer_543 (
        .din(new_Jinkela_wire_708),
        .dout(new_Jinkela_wire_709)
    );

    spl4L new_Jinkela_splitter_120 (
        .a(new_Jinkela_wire_1202),
        .d(new_Jinkela_wire_1203),
        .e(new_Jinkela_wire_1204),
        .b(new_Jinkela_wire_1205),
        .c(new_Jinkela_wire_1206)
    );

    bfr new_Jinkela_buffer_526 (
        .din(new_Jinkela_wire_683),
        .dout(new_Jinkela_wire_684)
    );

    bfr new_Jinkela_buffer_907 (
        .din(_116_),
        .dout(new_Jinkela_wire_1235)
    );

    bfr new_Jinkela_buffer_566 (
        .din(new_Jinkela_wire_739),
        .dout(new_Jinkela_wire_740)
    );

    bfr new_Jinkela_buffer_527 (
        .din(new_Jinkela_wire_684),
        .dout(new_Jinkela_wire_685)
    );

    bfr new_Jinkela_buffer_898 (
        .din(new_Jinkela_wire_1217),
        .dout(new_Jinkela_wire_1218)
    );

    bfr new_Jinkela_buffer_544 (
        .din(new_Jinkela_wire_709),
        .dout(new_Jinkela_wire_710)
    );

    bfr new_Jinkela_buffer_528 (
        .din(new_Jinkela_wire_685),
        .dout(new_Jinkela_wire_686)
    );

    spl4L new_Jinkela_splitter_129 (
        .a(new_Jinkela_wire_1257),
        .d(new_Jinkela_wire_1258),
        .e(new_Jinkela_wire_1259),
        .b(new_Jinkela_wire_1260),
        .c(new_Jinkela_wire_1261)
    );

    bfr new_Jinkela_buffer_595 (
        .din(new_Jinkela_wire_771),
        .dout(new_Jinkela_wire_772)
    );

    bfr new_Jinkela_buffer_899 (
        .din(new_Jinkela_wire_1218),
        .dout(new_Jinkela_wire_1219)
    );

    spl2 new_Jinkela_splitter_128 (
        .a(_243_),
        .b(new_Jinkela_wire_1255),
        .c(new_Jinkela_wire_1256)
    );

    bfr new_Jinkela_buffer_529 (
        .din(new_Jinkela_wire_686),
        .dout(new_Jinkela_wire_687)
    );

    bfr new_Jinkela_buffer_900 (
        .din(new_Jinkela_wire_1219),
        .dout(new_Jinkela_wire_1220)
    );

    bfr new_Jinkela_buffer_545 (
        .din(new_Jinkela_wire_710),
        .dout(new_Jinkela_wire_711)
    );

    spl4L new_Jinkela_splitter_126 (
        .a(new_Jinkela_wire_1235),
        .d(new_Jinkela_wire_1236),
        .e(new_Jinkela_wire_1237),
        .b(new_Jinkela_wire_1238),
        .c(new_Jinkela_wire_1239)
    );

    spl2 new_Jinkela_splitter_131 (
        .a(_263_),
        .b(new_Jinkela_wire_1276),
        .c(new_Jinkela_wire_1277)
    );

    bfr new_Jinkela_buffer_530 (
        .din(new_Jinkela_wire_687),
        .dout(new_Jinkela_wire_688)
    );

    bfr new_Jinkela_buffer_901 (
        .din(new_Jinkela_wire_1220),
        .dout(new_Jinkela_wire_1221)
    );

    bfr new_Jinkela_buffer_567 (
        .din(new_Jinkela_wire_740),
        .dout(new_Jinkela_wire_741)
    );

    bfr new_Jinkela_buffer_920 (
        .din(new_Jinkela_wire_1261),
        .dout(new_Jinkela_wire_1262)
    );

    bfr new_Jinkela_buffer_531 (
        .din(new_Jinkela_wire_688),
        .dout(new_Jinkela_wire_689)
    );

    bfr new_Jinkela_buffer_902 (
        .din(new_Jinkela_wire_1221),
        .dout(new_Jinkela_wire_1222)
    );

    bfr new_Jinkela_buffer_546 (
        .din(new_Jinkela_wire_711),
        .dout(new_Jinkela_wire_712)
    );

    spl2 new_Jinkela_splitter_133 (
        .a(_076_),
        .b(new_Jinkela_wire_1280),
        .c(new_Jinkela_wire_1281)
    );

    bfr new_Jinkela_buffer_532 (
        .din(new_Jinkela_wire_689),
        .dout(new_Jinkela_wire_690)
    );

    spl2 new_Jinkela_splitter_132 (
        .a(_138_),
        .b(new_Jinkela_wire_1278),
        .c(new_Jinkela_wire_1279)
    );

    bfr new_Jinkela_buffer_903 (
        .din(new_Jinkela_wire_1222),
        .dout(new_Jinkela_wire_1223)
    );

    spl2 new_Jinkela_splitter_72 (
        .a(N53),
        .b(new_Jinkela_wire_839),
        .c(new_Jinkela_wire_841)
    );

    bfr new_Jinkela_buffer_909 (
        .din(new_Jinkela_wire_1240),
        .dout(new_Jinkela_wire_1241)
    );

    bfr new_Jinkela_buffer_533 (
        .din(new_Jinkela_wire_690),
        .dout(new_Jinkela_wire_691)
    );

    bfr new_Jinkela_buffer_904 (
        .din(new_Jinkela_wire_1223),
        .dout(new_Jinkela_wire_1224)
    );

    bfr new_Jinkela_buffer_547 (
        .din(new_Jinkela_wire_712),
        .dout(new_Jinkela_wire_713)
    );

    bfr new_Jinkela_buffer_534 (
        .din(new_Jinkela_wire_691),
        .dout(new_Jinkela_wire_692)
    );

    bfr new_Jinkela_buffer_905 (
        .din(new_Jinkela_wire_1224),
        .dout(new_Jinkela_wire_1225)
    );

    bfr new_Jinkela_buffer_568 (
        .din(new_Jinkela_wire_741),
        .dout(new_Jinkela_wire_742)
    );

    bfr new_Jinkela_buffer_910 (
        .din(new_Jinkela_wire_1241),
        .dout(new_Jinkela_wire_1242)
    );

    bfr new_Jinkela_buffer_535 (
        .din(new_Jinkela_wire_692),
        .dout(new_Jinkela_wire_693)
    );

    spl4L new_Jinkela_splitter_123 (
        .a(new_Jinkela_wire_1225),
        .d(new_Jinkela_wire_1226),
        .e(new_Jinkela_wire_1227),
        .b(new_Jinkela_wire_1228),
        .c(new_Jinkela_wire_1229)
    );

    bfr new_Jinkela_buffer_548 (
        .din(new_Jinkela_wire_713),
        .dout(new_Jinkela_wire_714)
    );

    bfr new_Jinkela_buffer_919 (
        .din(_047_),
        .dout(new_Jinkela_wire_1257)
    );

    bfr new_Jinkela_buffer_536 (
        .din(new_Jinkela_wire_693),
        .dout(new_Jinkela_wire_694)
    );

    spl4L new_Jinkela_splitter_67 (
        .a(new_Jinkela_wire_773),
        .d(new_Jinkela_wire_774),
        .e(new_Jinkela_wire_775),
        .b(new_Jinkela_wire_776),
        .c(new_Jinkela_wire_777)
    );

    spl2 new_Jinkela_splitter_59 (
        .a(new_Jinkela_wire_694),
        .b(new_Jinkela_wire_695),
        .c(new_Jinkela_wire_696)
    );

    bfr new_Jinkela_buffer_911 (
        .din(new_Jinkela_wire_1242),
        .dout(new_Jinkela_wire_1243)
    );

    bfr new_Jinkela_buffer_569 (
        .din(new_Jinkela_wire_742),
        .dout(new_Jinkela_wire_743)
    );

    bfr new_Jinkela_buffer_908 (
        .din(new_Jinkela_wire_1239),
        .dout(new_Jinkela_wire_1240)
    );

    bfr new_Jinkela_buffer_912 (
        .din(new_Jinkela_wire_1243),
        .dout(new_Jinkela_wire_1244)
    );

    bfr new_Jinkela_buffer_549 (
        .din(new_Jinkela_wire_714),
        .dout(new_Jinkela_wire_715)
    );

    bfr new_Jinkela_buffer_921 (
        .din(new_Jinkela_wire_1262),
        .dout(new_Jinkela_wire_1263)
    );

    bfr new_Jinkela_buffer_550 (
        .din(new_Jinkela_wire_715),
        .dout(new_Jinkela_wire_716)
    );

    bfr new_Jinkela_buffer_913 (
        .din(new_Jinkela_wire_1244),
        .dout(new_Jinkela_wire_1245)
    );

    spl4L new_Jinkela_splitter_70 (
        .a(new_Jinkela_wire_807),
        .d(new_Jinkela_wire_808),
        .e(new_Jinkela_wire_809),
        .b(new_Jinkela_wire_810),
        .c(new_Jinkela_wire_811)
    );

    spl2 new_Jinkela_splitter_134 (
        .a(_312_),
        .b(new_Jinkela_wire_1282),
        .c(new_Jinkela_wire_1283)
    );

    bfr new_Jinkela_buffer_551 (
        .din(new_Jinkela_wire_716),
        .dout(new_Jinkela_wire_717)
    );

    spl2 new_Jinkela_splitter_136 (
        .a(_038_),
        .b(new_Jinkela_wire_1287),
        .c(new_Jinkela_wire_1288)
    );

    bfr new_Jinkela_buffer_914 (
        .din(new_Jinkela_wire_1245),
        .dout(new_Jinkela_wire_1246)
    );

    bfr new_Jinkela_buffer_570 (
        .din(new_Jinkela_wire_743),
        .dout(new_Jinkela_wire_744)
    );

    bfr new_Jinkela_buffer_922 (
        .din(new_Jinkela_wire_1263),
        .dout(new_Jinkela_wire_1264)
    );

    bfr new_Jinkela_buffer_552 (
        .din(new_Jinkela_wire_717),
        .dout(new_Jinkela_wire_718)
    );

    bfr new_Jinkela_buffer_915 (
        .din(new_Jinkela_wire_1246),
        .dout(new_Jinkela_wire_1247)
    );

    bfr new_Jinkela_buffer_553 (
        .din(new_Jinkela_wire_718),
        .dout(new_Jinkela_wire_719)
    );

    bfr new_Jinkela_buffer_916 (
        .din(new_Jinkela_wire_1247),
        .dout(new_Jinkela_wire_1248)
    );

    bfr new_Jinkela_buffer_571 (
        .din(new_Jinkela_wire_744),
        .dout(new_Jinkela_wire_745)
    );

    bfr new_Jinkela_buffer_930 (
        .din(_120_),
        .dout(new_Jinkela_wire_1284)
    );

    bfr new_Jinkela_buffer_99 (
        .din(new_Jinkela_wire_128),
        .dout(new_Jinkela_wire_129)
    );

    bfr new_Jinkela_buffer_136 (
        .din(new_Jinkela_wire_181),
        .dout(new_Jinkela_wire_182)
    );

    bfr new_Jinkela_buffer_100 (
        .din(new_Jinkela_wire_129),
        .dout(new_Jinkela_wire_130)
    );

    bfr new_Jinkela_buffer_116 (
        .din(new_Jinkela_wire_153),
        .dout(new_Jinkela_wire_154)
    );

    bfr new_Jinkela_buffer_101 (
        .din(new_Jinkela_wire_130),
        .dout(new_Jinkela_wire_131)
    );

    bfr new_Jinkela_buffer_192 (
        .din(new_Jinkela_wire_253),
        .dout(new_Jinkela_wire_254)
    );

    bfr new_Jinkela_buffer_102 (
        .din(new_Jinkela_wire_131),
        .dout(new_Jinkela_wire_132)
    );

    bfr new_Jinkela_buffer_117 (
        .din(new_Jinkela_wire_154),
        .dout(new_Jinkela_wire_155)
    );

    bfr new_Jinkela_buffer_103 (
        .din(new_Jinkela_wire_132),
        .dout(new_Jinkela_wire_133)
    );

    bfr new_Jinkela_buffer_137 (
        .din(new_Jinkela_wire_182),
        .dout(new_Jinkela_wire_183)
    );

    bfr new_Jinkela_buffer_104 (
        .din(new_Jinkela_wire_133),
        .dout(new_Jinkela_wire_134)
    );

    bfr new_Jinkela_buffer_118 (
        .din(new_Jinkela_wire_155),
        .dout(new_Jinkela_wire_156)
    );

    bfr new_Jinkela_buffer_105 (
        .din(new_Jinkela_wire_134),
        .dout(new_Jinkela_wire_135)
    );

    bfr new_Jinkela_buffer_161 (
        .din(new_Jinkela_wire_214),
        .dout(new_Jinkela_wire_215)
    );

    bfr new_Jinkela_buffer_106 (
        .din(new_Jinkela_wire_135),
        .dout(new_Jinkela_wire_136)
    );

    bfr new_Jinkela_buffer_119 (
        .din(new_Jinkela_wire_156),
        .dout(new_Jinkela_wire_157)
    );

    spl2 new_Jinkela_splitter_11 (
        .a(new_Jinkela_wire_136),
        .b(new_Jinkela_wire_137),
        .c(new_Jinkela_wire_138)
    );

    bfr new_Jinkela_buffer_120 (
        .din(new_Jinkela_wire_157),
        .dout(new_Jinkela_wire_158)
    );

    bfr new_Jinkela_buffer_138 (
        .din(new_Jinkela_wire_183),
        .dout(new_Jinkela_wire_184)
    );

    spl2 new_Jinkela_splitter_30 (
        .a(N109),
        .b(new_Jinkela_wire_349),
        .c(new_Jinkela_wire_351)
    );

    bfr new_Jinkela_buffer_193 (
        .din(new_Jinkela_wire_254),
        .dout(new_Jinkela_wire_255)
    );

    bfr new_Jinkela_buffer_121 (
        .din(new_Jinkela_wire_158),
        .dout(new_Jinkela_wire_159)
    );

    bfr new_Jinkela_buffer_139 (
        .din(new_Jinkela_wire_184),
        .dout(new_Jinkela_wire_185)
    );

    bfr new_Jinkela_buffer_122 (
        .din(new_Jinkela_wire_159),
        .dout(new_Jinkela_wire_160)
    );

    bfr new_Jinkela_buffer_162 (
        .din(new_Jinkela_wire_215),
        .dout(new_Jinkela_wire_216)
    );

    bfr new_Jinkela_buffer_123 (
        .din(new_Jinkela_wire_160),
        .dout(new_Jinkela_wire_161)
    );

    bfr new_Jinkela_buffer_140 (
        .din(new_Jinkela_wire_185),
        .dout(new_Jinkela_wire_186)
    );

    bfr new_Jinkela_buffer_124 (
        .din(new_Jinkela_wire_161),
        .dout(new_Jinkela_wire_162)
    );

    bfr new_Jinkela_buffer_125 (
        .din(new_Jinkela_wire_162),
        .dout(new_Jinkela_wire_163)
    );

    bfr new_Jinkela_buffer_141 (
        .din(new_Jinkela_wire_186),
        .dout(new_Jinkela_wire_187)
    );

    bfr new_Jinkela_buffer_126 (
        .din(new_Jinkela_wire_163),
        .dout(new_Jinkela_wire_164)
    );

    bfr new_Jinkela_buffer_163 (
        .din(new_Jinkela_wire_216),
        .dout(new_Jinkela_wire_217)
    );

    bfr new_Jinkela_buffer_127 (
        .din(new_Jinkela_wire_164),
        .dout(new_Jinkela_wire_165)
    );

    bfr new_Jinkela_buffer_142 (
        .din(new_Jinkela_wire_187),
        .dout(new_Jinkela_wire_188)
    );

    bfr new_Jinkela_buffer_128 (
        .din(new_Jinkela_wire_165),
        .dout(new_Jinkela_wire_166)
    );

    bfr new_Jinkela_buffer_215 (
        .din(new_Jinkela_wire_284),
        .dout(new_Jinkela_wire_285)
    );

    bfr new_Jinkela_buffer_129 (
        .din(new_Jinkela_wire_166),
        .dout(new_Jinkela_wire_167)
    );

    bfr new_Jinkela_buffer_143 (
        .din(new_Jinkela_wire_188),
        .dout(new_Jinkela_wire_189)
    );

    bfr new_Jinkela_buffer_130 (
        .din(new_Jinkela_wire_167),
        .dout(new_Jinkela_wire_168)
    );

    bfr new_Jinkela_buffer_164 (
        .din(new_Jinkela_wire_217),
        .dout(new_Jinkela_wire_218)
    );

    bfr new_Jinkela_buffer_131 (
        .din(new_Jinkela_wire_168),
        .dout(new_Jinkela_wire_169)
    );

    bfr new_Jinkela_buffer_144 (
        .din(new_Jinkela_wire_189),
        .dout(new_Jinkela_wire_190)
    );

    and_bi _601_ (
        .a(new_Jinkela_wire_1622),
        .b(new_Jinkela_wire_1703),
        .c(_213_)
    );

    bfr new_Jinkela_buffer_321 (
        .din(new_Jinkela_wire_414),
        .dout(new_Jinkela_wire_415)
    );

    or_bi _602_ (
        .a(new_Jinkela_wire_1539),
        .b(new_Jinkela_wire_1655),
        .c(_214_)
    );

    bfr new_Jinkela_buffer_336 (
        .din(new_Jinkela_wire_437),
        .dout(new_Jinkela_wire_438)
    );

    or_bb _603_ (
        .a(new_Jinkela_wire_1290),
        .b(new_Jinkela_wire_1215),
        .c(_215_)
    );

    spl2 new_Jinkela_splitter_35 (
        .a(new_Jinkela_wire_415),
        .b(new_Jinkela_wire_416),
        .c(new_Jinkela_wire_417)
    );

    or_bb _604_ (
        .a(new_Jinkela_wire_1650),
        .b(new_Jinkela_wire_1708),
        .c(_216_)
    );

    bfr new_Jinkela_buffer_337 (
        .din(new_Jinkela_wire_438),
        .dout(new_Jinkela_wire_439)
    );

    or_bb _605_ (
        .a(new_Jinkela_wire_1531),
        .b(new_Jinkela_wire_1186),
        .c(_217_)
    );

    bfr new_Jinkela_buffer_357 (
        .din(new_Jinkela_wire_466),
        .dout(new_Jinkela_wire_467)
    );

    or_bb _606_ (
        .a(new_Jinkela_wire_1164),
        .b(new_Jinkela_wire_1608),
        .c(_218_)
    );

    bfr new_Jinkela_buffer_380 (
        .din(new_Jinkela_wire_497),
        .dout(new_Jinkela_wire_498)
    );

    and_bi _607_ (
        .a(new_Jinkela_wire_1011),
        .b(new_Jinkela_wire_1643),
        .c(_219_)
    );

    bfr new_Jinkela_buffer_405 (
        .din(new_Jinkela_wire_525),
        .dout(new_Jinkela_wire_526)
    );

    bfr new_Jinkela_buffer_338 (
        .din(new_Jinkela_wire_439),
        .dout(new_Jinkela_wire_440)
    );

    and_bi _608_ (
        .a(new_Jinkela_wire_1642),
        .b(new_Jinkela_wire_1010),
        .c(_220_)
    );

    bfr new_Jinkela_buffer_358 (
        .din(new_Jinkela_wire_467),
        .dout(new_Jinkela_wire_468)
    );

    and_ii _609_ (
        .a(_220_),
        .b(_219_),
        .c(N726)
    );

    bfr new_Jinkela_buffer_339 (
        .din(new_Jinkela_wire_440),
        .dout(new_Jinkela_wire_441)
    );

    or_bi _610_ (
        .a(new_Jinkela_wire_1162),
        .b(new_Jinkela_wire_1251),
        .c(_221_)
    );

    spl2 new_Jinkela_splitter_51 (
        .a(N101),
        .b(new_Jinkela_wire_595),
        .c(new_Jinkela_wire_597)
    );

    and_bi _611_ (
        .a(new_Jinkela_wire_1702),
        .b(new_Jinkela_wire_311),
        .c(_222_)
    );

    bfr new_Jinkela_buffer_406 (
        .din(new_Jinkela_wire_531),
        .dout(new_Jinkela_wire_532)
    );

    bfr new_Jinkela_buffer_340 (
        .din(new_Jinkela_wire_441),
        .dout(new_Jinkela_wire_442)
    );

    and_bi _612_ (
        .a(new_Jinkela_wire_310),
        .b(new_Jinkela_wire_1701),
        .c(_223_)
    );

    bfr new_Jinkela_buffer_359 (
        .din(new_Jinkela_wire_468),
        .dout(new_Jinkela_wire_469)
    );

    and_ii _613_ (
        .a(_223_),
        .b(_222_),
        .c(N724)
    );

    bfr new_Jinkela_buffer_341 (
        .din(new_Jinkela_wire_442),
        .dout(new_Jinkela_wire_443)
    );

    and_bi _614_ (
        .a(new_Jinkela_wire_1451),
        .b(new_Jinkela_wire_1258),
        .c(_224_)
    );

    bfr new_Jinkela_buffer_381 (
        .din(new_Jinkela_wire_498),
        .dout(new_Jinkela_wire_499)
    );

    inv _615_ (
        .din(new_Jinkela_wire_1413),
        .dout(_225_)
    );

    bfr new_Jinkela_buffer_342 (
        .din(new_Jinkela_wire_443),
        .dout(new_Jinkela_wire_444)
    );

    or_bb _616_ (
        .a(new_Jinkela_wire_1553),
        .b(new_Jinkela_wire_1530),
        .c(_226_)
    );

    bfr new_Jinkela_buffer_360 (
        .din(new_Jinkela_wire_469),
        .dout(new_Jinkela_wire_470)
    );

    or_bi _617_ (
        .a(new_Jinkela_wire_1426),
        .b(new_Jinkela_wire_1254),
        .c(_227_)
    );

    bfr new_Jinkela_buffer_343 (
        .din(new_Jinkela_wire_444),
        .dout(new_Jinkela_wire_445)
    );

    and_bi _618_ (
        .a(new_Jinkela_wire_1557),
        .b(new_Jinkela_wire_206),
        .c(_228_)
    );

    and_bi _619_ (
        .a(new_Jinkela_wire_207),
        .b(new_Jinkela_wire_1556),
        .c(_229_)
    );

    bfr new_Jinkela_buffer_344 (
        .din(new_Jinkela_wire_445),
        .dout(new_Jinkela_wire_446)
    );

    and_ii _620_ (
        .a(_229_),
        .b(_228_),
        .c(N728)
    );

    bfr new_Jinkela_buffer_361 (
        .din(new_Jinkela_wire_470),
        .dout(new_Jinkela_wire_471)
    );

    or_bi _621_ (
        .a(new_Jinkela_wire_1163),
        .b(new_Jinkela_wire_1364),
        .c(_230_)
    );

    bfr new_Jinkela_buffer_345 (
        .din(new_Jinkela_wire_446),
        .dout(new_Jinkela_wire_447)
    );

    and_bi _622_ (
        .a(new_Jinkela_wire_1234),
        .b(new_Jinkela_wire_765),
        .c(_231_)
    );

    bfr new_Jinkela_buffer_382 (
        .din(new_Jinkela_wire_499),
        .dout(new_Jinkela_wire_500)
    );

    and_bi _623_ (
        .a(new_Jinkela_wire_766),
        .b(new_Jinkela_wire_1233),
        .c(_232_)
    );

    bfr new_Jinkela_buffer_346 (
        .din(new_Jinkela_wire_447),
        .dout(new_Jinkela_wire_448)
    );

    and_ii _624_ (
        .a(_232_),
        .b(_231_),
        .c(N725)
    );

    bfr new_Jinkela_buffer_362 (
        .din(new_Jinkela_wire_471),
        .dout(new_Jinkela_wire_472)
    );

    or_bi _625_ (
        .a(new_Jinkela_wire_1512),
        .b(new_Jinkela_wire_1297),
        .c(_233_)
    );

    bfr new_Jinkela_buffer_347 (
        .din(new_Jinkela_wire_448),
        .dout(new_Jinkela_wire_449)
    );

    and_bi _626_ (
        .a(new_Jinkela_wire_1654),
        .b(new_Jinkela_wire_1538),
        .c(_234_)
    );

    or_bb _627_ (
        .a(new_Jinkela_wire_1192),
        .b(new_Jinkela_wire_1367),
        .c(_235_)
    );

    bfr new_Jinkela_buffer_348 (
        .din(new_Jinkela_wire_449),
        .dout(new_Jinkela_wire_450)
    );

    and_bb _628_ (
        .a(new_Jinkela_wire_1565),
        .b(new_Jinkela_wire_1644),
        .c(_236_)
    );

    bfr new_Jinkela_buffer_363 (
        .din(new_Jinkela_wire_472),
        .dout(new_Jinkela_wire_473)
    );

    or_bb _629_ (
        .a(new_Jinkela_wire_1450),
        .b(new_Jinkela_wire_1259),
        .c(_237_)
    );

    bfr new_Jinkela_buffer_349 (
        .din(new_Jinkela_wire_450),
        .dout(new_Jinkela_wire_451)
    );

    or_bb _630_ (
        .a(new_Jinkela_wire_1527),
        .b(_236_),
        .c(_238_)
    );

    bfr new_Jinkela_buffer_383 (
        .din(new_Jinkela_wire_500),
        .dout(new_Jinkela_wire_501)
    );

    or_bb _631_ (
        .a(new_Jinkela_wire_1412),
        .b(new_Jinkela_wire_1611),
        .c(_239_)
    );

    bfr new_Jinkela_buffer_350 (
        .din(new_Jinkela_wire_451),
        .dout(new_Jinkela_wire_452)
    );

    or_bb _632_ (
        .a(new_Jinkela_wire_1289),
        .b(new_Jinkela_wire_1366),
        .c(_240_)
    );

    bfr new_Jinkela_buffer_364 (
        .din(new_Jinkela_wire_473),
        .dout(new_Jinkela_wire_474)
    );

    and_bi _633_ (
        .a(_239_),
        .b(new_Jinkela_wire_1136),
        .c(_241_)
    );

    bfr new_Jinkela_buffer_351 (
        .din(new_Jinkela_wire_452),
        .dout(new_Jinkela_wire_453)
    );

    and_bi _634_ (
        .a(_238_),
        .b(new_Jinkela_wire_1394),
        .c(_242_)
    );

    spl4L new_Jinkela_splitter_49 (
        .a(new_Jinkela_wire_562),
        .d(new_Jinkela_wire_563),
        .e(new_Jinkela_wire_564),
        .b(new_Jinkela_wire_565),
        .c(new_Jinkela_wire_566)
    );

    or_bb _635_ (
        .a(new_Jinkela_wire_1555),
        .b(new_Jinkela_wire_1509),
        .c(_243_)
    );

    spl4L new_Jinkela_splitter_52 (
        .a(new_Jinkela_wire_597),
        .d(new_Jinkela_wire_598),
        .e(new_Jinkela_wire_599),
        .b(new_Jinkela_wire_600),
        .c(new_Jinkela_wire_601)
    );

    bfr new_Jinkela_buffer_352 (
        .din(new_Jinkela_wire_453),
        .dout(new_Jinkela_wire_454)
    );

    or_bb _636_ (
        .a(new_Jinkela_wire_1256),
        .b(new_Jinkela_wire_1580),
        .c(_244_)
    );

    bfr new_Jinkela_buffer_365 (
        .din(new_Jinkela_wire_474),
        .dout(new_Jinkela_wire_475)
    );

    or_bi _637_ (
        .a(new_Jinkela_wire_1393),
        .b(new_Jinkela_wire_1467),
        .c(_245_)
    );

    spl2 new_Jinkela_splitter_38 (
        .a(new_Jinkela_wire_454),
        .b(new_Jinkela_wire_455),
        .c(new_Jinkela_wire_456)
    );

    and_bi _638_ (
        .a(new_Jinkela_wire_172),
        .b(new_Jinkela_wire_1294),
        .c(_246_)
    );

    bfr new_Jinkela_buffer_366 (
        .din(new_Jinkela_wire_475),
        .dout(new_Jinkela_wire_476)
    );

    and_bi _639_ (
        .a(new_Jinkela_wire_1293),
        .b(new_Jinkela_wire_171),
        .c(_247_)
    );

    bfr new_Jinkela_buffer_384 (
        .din(new_Jinkela_wire_501),
        .dout(new_Jinkela_wire_502)
    );

    and_ii _640_ (
        .a(_247_),
        .b(_246_),
        .c(new_net_709)
    );

    or_bi _641_ (
        .a(new_Jinkela_wire_1554),
        .b(new_Jinkela_wire_1484),
        .c(_248_)
    );

    bfr new_Jinkela_buffer_432 (
        .din(new_Jinkela_wire_560),
        .dout(new_Jinkela_wire_561)
    );

    bfr new_Jinkela_buffer_367 (
        .din(new_Jinkela_wire_476),
        .dout(new_Jinkela_wire_477)
    );

    or_bb _642_ (
        .a(new_Jinkela_wire_1664),
        .b(new_Jinkela_wire_1564),
        .c(_249_)
    );

    bfr new_Jinkela_buffer_760 (
        .din(new_Jinkela_wire_989),
        .dout(new_Jinkela_wire_990)
    );

    bfr new_Jinkela_buffer_744 (
        .din(new_Jinkela_wire_965),
        .dout(new_Jinkela_wire_966)
    );

    bfr new_Jinkela_buffer_745 (
        .din(new_Jinkela_wire_966),
        .dout(new_Jinkela_wire_967)
    );

    bfr new_Jinkela_buffer_761 (
        .din(new_Jinkela_wire_990),
        .dout(new_Jinkela_wire_991)
    );

    bfr new_Jinkela_buffer_746 (
        .din(new_Jinkela_wire_967),
        .dout(new_Jinkela_wire_968)
    );

    bfr new_Jinkela_buffer_783 (
        .din(new_Jinkela_wire_1020),
        .dout(new_Jinkela_wire_1021)
    );

    bfr new_Jinkela_buffer_747 (
        .din(new_Jinkela_wire_968),
        .dout(new_Jinkela_wire_969)
    );

    bfr new_Jinkela_buffer_762 (
        .din(new_Jinkela_wire_991),
        .dout(new_Jinkela_wire_992)
    );

    bfr new_Jinkela_buffer_748 (
        .din(new_Jinkela_wire_969),
        .dout(new_Jinkela_wire_970)
    );

    bfr new_Jinkela_buffer_834 (
        .din(N136),
        .dout(new_Jinkela_wire_1092)
    );

    bfr new_Jinkela_buffer_808 (
        .din(new_Jinkela_wire_1063),
        .dout(new_Jinkela_wire_1064)
    );

    bfr new_Jinkela_buffer_749 (
        .din(new_Jinkela_wire_970),
        .dout(new_Jinkela_wire_971)
    );

    bfr new_Jinkela_buffer_763 (
        .din(new_Jinkela_wire_992),
        .dout(new_Jinkela_wire_993)
    );

    bfr new_Jinkela_buffer_750 (
        .din(new_Jinkela_wire_971),
        .dout(new_Jinkela_wire_972)
    );

    bfr new_Jinkela_buffer_784 (
        .din(new_Jinkela_wire_1021),
        .dout(new_Jinkela_wire_1022)
    );

    bfr new_Jinkela_buffer_751 (
        .din(new_Jinkela_wire_972),
        .dout(new_Jinkela_wire_973)
    );

    bfr new_Jinkela_buffer_764 (
        .din(new_Jinkela_wire_993),
        .dout(new_Jinkela_wire_994)
    );

    bfr new_Jinkela_buffer_752 (
        .din(new_Jinkela_wire_973),
        .dout(new_Jinkela_wire_974)
    );

    bfr new_Jinkela_buffer_835 (
        .din(new_Jinkela_wire_1092),
        .dout(new_Jinkela_wire_1093)
    );

    spl2 new_Jinkela_splitter_83 (
        .a(new_Jinkela_wire_974),
        .b(new_Jinkela_wire_975),
        .c(new_Jinkela_wire_976)
    );

    bfr new_Jinkela_buffer_785 (
        .din(new_Jinkela_wire_1022),
        .dout(new_Jinkela_wire_1023)
    );

    bfr new_Jinkela_buffer_765 (
        .din(new_Jinkela_wire_994),
        .dout(new_Jinkela_wire_995)
    );

    bfr new_Jinkela_buffer_766 (
        .din(new_Jinkela_wire_995),
        .dout(new_Jinkela_wire_996)
    );

    bfr new_Jinkela_buffer_767 (
        .din(new_Jinkela_wire_996),
        .dout(new_Jinkela_wire_997)
    );

    bfr new_Jinkela_buffer_786 (
        .din(new_Jinkela_wire_1023),
        .dout(new_Jinkela_wire_1024)
    );

    bfr new_Jinkela_buffer_768 (
        .din(new_Jinkela_wire_997),
        .dout(new_Jinkela_wire_998)
    );

    bfr new_Jinkela_buffer_836 (
        .din(N129),
        .dout(new_Jinkela_wire_1094)
    );

    bfr new_Jinkela_buffer_807 (
        .din(new_Jinkela_wire_1057),
        .dout(new_Jinkela_wire_1058)
    );

    bfr new_Jinkela_buffer_769 (
        .din(new_Jinkela_wire_998),
        .dout(new_Jinkela_wire_999)
    );

    bfr new_Jinkela_buffer_787 (
        .din(new_Jinkela_wire_1024),
        .dout(new_Jinkela_wire_1025)
    );

    bfr new_Jinkela_buffer_770 (
        .din(new_Jinkela_wire_999),
        .dout(new_Jinkela_wire_1000)
    );

    spl2 new_Jinkela_splitter_96 (
        .a(N65),
        .b(new_Jinkela_wire_1096),
        .c(new_Jinkela_wire_1098)
    );

    bfr new_Jinkela_buffer_771 (
        .din(new_Jinkela_wire_1000),
        .dout(new_Jinkela_wire_1001)
    );

    bfr new_Jinkela_buffer_788 (
        .din(new_Jinkela_wire_1025),
        .dout(new_Jinkela_wire_1026)
    );

    bfr new_Jinkela_buffer_772 (
        .din(new_Jinkela_wire_1001),
        .dout(new_Jinkela_wire_1002)
    );

    spl2 new_Jinkela_splitter_99 (
        .a(_075_),
        .b(new_Jinkela_wire_1130),
        .c(new_Jinkela_wire_1131)
    );

    bfr new_Jinkela_buffer_837 (
        .din(new_Jinkela_wire_1094),
        .dout(new_Jinkela_wire_1095)
    );

    bfr new_Jinkela_buffer_773 (
        .din(new_Jinkela_wire_1002),
        .dout(new_Jinkela_wire_1003)
    );

    bfr new_Jinkela_buffer_789 (
        .din(new_Jinkela_wire_1026),
        .dout(new_Jinkela_wire_1027)
    );

    bfr new_Jinkela_buffer_774 (
        .din(new_Jinkela_wire_1003),
        .dout(new_Jinkela_wire_1004)
    );

    bfr new_Jinkela_buffer_809 (
        .din(new_Jinkela_wire_1064),
        .dout(new_Jinkela_wire_1065)
    );

    bfr new_Jinkela_buffer_775 (
        .din(new_Jinkela_wire_1004),
        .dout(new_Jinkela_wire_1005)
    );

    bfr new_Jinkela_buffer_790 (
        .din(new_Jinkela_wire_1027),
        .dout(new_Jinkela_wire_1028)
    );

    spl2 new_Jinkela_splitter_214 (
        .a(_227_),
        .b(new_Jinkela_wire_1556),
        .c(new_Jinkela_wire_1557)
    );

    bfr new_Jinkela_buffer_1011 (
        .din(new_Jinkela_wire_1542),
        .dout(new_Jinkela_wire_1543)
    );

    bfr new_Jinkela_buffer_1013 (
        .din(new_Jinkela_wire_1546),
        .dout(new_Jinkela_wire_1547)
    );

    spl2 new_Jinkela_splitter_211 (
        .a(new_Jinkela_wire_1543),
        .b(new_Jinkela_wire_1544),
        .c(new_Jinkela_wire_1545)
    );

    bfr new_Jinkela_buffer_1014 (
        .din(new_Jinkela_wire_1547),
        .dout(new_Jinkela_wire_1548)
    );

    spl2 new_Jinkela_splitter_216 (
        .a(_235_),
        .b(new_Jinkela_wire_1565),
        .c(new_Jinkela_wire_1566)
    );

    spl2 new_Jinkela_splitter_215 (
        .a(_147_),
        .b(new_Jinkela_wire_1558),
        .c(new_Jinkela_wire_1559)
    );

    bfr new_Jinkela_buffer_1015 (
        .din(new_Jinkela_wire_1548),
        .dout(new_Jinkela_wire_1549)
    );

    bfr new_Jinkela_buffer_1018 (
        .din(new_Jinkela_wire_1559),
        .dout(new_Jinkela_wire_1560)
    );

    bfr new_Jinkela_buffer_1016 (
        .din(new_Jinkela_wire_1549),
        .dout(new_Jinkela_wire_1550)
    );

    spl2 new_Jinkela_splitter_217 (
        .a(_148_),
        .b(new_Jinkela_wire_1572),
        .c(new_Jinkela_wire_1573)
    );

    bfr new_Jinkela_buffer_1017 (
        .din(new_Jinkela_wire_1550),
        .dout(new_Jinkela_wire_1551)
    );

    spl2 new_Jinkela_splitter_212 (
        .a(new_Jinkela_wire_1551),
        .b(new_Jinkela_wire_1552),
        .c(new_Jinkela_wire_1553)
    );

    bfr new_Jinkela_buffer_1023 (
        .din(new_Jinkela_wire_1566),
        .dout(new_Jinkela_wire_1567)
    );

    bfr new_Jinkela_buffer_1035 (
        .din(_011_),
        .dout(new_Jinkela_wire_1581)
    );

    bfr new_Jinkela_buffer_1019 (
        .din(new_Jinkela_wire_1560),
        .dout(new_Jinkela_wire_1561)
    );

    bfr new_Jinkela_buffer_1020 (
        .din(new_Jinkela_wire_1561),
        .dout(new_Jinkela_wire_1562)
    );

    spl4L new_Jinkela_splitter_219 (
        .a(_032_),
        .d(new_Jinkela_wire_1587),
        .e(new_Jinkela_wire_1588),
        .b(new_Jinkela_wire_1589),
        .c(new_Jinkela_wire_1590)
    );

    bfr new_Jinkela_buffer_1021 (
        .din(new_Jinkela_wire_1562),
        .dout(new_Jinkela_wire_1563)
    );

    bfr new_Jinkela_buffer_1024 (
        .din(new_Jinkela_wire_1567),
        .dout(new_Jinkela_wire_1568)
    );

    bfr new_Jinkela_buffer_1022 (
        .din(new_Jinkela_wire_1563),
        .dout(new_Jinkela_wire_1564)
    );

    bfr new_Jinkela_buffer_1028 (
        .din(new_Jinkela_wire_1573),
        .dout(new_Jinkela_wire_1574)
    );

    bfr new_Jinkela_buffer_1025 (
        .din(new_Jinkela_wire_1568),
        .dout(new_Jinkela_wire_1569)
    );

    spl2 new_Jinkela_splitter_220 (
        .a(_342_),
        .b(new_Jinkela_wire_1591),
        .c(new_Jinkela_wire_1592)
    );

    bfr new_Jinkela_buffer_1026 (
        .din(new_Jinkela_wire_1569),
        .dout(new_Jinkela_wire_1570)
    );

    bfr new_Jinkela_buffer_1029 (
        .din(new_Jinkela_wire_1574),
        .dout(new_Jinkela_wire_1575)
    );

    bfr new_Jinkela_buffer_1027 (
        .din(new_Jinkela_wire_1570),
        .dout(new_Jinkela_wire_1571)
    );

    bfr new_Jinkela_buffer_1036 (
        .din(new_Jinkela_wire_1581),
        .dout(new_Jinkela_wire_1582)
    );

    bfr new_Jinkela_buffer_1030 (
        .din(new_Jinkela_wire_1575),
        .dout(new_Jinkela_wire_1576)
    );

    spl3L new_Jinkela_splitter_221 (
        .a(_010_),
        .d(new_Jinkela_wire_1593),
        .b(new_Jinkela_wire_1594),
        .c(new_Jinkela_wire_1595)
    );

    bfr new_Jinkela_buffer_1031 (
        .din(new_Jinkela_wire_1576),
        .dout(new_Jinkela_wire_1577)
    );

    bfr new_Jinkela_buffer_1037 (
        .din(new_Jinkela_wire_1582),
        .dout(new_Jinkela_wire_1583)
    );

    bfr new_Jinkela_buffer_1032 (
        .din(new_Jinkela_wire_1577),
        .dout(new_Jinkela_wire_1578)
    );

    spl2 new_Jinkela_splitter_225 (
        .a(_290_),
        .b(new_Jinkela_wire_1615),
        .c(new_Jinkela_wire_1616)
    );

    bfr new_Jinkela_buffer_1033 (
        .din(new_Jinkela_wire_1578),
        .dout(new_Jinkela_wire_1579)
    );

    bfr new_Jinkela_buffer_1038 (
        .din(new_Jinkela_wire_1583),
        .dout(new_Jinkela_wire_1584)
    );

    bfr new_Jinkela_buffer_1034 (
        .din(new_Jinkela_wire_1579),
        .dout(new_Jinkela_wire_1580)
    );

    spl2 new_Jinkela_splitter_226 (
        .a(_082_),
        .b(new_Jinkela_wire_1617),
        .c(new_Jinkela_wire_1618)
    );

    spl2 new_Jinkela_splitter_218 (
        .a(new_Jinkela_wire_1584),
        .b(new_Jinkela_wire_1585),
        .c(new_Jinkela_wire_1586)
    );

    spl2 new_Jinkela_splitter_224 (
        .a(_272_),
        .b(new_Jinkela_wire_1613),
        .c(new_Jinkela_wire_1614)
    );

    spl2 new_Jinkela_splitter_223 (
        .a(_086_),
        .b(new_Jinkela_wire_1611),
        .c(new_Jinkela_wire_1612)
    );

    bfr new_Jinkela_buffer_1039 (
        .din(new_Jinkela_wire_1595),
        .dout(new_Jinkela_wire_1596)
    );

    bfr new_Jinkela_buffer_1040 (
        .din(new_Jinkela_wire_1596),
        .dout(new_Jinkela_wire_1597)
    );

    bfr new_Jinkela_buffer_132 (
        .din(new_Jinkela_wire_169),
        .dout(new_Jinkela_wire_170)
    );

    and_bi _433_ (
        .a(new_Jinkela_wire_1371),
        .b(new_Jinkela_wire_1537),
        .c(_045_)
    );

    bfr new_Jinkela_buffer_187 (
        .din(new_Jinkela_wire_243),
        .dout(new_Jinkela_wire_244)
    );

    and_bi _434_ (
        .a(new_Jinkela_wire_1536),
        .b(new_Jinkela_wire_1370),
        .c(_046_)
    );

    spl2 new_Jinkela_splitter_14 (
        .a(new_Jinkela_wire_170),
        .b(new_Jinkela_wire_171),
        .c(new_Jinkela_wire_172)
    );

    or_bb _435_ (
        .a(_046_),
        .b(_045_),
        .c(_047_)
    );

    bfr new_Jinkela_buffer_165 (
        .din(new_Jinkela_wire_218),
        .dout(new_Jinkela_wire_219)
    );

    or_ii _436_ (
        .a(new_Jinkela_wire_1093),
        .b(new_Jinkela_wire_1053),
        .c(_048_)
    );

    bfr new_Jinkela_buffer_145 (
        .din(new_Jinkela_wire_190),
        .dout(new_Jinkela_wire_191)
    );

    or_bi _437_ (
        .a(new_Jinkela_wire_809),
        .b(new_Jinkela_wire_352),
        .c(_049_)
    );

    bfr new_Jinkela_buffer_146 (
        .din(new_Jinkela_wire_191),
        .dout(new_Jinkela_wire_192)
    );

    and_bi _438_ (
        .a(new_Jinkela_wire_810),
        .b(new_Jinkela_wire_353),
        .c(_050_)
    );

    bfr new_Jinkela_buffer_240 (
        .din(N131),
        .dout(new_Jinkela_wire_312)
    );

    or_bi _439_ (
        .a(_050_),
        .b(_049_),
        .c(_051_)
    );

    bfr new_Jinkela_buffer_147 (
        .din(new_Jinkela_wire_192),
        .dout(new_Jinkela_wire_193)
    );

    or_bi _440_ (
        .a(new_Jinkela_wire_246),
        .b(new_Jinkela_wire_144),
        .c(_052_)
    );

    bfr new_Jinkela_buffer_166 (
        .din(new_Jinkela_wire_219),
        .dout(new_Jinkela_wire_220)
    );

    and_bi _441_ (
        .a(new_Jinkela_wire_244),
        .b(new_Jinkela_wire_143),
        .c(_053_)
    );

    bfr new_Jinkela_buffer_148 (
        .din(new_Jinkela_wire_193),
        .dout(new_Jinkela_wire_194)
    );

    or_bi _442_ (
        .a(_053_),
        .b(_052_),
        .c(_054_)
    );

    or_bi _443_ (
        .a(new_Jinkela_wire_1695),
        .b(new_Jinkela_wire_1134),
        .c(_055_)
    );

    bfr new_Jinkela_buffer_188 (
        .din(new_Jinkela_wire_249),
        .dout(new_Jinkela_wire_250)
    );

    bfr new_Jinkela_buffer_149 (
        .din(new_Jinkela_wire_194),
        .dout(new_Jinkela_wire_195)
    );

    and_bi _444_ (
        .a(new_Jinkela_wire_1694),
        .b(new_Jinkela_wire_1133),
        .c(_056_)
    );

    bfr new_Jinkela_buffer_167 (
        .din(new_Jinkela_wire_220),
        .dout(new_Jinkela_wire_221)
    );

    or_bi _445_ (
        .a(_056_),
        .b(_055_),
        .c(_057_)
    );

    bfr new_Jinkela_buffer_150 (
        .din(new_Jinkela_wire_195),
        .dout(new_Jinkela_wire_196)
    );

    or_bi _446_ (
        .a(new_Jinkela_wire_1327),
        .b(new_Jinkela_wire_1533),
        .c(_058_)
    );

    and_bi _447_ (
        .a(new_Jinkela_wire_1326),
        .b(new_Jinkela_wire_1532),
        .c(_059_)
    );

    bfr new_Jinkela_buffer_241 (
        .din(new_Jinkela_wire_312),
        .dout(new_Jinkela_wire_313)
    );

    and_bi _410_ (
        .a(new_Jinkela_wire_1585),
        .b(new_Jinkela_wire_1139),
        .c(_022_)
    );

    bfr new_Jinkela_buffer_151 (
        .din(new_Jinkela_wire_196),
        .dout(new_Jinkela_wire_197)
    );

    and_bi _448_ (
        .a(_058_),
        .b(_059_),
        .c(_060_)
    );

    bfr new_Jinkela_buffer_168 (
        .din(new_Jinkela_wire_221),
        .dout(new_Jinkela_wire_222)
    );

    or_bb _449_ (
        .a(new_Jinkela_wire_911),
        .b(new_Jinkela_wire_315),
        .c(_061_)
    );

    bfr new_Jinkela_buffer_152 (
        .din(new_Jinkela_wire_197),
        .dout(new_Jinkela_wire_198)
    );

    and_bb _450_ (
        .a(new_Jinkela_wire_913),
        .b(new_Jinkela_wire_317),
        .c(_062_)
    );

    and_bi _451_ (
        .a(_061_),
        .b(_062_),
        .c(_063_)
    );

    bfr new_Jinkela_buffer_214 (
        .din(new_Jinkela_wire_283),
        .dout(new_Jinkela_wire_284)
    );

    bfr new_Jinkela_buffer_153 (
        .din(new_Jinkela_wire_198),
        .dout(new_Jinkela_wire_199)
    );

    or_bi _452_ (
        .a(new_Jinkela_wire_529),
        .b(new_Jinkela_wire_174),
        .c(_064_)
    );

    bfr new_Jinkela_buffer_169 (
        .din(new_Jinkela_wire_222),
        .dout(new_Jinkela_wire_223)
    );

    and_bi _453_ (
        .a(new_Jinkela_wire_528),
        .b(new_Jinkela_wire_176),
        .c(_065_)
    );

    bfr new_Jinkela_buffer_154 (
        .din(new_Jinkela_wire_199),
        .dout(new_Jinkela_wire_200)
    );

    or_bi _454_ (
        .a(_065_),
        .b(_064_),
        .c(_066_)
    );

    spl4L new_Jinkela_splitter_31 (
        .a(new_Jinkela_wire_351),
        .d(new_Jinkela_wire_352),
        .e(new_Jinkela_wire_353),
        .b(new_Jinkela_wire_354),
        .c(new_Jinkela_wire_355)
    );

    or_bi _455_ (
        .a(new_Jinkela_wire_1657),
        .b(new_Jinkela_wire_1502),
        .c(_067_)
    );

    bfr new_Jinkela_buffer_189 (
        .din(new_Jinkela_wire_250),
        .dout(new_Jinkela_wire_251)
    );

    bfr new_Jinkela_buffer_155 (
        .din(new_Jinkela_wire_200),
        .dout(new_Jinkela_wire_201)
    );

    and_bi _456_ (
        .a(new_Jinkela_wire_1656),
        .b(new_Jinkela_wire_1501),
        .c(_068_)
    );

    bfr new_Jinkela_buffer_170 (
        .din(new_Jinkela_wire_223),
        .dout(new_Jinkela_wire_224)
    );

    and_bi _457_ (
        .a(_067_),
        .b(_068_),
        .c(_069_)
    );

    bfr new_Jinkela_buffer_156 (
        .din(new_Jinkela_wire_201),
        .dout(new_Jinkela_wire_202)
    );

    or_bb _458_ (
        .a(new_Jinkela_wire_426),
        .b(new_Jinkela_wire_109),
        .c(_070_)
    );

    and_bb _459_ (
        .a(new_Jinkela_wire_423),
        .b(new_Jinkela_wire_107),
        .c(_071_)
    );

    bfr new_Jinkela_buffer_157 (
        .din(new_Jinkela_wire_202),
        .dout(new_Jinkela_wire_203)
    );

    and_bi _460_ (
        .a(_070_),
        .b(_071_),
        .c(_072_)
    );

    bfr new_Jinkela_buffer_171 (
        .din(new_Jinkela_wire_224),
        .dout(new_Jinkela_wire_225)
    );

    or_bi _461_ (
        .a(new_Jinkela_wire_844),
        .b(new_Jinkela_wire_212),
        .c(_073_)
    );

    bfr new_Jinkela_buffer_158 (
        .din(new_Jinkela_wire_203),
        .dout(new_Jinkela_wire_204)
    );

    and_bi _462_ (
        .a(new_Jinkela_wire_842),
        .b(new_Jinkela_wire_213),
        .c(_074_)
    );

    or_bi _463_ (
        .a(_074_),
        .b(_073_),
        .c(_075_)
    );

    bfr new_Jinkela_buffer_190 (
        .din(new_Jinkela_wire_251),
        .dout(new_Jinkela_wire_252)
    );

    bfr new_Jinkela_buffer_159 (
        .din(new_Jinkela_wire_204),
        .dout(new_Jinkela_wire_205)
    );

    or_bi _464_ (
        .a(new_Jinkela_wire_1332),
        .b(new_Jinkela_wire_1131),
        .c(_076_)
    );

    bfr new_Jinkela_buffer_172 (
        .din(new_Jinkela_wire_225),
        .dout(new_Jinkela_wire_226)
    );

    and_bi _465_ (
        .a(new_Jinkela_wire_1331),
        .b(new_Jinkela_wire_1130),
        .c(_077_)
    );

    spl2 new_Jinkela_splitter_17 (
        .a(new_Jinkela_wire_205),
        .b(new_Jinkela_wire_206),
        .c(new_Jinkela_wire_207)
    );

    and_bi _466_ (
        .a(new_Jinkela_wire_1281),
        .b(new_Jinkela_wire_1672),
        .c(_078_)
    );

    bfr new_Jinkela_buffer_173 (
        .din(new_Jinkela_wire_226),
        .dout(new_Jinkela_wire_227)
    );

    or_bb _467_ (
        .a(new_Jinkela_wire_1379),
        .b(new_Jinkela_wire_1630),
        .c(_079_)
    );

    or_bi _468_ (
        .a(new_Jinkela_wire_1671),
        .b(new_Jinkela_wire_1280),
        .c(_080_)
    );

    spl2 new_Jinkela_splitter_27 (
        .a(N25),
        .b(new_Jinkela_wire_314),
        .c(new_Jinkela_wire_316)
    );

    bfr new_Jinkela_buffer_213 (
        .din(new_Jinkela_wire_277),
        .dout(new_Jinkela_wire_278)
    );

    and_bi _469_ (
        .a(new_Jinkela_wire_1629),
        .b(new_Jinkela_wire_1680),
        .c(_081_)
    );

    bfr new_Jinkela_buffer_191 (
        .din(new_Jinkela_wire_252),
        .dout(new_Jinkela_wire_253)
    );

    bfr new_Jinkela_buffer_174 (
        .din(new_Jinkela_wire_227),
        .dout(new_Jinkela_wire_228)
    );

    and_bi _470_ (
        .a(_079_),
        .b(_081_),
        .c(_082_)
    );

    and_bi _471_ (
        .a(new_Jinkela_wire_1618),
        .b(new_Jinkela_wire_1449),
        .c(_083_)
    );

    bfr new_Jinkela_buffer_175 (
        .din(new_Jinkela_wire_228),
        .dout(new_Jinkela_wire_229)
    );

    and_bi _472_ (
        .a(new_Jinkela_wire_1448),
        .b(new_Jinkela_wire_1617),
        .c(_084_)
    );

    or_bb _473_ (
        .a(_084_),
        .b(_083_),
        .c(_085_)
    );

    spl4L new_Jinkela_splitter_25 (
        .a(new_Jinkela_wire_279),
        .d(new_Jinkela_wire_280),
        .e(new_Jinkela_wire_281),
        .b(new_Jinkela_wire_282),
        .c(new_Jinkela_wire_283)
    );

    bfr new_Jinkela_buffer_176 (
        .din(new_Jinkela_wire_229),
        .dout(new_Jinkela_wire_230)
    );

    and_bi _474_ (
        .a(new_Jinkela_wire_1260),
        .b(new_Jinkela_wire_1452),
        .c(_086_)
    );

    bfr new_Jinkela_buffer_554 (
        .din(new_Jinkela_wire_719),
        .dout(new_Jinkela_wire_720)
    );

    bfr new_Jinkela_buffer_596 (
        .din(new_Jinkela_wire_777),
        .dout(new_Jinkela_wire_778)
    );

    bfr new_Jinkela_buffer_555 (
        .din(new_Jinkela_wire_720),
        .dout(new_Jinkela_wire_721)
    );

    bfr new_Jinkela_buffer_572 (
        .din(new_Jinkela_wire_745),
        .dout(new_Jinkela_wire_746)
    );

    bfr new_Jinkela_buffer_556 (
        .din(new_Jinkela_wire_721),
        .dout(new_Jinkela_wire_722)
    );

    bfr new_Jinkela_buffer_621 (
        .din(new_Jinkela_wire_805),
        .dout(new_Jinkela_wire_806)
    );

    bfr new_Jinkela_buffer_557 (
        .din(new_Jinkela_wire_722),
        .dout(new_Jinkela_wire_723)
    );

    bfr new_Jinkela_buffer_573 (
        .din(new_Jinkela_wire_746),
        .dout(new_Jinkela_wire_747)
    );

    bfr new_Jinkela_buffer_558 (
        .din(new_Jinkela_wire_723),
        .dout(new_Jinkela_wire_724)
    );

    spl2 new_Jinkela_splitter_75 (
        .a(N69),
        .b(new_Jinkela_wire_874),
        .c(new_Jinkela_wire_876)
    );

    bfr new_Jinkela_buffer_622 (
        .din(new_Jinkela_wire_811),
        .dout(new_Jinkela_wire_812)
    );

    bfr new_Jinkela_buffer_559 (
        .din(new_Jinkela_wire_724),
        .dout(new_Jinkela_wire_725)
    );

    bfr new_Jinkela_buffer_574 (
        .din(new_Jinkela_wire_747),
        .dout(new_Jinkela_wire_748)
    );

    bfr new_Jinkela_buffer_560 (
        .din(new_Jinkela_wire_725),
        .dout(new_Jinkela_wire_726)
    );

    bfr new_Jinkela_buffer_597 (
        .din(new_Jinkela_wire_778),
        .dout(new_Jinkela_wire_779)
    );

    bfr new_Jinkela_buffer_561 (
        .din(new_Jinkela_wire_726),
        .dout(new_Jinkela_wire_727)
    );

    bfr new_Jinkela_buffer_575 (
        .din(new_Jinkela_wire_748),
        .dout(new_Jinkela_wire_749)
    );

    bfr new_Jinkela_buffer_562 (
        .din(new_Jinkela_wire_727),
        .dout(new_Jinkela_wire_728)
    );

    bfr new_Jinkela_buffer_563 (
        .din(new_Jinkela_wire_728),
        .dout(new_Jinkela_wire_729)
    );

    bfr new_Jinkela_buffer_576 (
        .din(new_Jinkela_wire_749),
        .dout(new_Jinkela_wire_750)
    );

    spl2 new_Jinkela_splitter_62 (
        .a(new_Jinkela_wire_729),
        .b(new_Jinkela_wire_730),
        .c(new_Jinkela_wire_731)
    );

    bfr new_Jinkela_buffer_577 (
        .din(new_Jinkela_wire_750),
        .dout(new_Jinkela_wire_751)
    );

    bfr new_Jinkela_buffer_598 (
        .din(new_Jinkela_wire_779),
        .dout(new_Jinkela_wire_780)
    );

    bfr new_Jinkela_buffer_578 (
        .din(new_Jinkela_wire_751),
        .dout(new_Jinkela_wire_752)
    );

    bfr new_Jinkela_buffer_599 (
        .din(new_Jinkela_wire_780),
        .dout(new_Jinkela_wire_781)
    );

    bfr new_Jinkela_buffer_579 (
        .din(new_Jinkela_wire_752),
        .dout(new_Jinkela_wire_753)
    );

    spl4L new_Jinkela_splitter_73 (
        .a(new_Jinkela_wire_841),
        .d(new_Jinkela_wire_842),
        .e(new_Jinkela_wire_843),
        .b(new_Jinkela_wire_844),
        .c(new_Jinkela_wire_845)
    );

    bfr new_Jinkela_buffer_580 (
        .din(new_Jinkela_wire_753),
        .dout(new_Jinkela_wire_754)
    );

    bfr new_Jinkela_buffer_600 (
        .din(new_Jinkela_wire_781),
        .dout(new_Jinkela_wire_782)
    );

    bfr new_Jinkela_buffer_581 (
        .din(new_Jinkela_wire_754),
        .dout(new_Jinkela_wire_755)
    );

    bfr new_Jinkela_buffer_647 (
        .din(new_Jinkela_wire_839),
        .dout(new_Jinkela_wire_840)
    );

    bfr new_Jinkela_buffer_582 (
        .din(new_Jinkela_wire_755),
        .dout(new_Jinkela_wire_756)
    );

    bfr new_Jinkela_buffer_601 (
        .din(new_Jinkela_wire_782),
        .dout(new_Jinkela_wire_783)
    );

    bfr new_Jinkela_buffer_583 (
        .din(new_Jinkela_wire_756),
        .dout(new_Jinkela_wire_757)
    );

    bfr new_Jinkela_buffer_623 (
        .din(new_Jinkela_wire_812),
        .dout(new_Jinkela_wire_813)
    );

    bfr new_Jinkela_buffer_584 (
        .din(new_Jinkela_wire_757),
        .dout(new_Jinkela_wire_758)
    );

    bfr new_Jinkela_buffer_602 (
        .din(new_Jinkela_wire_783),
        .dout(new_Jinkela_wire_784)
    );

    bfr new_Jinkela_buffer_585 (
        .din(new_Jinkela_wire_758),
        .dout(new_Jinkela_wire_759)
    );

    spl4L new_Jinkela_splitter_76 (
        .a(new_Jinkela_wire_876),
        .d(new_Jinkela_wire_877),
        .e(new_Jinkela_wire_878),
        .b(new_Jinkela_wire_879),
        .c(new_Jinkela_wire_880)
    );

    spl2 new_Jinkela_splitter_78 (
        .a(N29),
        .b(new_Jinkela_wire_908),
        .c(new_Jinkela_wire_910)
    );

    bfr new_Jinkela_buffer_586 (
        .din(new_Jinkela_wire_759),
        .dout(new_Jinkela_wire_760)
    );

    bfr new_Jinkela_buffer_603 (
        .din(new_Jinkela_wire_784),
        .dout(new_Jinkela_wire_785)
    );

    bfr new_Jinkela_buffer_776 (
        .din(new_Jinkela_wire_1005),
        .dout(new_Jinkela_wire_1006)
    );

    bfr new_Jinkela_buffer_864 (
        .din(new_net_711),
        .dout(new_Jinkela_wire_1132)
    );

    bfr new_Jinkela_buffer_777 (
        .din(new_Jinkela_wire_1006),
        .dout(new_Jinkela_wire_1007)
    );

    bfr new_Jinkela_buffer_791 (
        .din(new_Jinkela_wire_1028),
        .dout(new_Jinkela_wire_1029)
    );

    bfr new_Jinkela_buffer_778 (
        .din(new_Jinkela_wire_1007),
        .dout(new_Jinkela_wire_1008)
    );

    bfr new_Jinkela_buffer_810 (
        .din(new_Jinkela_wire_1065),
        .dout(new_Jinkela_wire_1066)
    );

    bfr new_Jinkela_buffer_779 (
        .din(new_Jinkela_wire_1008),
        .dout(new_Jinkela_wire_1009)
    );

    bfr new_Jinkela_buffer_792 (
        .din(new_Jinkela_wire_1029),
        .dout(new_Jinkela_wire_1030)
    );

    spl2 new_Jinkela_splitter_86 (
        .a(new_Jinkela_wire_1009),
        .b(new_Jinkela_wire_1010),
        .c(new_Jinkela_wire_1011)
    );

    bfr new_Jinkela_buffer_793 (
        .din(new_Jinkela_wire_1030),
        .dout(new_Jinkela_wire_1031)
    );

    bfr new_Jinkela_buffer_838 (
        .din(new_Jinkela_wire_1096),
        .dout(new_Jinkela_wire_1097)
    );

    bfr new_Jinkela_buffer_811 (
        .din(new_Jinkela_wire_1066),
        .dout(new_Jinkela_wire_1067)
    );

    bfr new_Jinkela_buffer_794 (
        .din(new_Jinkela_wire_1031),
        .dout(new_Jinkela_wire_1032)
    );

    bfr new_Jinkela_buffer_795 (
        .din(new_Jinkela_wire_1032),
        .dout(new_Jinkela_wire_1033)
    );

    bfr new_Jinkela_buffer_812 (
        .din(new_Jinkela_wire_1067),
        .dout(new_Jinkela_wire_1068)
    );

    bfr new_Jinkela_buffer_796 (
        .din(new_Jinkela_wire_1033),
        .dout(new_Jinkela_wire_1034)
    );

    spl4L new_Jinkela_splitter_97 (
        .a(new_Jinkela_wire_1098),
        .d(new_Jinkela_wire_1099),
        .e(new_Jinkela_wire_1100),
        .b(new_Jinkela_wire_1101),
        .c(new_Jinkela_wire_1102)
    );

    bfr new_Jinkela_buffer_797 (
        .din(new_Jinkela_wire_1034),
        .dout(new_Jinkela_wire_1035)
    );

    bfr new_Jinkela_buffer_813 (
        .din(new_Jinkela_wire_1068),
        .dout(new_Jinkela_wire_1069)
    );

    bfr new_Jinkela_buffer_798 (
        .din(new_Jinkela_wire_1035),
        .dout(new_Jinkela_wire_1036)
    );

    bfr new_Jinkela_buffer_865 (
        .din(new_net_697),
        .dout(new_Jinkela_wire_1135)
    );

    bfr new_Jinkela_buffer_799 (
        .din(new_Jinkela_wire_1036),
        .dout(new_Jinkela_wire_1037)
    );

    bfr new_Jinkela_buffer_814 (
        .din(new_Jinkela_wire_1069),
        .dout(new_Jinkela_wire_1070)
    );

    bfr new_Jinkela_buffer_800 (
        .din(new_Jinkela_wire_1037),
        .dout(new_Jinkela_wire_1038)
    );

    bfr new_Jinkela_buffer_839 (
        .din(new_Jinkela_wire_1102),
        .dout(new_Jinkela_wire_1103)
    );

    bfr new_Jinkela_buffer_801 (
        .din(new_Jinkela_wire_1038),
        .dout(new_Jinkela_wire_1039)
    );

    bfr new_Jinkela_buffer_815 (
        .din(new_Jinkela_wire_1070),
        .dout(new_Jinkela_wire_1071)
    );

    bfr new_Jinkela_buffer_802 (
        .din(new_Jinkela_wire_1039),
        .dout(new_Jinkela_wire_1040)
    );

    spl2 new_Jinkela_splitter_100 (
        .a(_054_),
        .b(new_Jinkela_wire_1133),
        .c(new_Jinkela_wire_1134)
    );

    bfr new_Jinkela_buffer_803 (
        .din(new_Jinkela_wire_1040),
        .dout(new_Jinkela_wire_1041)
    );

    bfr new_Jinkela_buffer_816 (
        .din(new_Jinkela_wire_1071),
        .dout(new_Jinkela_wire_1072)
    );

    bfr new_Jinkela_buffer_804 (
        .din(new_Jinkela_wire_1041),
        .dout(new_Jinkela_wire_1042)
    );

    bfr new_Jinkela_buffer_867 (
        .din(_174_),
        .dout(new_Jinkela_wire_1137)
    );

    bfr new_Jinkela_buffer_805 (
        .din(new_Jinkela_wire_1042),
        .dout(new_Jinkela_wire_1043)
    );

    bfr new_Jinkela_buffer_817 (
        .din(new_Jinkela_wire_1072),
        .dout(new_Jinkela_wire_1073)
    );

    bfr new_Jinkela_buffer_806 (
        .din(new_Jinkela_wire_1043),
        .dout(new_Jinkela_wire_1044)
    );

    bfr new_Jinkela_buffer_840 (
        .din(new_Jinkela_wire_1103),
        .dout(new_Jinkela_wire_1104)
    );

    spl2 new_Jinkela_splitter_89 (
        .a(new_Jinkela_wire_1044),
        .b(new_Jinkela_wire_1045),
        .c(new_Jinkela_wire_1046)
    );

    bfr new_Jinkela_buffer_866 (
        .din(_240_),
        .dout(new_Jinkela_wire_1136)
    );

    bfr new_Jinkela_buffer_818 (
        .din(new_Jinkela_wire_1073),
        .dout(new_Jinkela_wire_1074)
    );

    bfr new_Jinkela_buffer_819 (
        .din(new_Jinkela_wire_1074),
        .dout(new_Jinkela_wire_1075)
    );

    bfr new_Jinkela_buffer_385 (
        .din(new_Jinkela_wire_502),
        .dout(new_Jinkela_wire_503)
    );

    bfr new_Jinkela_buffer_917 (
        .din(new_Jinkela_wire_1248),
        .dout(new_Jinkela_wire_1249)
    );

    bfr new_Jinkela_buffer_368 (
        .din(new_Jinkela_wire_477),
        .dout(new_Jinkela_wire_478)
    );

    spl2 new_Jinkela_splitter_137 (
        .a(_214_),
        .b(new_Jinkela_wire_1289),
        .c(new_Jinkela_wire_1290)
    );

    bfr new_Jinkela_buffer_1041 (
        .din(new_Jinkela_wire_1597),
        .dout(new_Jinkela_wire_1598)
    );

    bfr new_Jinkela_buffer_407 (
        .din(new_Jinkela_wire_532),
        .dout(new_Jinkela_wire_533)
    );

    bfr new_Jinkela_buffer_923 (
        .din(new_Jinkela_wire_1264),
        .dout(new_Jinkela_wire_1265)
    );

    bfr new_Jinkela_buffer_918 (
        .din(new_Jinkela_wire_1249),
        .dout(new_Jinkela_wire_1250)
    );

    bfr new_Jinkela_buffer_369 (
        .din(new_Jinkela_wire_478),
        .dout(new_Jinkela_wire_479)
    );

    spl2 new_Jinkela_splitter_227 (
        .a(_160_),
        .b(new_Jinkela_wire_1619),
        .c(new_Jinkela_wire_1620)
    );

    bfr new_Jinkela_buffer_1042 (
        .din(new_Jinkela_wire_1598),
        .dout(new_Jinkela_wire_1599)
    );

    bfr new_Jinkela_buffer_386 (
        .din(new_Jinkela_wire_503),
        .dout(new_Jinkela_wire_504)
    );

    spl2 new_Jinkela_splitter_135 (
        .a(new_Jinkela_wire_1284),
        .b(new_Jinkela_wire_1285),
        .c(new_Jinkela_wire_1286)
    );

    spl4L new_Jinkela_splitter_127 (
        .a(new_Jinkela_wire_1250),
        .d(new_Jinkela_wire_1251),
        .e(new_Jinkela_wire_1252),
        .b(new_Jinkela_wire_1253),
        .c(new_Jinkela_wire_1254)
    );

    bfr new_Jinkela_buffer_370 (
        .din(new_Jinkela_wire_479),
        .dout(new_Jinkela_wire_480)
    );

    bfr new_Jinkela_buffer_1050 (
        .din(_208_),
        .dout(new_Jinkela_wire_1621)
    );

    bfr new_Jinkela_buffer_1043 (
        .din(new_Jinkela_wire_1599),
        .dout(new_Jinkela_wire_1600)
    );

    spl2 new_Jinkela_splitter_138 (
        .a(_354_),
        .b(new_Jinkela_wire_1291),
        .c(new_Jinkela_wire_1292)
    );

    bfr new_Jinkela_buffer_924 (
        .din(new_Jinkela_wire_1265),
        .dout(new_Jinkela_wire_1266)
    );

    spl2 new_Jinkela_splitter_228 (
        .a(new_Jinkela_wire_1621),
        .b(new_Jinkela_wire_1622),
        .c(new_Jinkela_wire_1623)
    );

    bfr new_Jinkela_buffer_371 (
        .din(new_Jinkela_wire_480),
        .dout(new_Jinkela_wire_481)
    );

    bfr new_Jinkela_buffer_925 (
        .din(new_Jinkela_wire_1266),
        .dout(new_Jinkela_wire_1267)
    );

    bfr new_Jinkela_buffer_1044 (
        .din(new_Jinkela_wire_1600),
        .dout(new_Jinkela_wire_1601)
    );

    bfr new_Jinkela_buffer_387 (
        .din(new_Jinkela_wire_504),
        .dout(new_Jinkela_wire_505)
    );

    spl2 new_Jinkela_splitter_141 (
        .a(_193_),
        .b(new_Jinkela_wire_1297),
        .c(new_Jinkela_wire_1298)
    );

    spl2 new_Jinkela_splitter_229 (
        .a(_266_),
        .b(new_Jinkela_wire_1624),
        .c(new_Jinkela_wire_1625)
    );

    bfr new_Jinkela_buffer_372 (
        .din(new_Jinkela_wire_481),
        .dout(new_Jinkela_wire_482)
    );

    bfr new_Jinkela_buffer_926 (
        .din(new_Jinkela_wire_1267),
        .dout(new_Jinkela_wire_1268)
    );

    bfr new_Jinkela_buffer_1045 (
        .din(new_Jinkela_wire_1601),
        .dout(new_Jinkela_wire_1602)
    );

    bfr new_Jinkela_buffer_408 (
        .din(new_Jinkela_wire_533),
        .dout(new_Jinkela_wire_534)
    );

    spl3L new_Jinkela_splitter_230 (
        .a(_069_),
        .d(new_Jinkela_wire_1626),
        .b(new_Jinkela_wire_1627),
        .c(new_Jinkela_wire_1628)
    );

    bfr new_Jinkela_buffer_373 (
        .din(new_Jinkela_wire_482),
        .dout(new_Jinkela_wire_483)
    );

    spl2 new_Jinkela_splitter_139 (
        .a(_245_),
        .b(new_Jinkela_wire_1293),
        .c(new_Jinkela_wire_1294)
    );

    bfr new_Jinkela_buffer_1051 (
        .din(_199_),
        .dout(new_Jinkela_wire_1631)
    );

    bfr new_Jinkela_buffer_927 (
        .din(new_Jinkela_wire_1268),
        .dout(new_Jinkela_wire_1269)
    );

    bfr new_Jinkela_buffer_1046 (
        .din(new_Jinkela_wire_1602),
        .dout(new_Jinkela_wire_1603)
    );

    bfr new_Jinkela_buffer_388 (
        .din(new_Jinkela_wire_505),
        .dout(new_Jinkela_wire_506)
    );

    spl2 new_Jinkela_splitter_233 (
        .a(_321_),
        .b(new_Jinkela_wire_1634),
        .c(new_Jinkela_wire_1635)
    );

    bfr new_Jinkela_buffer_374 (
        .din(new_Jinkela_wire_483),
        .dout(new_Jinkela_wire_484)
    );

    bfr new_Jinkela_buffer_928 (
        .din(new_Jinkela_wire_1269),
        .dout(new_Jinkela_wire_1270)
    );

    bfr new_Jinkela_buffer_1047 (
        .din(new_Jinkela_wire_1603),
        .dout(new_Jinkela_wire_1604)
    );

    spl2 new_Jinkela_splitter_54 (
        .a(N81),
        .b(new_Jinkela_wire_629),
        .c(new_Jinkela_wire_631)
    );

    spl2 new_Jinkela_splitter_140 (
        .a(_260_),
        .b(new_Jinkela_wire_1295),
        .c(new_Jinkela_wire_1296)
    );

    bfr new_Jinkela_buffer_375 (
        .din(new_Jinkela_wire_484),
        .dout(new_Jinkela_wire_485)
    );

    spl2 new_Jinkela_splitter_235 (
        .a(_095_),
        .b(new_Jinkela_wire_1638),
        .c(new_Jinkela_wire_1639)
    );

    bfr new_Jinkela_buffer_929 (
        .din(new_Jinkela_wire_1270),
        .dout(new_Jinkela_wire_1271)
    );

    bfr new_Jinkela_buffer_1048 (
        .din(new_Jinkela_wire_1604),
        .dout(new_Jinkela_wire_1605)
    );

    bfr new_Jinkela_buffer_389 (
        .din(new_Jinkela_wire_506),
        .dout(new_Jinkela_wire_507)
    );

    spl2 new_Jinkela_splitter_145 (
        .a(_282_),
        .b(new_Jinkela_wire_1310),
        .c(new_Jinkela_wire_1311)
    );

    spl2 new_Jinkela_splitter_231 (
        .a(new_Jinkela_wire_1628),
        .b(new_Jinkela_wire_1629),
        .c(new_Jinkela_wire_1630)
    );

    bfr new_Jinkela_buffer_376 (
        .din(new_Jinkela_wire_485),
        .dout(new_Jinkela_wire_486)
    );

    spl4L new_Jinkela_splitter_142 (
        .a(_289_),
        .d(new_Jinkela_wire_1299),
        .e(new_Jinkela_wire_1300),
        .b(new_Jinkela_wire_1301),
        .c(new_Jinkela_wire_1302)
    );

    spl2 new_Jinkela_splitter_234 (
        .a(_351_),
        .b(new_Jinkela_wire_1636),
        .c(new_Jinkela_wire_1637)
    );

    spl4L new_Jinkela_splitter_130 (
        .a(new_Jinkela_wire_1271),
        .d(new_Jinkela_wire_1272),
        .e(new_Jinkela_wire_1273),
        .b(new_Jinkela_wire_1274),
        .c(new_Jinkela_wire_1275)
    );

    bfr new_Jinkela_buffer_1049 (
        .din(new_Jinkela_wire_1605),
        .dout(new_Jinkela_wire_1606)
    );

    bfr new_Jinkela_buffer_409 (
        .din(new_Jinkela_wire_534),
        .dout(new_Jinkela_wire_535)
    );

    spl2 new_Jinkela_splitter_143 (
        .a(_132_),
        .b(new_Jinkela_wire_1303),
        .c(new_Jinkela_wire_1304)
    );

    bfr new_Jinkela_buffer_377 (
        .din(new_Jinkela_wire_486),
        .dout(new_Jinkela_wire_487)
    );

    spl4L new_Jinkela_splitter_222 (
        .a(new_Jinkela_wire_1606),
        .d(new_Jinkela_wire_1607),
        .e(new_Jinkela_wire_1608),
        .b(new_Jinkela_wire_1609),
        .c(new_Jinkela_wire_1610)
    );

    bfr new_Jinkela_buffer_390 (
        .din(new_Jinkela_wire_507),
        .dout(new_Jinkela_wire_508)
    );

    bfr new_Jinkela_buffer_931 (
        .din(new_net_687),
        .dout(new_Jinkela_wire_1305)
    );

    bfr new_Jinkela_buffer_378 (
        .din(new_Jinkela_wire_487),
        .dout(new_Jinkela_wire_488)
    );

    bfr new_Jinkela_buffer_433 (
        .din(new_Jinkela_wire_566),
        .dout(new_Jinkela_wire_567)
    );

    spl4L new_Jinkela_splitter_144 (
        .a(_275_),
        .d(new_Jinkela_wire_1306),
        .e(new_Jinkela_wire_1307),
        .b(new_Jinkela_wire_1308),
        .c(new_Jinkela_wire_1309)
    );

    spl2 new_Jinkela_splitter_232 (
        .a(new_Jinkela_wire_1631),
        .b(new_Jinkela_wire_1632),
        .c(new_Jinkela_wire_1633)
    );

    bfr new_Jinkela_buffer_932 (
        .din(_048_),
        .dout(new_Jinkela_wire_1322)
    );

    spl2 new_Jinkela_splitter_41 (
        .a(new_Jinkela_wire_488),
        .b(new_Jinkela_wire_489),
        .c(new_Jinkela_wire_490)
    );

    spl2 new_Jinkela_splitter_147 (
        .a(_126_),
        .b(new_Jinkela_wire_1314),
        .c(new_Jinkela_wire_1315)
    );

    spl2 new_Jinkela_splitter_236 (
        .a(_360_),
        .b(new_Jinkela_wire_1640),
        .c(new_Jinkela_wire_1641)
    );

    bfr new_Jinkela_buffer_410 (
        .din(new_Jinkela_wire_535),
        .dout(new_Jinkela_wire_536)
    );

    spl2 new_Jinkela_splitter_146 (
        .a(_254_),
        .b(new_Jinkela_wire_1312),
        .c(new_Jinkela_wire_1313)
    );

    bfr new_Jinkela_buffer_1057 (
        .din(new_net_715),
        .dout(new_Jinkela_wire_1651)
    );

    spl2 new_Jinkela_splitter_237 (
        .a(_218_),
        .b(new_Jinkela_wire_1642),
        .c(new_Jinkela_wire_1643)
    );

    bfr new_Jinkela_buffer_391 (
        .din(new_Jinkela_wire_508),
        .dout(new_Jinkela_wire_509)
    );

    spl2 new_Jinkela_splitter_148 (
        .a(_293_),
        .b(new_Jinkela_wire_1316),
        .c(new_Jinkela_wire_1317)
    );

    spl2 new_Jinkela_splitter_238 (
        .a(_215_),
        .b(new_Jinkela_wire_1644),
        .c(new_Jinkela_wire_1645)
    );

    bfr new_Jinkela_buffer_392 (
        .din(new_Jinkela_wire_509),
        .dout(new_Jinkela_wire_510)
    );

    spl4L new_Jinkela_splitter_149 (
        .a(_308_),
        .d(new_Jinkela_wire_1318),
        .e(new_Jinkela_wire_1319),
        .b(new_Jinkela_wire_1320),
        .c(new_Jinkela_wire_1321)
    );

    bfr new_Jinkela_buffer_1052 (
        .din(new_Jinkela_wire_1645),
        .dout(new_Jinkela_wire_1646)
    );

    bfr new_Jinkela_buffer_936 (
        .din(new_net_695),
        .dout(new_Jinkela_wire_1328)
    );

    bfr new_Jinkela_buffer_459 (
        .din(new_Jinkela_wire_595),
        .dout(new_Jinkela_wire_596)
    );

    spl2 new_Jinkela_splitter_239 (
        .a(_009_),
        .b(new_Jinkela_wire_1652),
        .c(new_Jinkela_wire_1653)
    );

    bfr new_Jinkela_buffer_393 (
        .din(new_Jinkela_wire_510),
        .dout(new_Jinkela_wire_511)
    );

    spl2 new_Jinkela_splitter_151 (
        .a(_202_),
        .b(new_Jinkela_wire_1329),
        .c(new_Jinkela_wire_1330)
    );

    spl2 new_Jinkela_splitter_240 (
        .a(_212_),
        .b(new_Jinkela_wire_1654),
        .c(new_Jinkela_wire_1655)
    );

    bfr new_Jinkela_buffer_411 (
        .din(new_Jinkela_wire_536),
        .dout(new_Jinkela_wire_537)
    );

    spl2 new_Jinkela_splitter_152 (
        .a(_072_),
        .b(new_Jinkela_wire_1331),
        .c(new_Jinkela_wire_1332)
    );

    bfr new_Jinkela_buffer_1053 (
        .din(new_Jinkela_wire_1646),
        .dout(new_Jinkela_wire_1647)
    );

    bfr new_Jinkela_buffer_933 (
        .din(new_Jinkela_wire_1322),
        .dout(new_Jinkela_wire_1323)
    );

    bfr new_Jinkela_buffer_394 (
        .din(new_Jinkela_wire_511),
        .dout(new_Jinkela_wire_512)
    );

    spl2 new_Jinkela_splitter_242 (
        .a(_299_),
        .b(new_Jinkela_wire_1658),
        .c(new_Jinkela_wire_1659)
    );

    bfr new_Jinkela_buffer_434 (
        .din(new_Jinkela_wire_567),
        .dout(new_Jinkela_wire_568)
    );

    bfr new_Jinkela_buffer_934 (
        .din(new_Jinkela_wire_1323),
        .dout(new_Jinkela_wire_1324)
    );

    bfr new_Jinkela_buffer_1054 (
        .din(new_Jinkela_wire_1647),
        .dout(new_Jinkela_wire_1648)
    );

    bfr new_Jinkela_buffer_395 (
        .din(new_Jinkela_wire_512),
        .dout(new_Jinkela_wire_513)
    );

    spl4L new_Jinkela_splitter_155 (
        .a(_249_),
        .d(new_Jinkela_wire_1338),
        .e(new_Jinkela_wire_1339),
        .b(new_Jinkela_wire_1340),
        .c(new_Jinkela_wire_1341)
    );

    spl2 new_Jinkela_splitter_241 (
        .a(_063_),
        .b(new_Jinkela_wire_1656),
        .c(new_Jinkela_wire_1657)
    );

    bfr new_Jinkela_buffer_412 (
        .din(new_Jinkela_wire_537),
        .dout(new_Jinkela_wire_538)
    );

    bfr new_Jinkela_buffer_935 (
        .din(new_Jinkela_wire_1324),
        .dout(new_Jinkela_wire_1325)
    );

    bfr new_Jinkela_buffer_1055 (
        .din(new_Jinkela_wire_1648),
        .dout(new_Jinkela_wire_1649)
    );

    bfr new_Jinkela_buffer_396 (
        .din(new_Jinkela_wire_513),
        .dout(new_Jinkela_wire_514)
    );

    spl3L new_Jinkela_splitter_153 (
        .a(_110_),
        .d(new_Jinkela_wire_1333),
        .b(new_Jinkela_wire_1334),
        .c(new_Jinkela_wire_1335)
    );

    spl4L new_Jinkela_splitter_55 (
        .a(new_Jinkela_wire_631),
        .d(new_Jinkela_wire_632),
        .e(new_Jinkela_wire_633),
        .b(new_Jinkela_wire_634),
        .c(new_Jinkela_wire_635)
    );

    spl2 new_Jinkela_splitter_150 (
        .a(new_Jinkela_wire_1325),
        .b(new_Jinkela_wire_1326),
        .c(new_Jinkela_wire_1327)
    );

    bfr new_Jinkela_buffer_1056 (
        .din(new_Jinkela_wire_1649),
        .dout(new_Jinkela_wire_1650)
    );

    spl2 new_Jinkela_splitter_57 (
        .a(N105),
        .b(new_Jinkela_wire_663),
        .c(new_Jinkela_wire_665)
    );

    bfr new_Jinkela_buffer_397 (
        .din(new_Jinkela_wire_514),
        .dout(new_Jinkela_wire_515)
    );

    spl2 new_Jinkela_splitter_160 (
        .a(_302_),
        .b(new_Jinkela_wire_1368),
        .c(new_Jinkela_wire_1369)
    );

    bfr new_Jinkela_buffer_1058 (
        .din(_172_),
        .dout(new_Jinkela_wire_1660)
    );

    spl2 new_Jinkela_splitter_154 (
        .a(new_Jinkela_wire_1335),
        .b(new_Jinkela_wire_1336),
        .c(new_Jinkela_wire_1337)
    );

    spl2 new_Jinkela_splitter_244 (
        .a(_248_),
        .b(new_Jinkela_wire_1663),
        .c(new_Jinkela_wire_1664)
    );

    bfr new_Jinkela_buffer_413 (
        .din(new_Jinkela_wire_538),
        .dout(new_Jinkela_wire_539)
    );

    bfr new_Jinkela_buffer_937 (
        .din(_180_),
        .dout(new_Jinkela_wire_1342)
    );

    spl2 new_Jinkela_splitter_243 (
        .a(_192_),
        .b(new_Jinkela_wire_1661),
        .c(new_Jinkela_wire_1662)
    );

    bfr new_Jinkela_buffer_398 (
        .din(new_Jinkela_wire_515),
        .dout(new_Jinkela_wire_516)
    );

    spl2 new_Jinkela_splitter_156 (
        .a(new_Jinkela_wire_1342),
        .b(new_Jinkela_wire_1343),
        .c(new_Jinkela_wire_1344)
    );

    bfr new_Jinkela_buffer_435 (
        .din(new_Jinkela_wire_568),
        .dout(new_Jinkela_wire_569)
    );

    bfr new_Jinkela_buffer_938 (
        .din(new_net_707),
        .dout(new_Jinkela_wire_1345)
    );

    spl2 new_Jinkela_splitter_245 (
        .a(_324_),
        .b(new_Jinkela_wire_1665),
        .c(new_Jinkela_wire_1666)
    );

    bfr new_Jinkela_buffer_399 (
        .din(new_Jinkela_wire_516),
        .dout(new_Jinkela_wire_517)
    );

    spl2 new_Jinkela_splitter_246 (
        .a(_257_),
        .b(new_Jinkela_wire_1667),
        .c(new_Jinkela_wire_1668)
    );

    spl4L new_Jinkela_splitter_157 (
        .a(_145_),
        .d(new_Jinkela_wire_1346),
        .e(new_Jinkela_wire_1347),
        .b(new_Jinkela_wire_1348),
        .c(new_Jinkela_wire_1349)
    );

    spl2 new_Jinkela_splitter_248 (
        .a(_077_),
        .b(new_Jinkela_wire_1671),
        .c(new_Jinkela_wire_1672)
    );

    bfr new_Jinkela_buffer_414 (
        .din(new_Jinkela_wire_539),
        .dout(new_Jinkela_wire_540)
    );

    spl2 new_Jinkela_splitter_247 (
        .a(_315_),
        .b(new_Jinkela_wire_1669),
        .c(new_Jinkela_wire_1670)
    );

    bfr new_Jinkela_buffer_950 (
        .din(_233_),
        .dout(new_Jinkela_wire_1365)
    );

    bfr new_Jinkela_buffer_587 (
        .din(new_Jinkela_wire_760),
        .dout(new_Jinkela_wire_761)
    );

    or_bb _643_ (
        .a(new_Jinkela_wire_1341),
        .b(new_Jinkela_wire_1228),
        .c(_250_)
    );

    bfr new_Jinkela_buffer_624 (
        .din(new_Jinkela_wire_813),
        .dout(new_Jinkela_wire_814)
    );

    or_bi _644_ (
        .a(new_Jinkela_wire_66),
        .b(new_Jinkela_wire_1151),
        .c(_251_)
    );

    bfr new_Jinkela_buffer_588 (
        .din(new_Jinkela_wire_761),
        .dout(new_Jinkela_wire_762)
    );

    and_bi _645_ (
        .a(new_Jinkela_wire_67),
        .b(new_Jinkela_wire_1150),
        .c(_252_)
    );

    bfr new_Jinkela_buffer_604 (
        .din(new_Jinkela_wire_785),
        .dout(new_Jinkela_wire_786)
    );

    and_bi _646_ (
        .a(_251_),
        .b(_252_),
        .c(new_net_707)
    );

    bfr new_Jinkela_buffer_589 (
        .din(new_Jinkela_wire_762),
        .dout(new_Jinkela_wire_763)
    );

    or_bb _647_ (
        .a(new_Jinkela_wire_1663),
        .b(new_Jinkela_wire_1213),
        .c(_253_)
    );

    or_bb _648_ (
        .a(new_Jinkela_wire_1444),
        .b(new_Jinkela_wire_1229),
        .c(_254_)
    );

    bfr new_Jinkela_buffer_590 (
        .din(new_Jinkela_wire_763),
        .dout(new_Jinkela_wire_764)
    );

    and_bi _649_ (
        .a(new_Jinkela_wire_1313),
        .b(new_Jinkela_wire_662),
        .c(_255_)
    );

    bfr new_Jinkela_buffer_605 (
        .din(new_Jinkela_wire_786),
        .dout(new_Jinkela_wire_787)
    );

    and_bi _650_ (
        .a(new_Jinkela_wire_661),
        .b(new_Jinkela_wire_1312),
        .c(_256_)
    );

    spl2 new_Jinkela_splitter_65 (
        .a(new_Jinkela_wire_764),
        .b(new_Jinkela_wire_765),
        .c(new_Jinkela_wire_766)
    );

    and_ii _651_ (
        .a(_256_),
        .b(_255_),
        .c(new_net_715)
    );

    bfr new_Jinkela_buffer_606 (
        .din(new_Jinkela_wire_787),
        .dout(new_Jinkela_wire_788)
    );

    or_bb _652_ (
        .a(new_Jinkela_wire_1340),
        .b(new_Jinkela_wire_1204),
        .c(_257_)
    );

    bfr new_Jinkela_buffer_625 (
        .din(new_Jinkela_wire_814),
        .dout(new_Jinkela_wire_815)
    );

    and_bi _653_ (
        .a(new_Jinkela_wire_1668),
        .b(new_Jinkela_wire_524),
        .c(_258_)
    );

    bfr new_Jinkela_buffer_648 (
        .din(new_Jinkela_wire_845),
        .dout(new_Jinkela_wire_846)
    );

    and_bi _654_ (
        .a(new_Jinkela_wire_523),
        .b(new_Jinkela_wire_1667),
        .c(_259_)
    );

    bfr new_Jinkela_buffer_674 (
        .din(new_Jinkela_wire_874),
        .dout(new_Jinkela_wire_875)
    );

    bfr new_Jinkela_buffer_607 (
        .din(new_Jinkela_wire_788),
        .dout(new_Jinkela_wire_789)
    );

    and_ii _655_ (
        .a(_259_),
        .b(_258_),
        .c(new_net_691)
    );

    bfr new_Jinkela_buffer_626 (
        .din(new_Jinkela_wire_815),
        .dout(new_Jinkela_wire_816)
    );

    or_bb _656_ (
        .a(new_Jinkela_wire_1443),
        .b(new_Jinkela_wire_1205),
        .c(_260_)
    );

    bfr new_Jinkela_buffer_608 (
        .din(new_Jinkela_wire_789),
        .dout(new_Jinkela_wire_790)
    );

    and_bi _657_ (
        .a(new_Jinkela_wire_1296),
        .b(new_Jinkela_wire_490),
        .c(_261_)
    );

    spl2 new_Jinkela_splitter_81 (
        .a(N121),
        .b(new_Jinkela_wire_943),
        .c(new_Jinkela_wire_945)
    );

    and_bi _658_ (
        .a(new_Jinkela_wire_489),
        .b(new_Jinkela_wire_1295),
        .c(_262_)
    );

    bfr new_Jinkela_buffer_675 (
        .din(new_Jinkela_wire_880),
        .dout(new_Jinkela_wire_881)
    );

    bfr new_Jinkela_buffer_609 (
        .din(new_Jinkela_wire_790),
        .dout(new_Jinkela_wire_791)
    );

    and_ii _659_ (
        .a(_262_),
        .b(_261_),
        .c(new_net_693)
    );

    bfr new_Jinkela_buffer_627 (
        .din(new_Jinkela_wire_816),
        .dout(new_Jinkela_wire_817)
    );

    or_bi _660_ (
        .a(new_Jinkela_wire_1339),
        .b(new_Jinkela_wire_1273),
        .c(_263_)
    );

    bfr new_Jinkela_buffer_610 (
        .din(new_Jinkela_wire_791),
        .dout(new_Jinkela_wire_792)
    );

    and_bi _661_ (
        .a(new_Jinkela_wire_976),
        .b(new_Jinkela_wire_1277),
        .c(_264_)
    );

    bfr new_Jinkela_buffer_649 (
        .din(new_Jinkela_wire_846),
        .dout(new_Jinkela_wire_847)
    );

    and_bi _662_ (
        .a(new_Jinkela_wire_1276),
        .b(new_Jinkela_wire_975),
        .c(_265_)
    );

    bfr new_Jinkela_buffer_611 (
        .din(new_Jinkela_wire_792),
        .dout(new_Jinkela_wire_793)
    );

    and_ii _663_ (
        .a(_265_),
        .b(_264_),
        .c(new_net_687)
    );

    bfr new_Jinkela_buffer_628 (
        .din(new_Jinkela_wire_817),
        .dout(new_Jinkela_wire_818)
    );

    or_bi _664_ (
        .a(new_Jinkela_wire_1442),
        .b(new_Jinkela_wire_1274),
        .c(_266_)
    );

    bfr new_Jinkela_buffer_612 (
        .din(new_Jinkela_wire_793),
        .dout(new_Jinkela_wire_794)
    );

    and_bi _665_ (
        .a(new_Jinkela_wire_804),
        .b(new_Jinkela_wire_1625),
        .c(_267_)
    );

    and_bi _666_ (
        .a(new_Jinkela_wire_1624),
        .b(new_Jinkela_wire_803),
        .c(_268_)
    );

    bfr new_Jinkela_buffer_613 (
        .din(new_Jinkela_wire_794),
        .dout(new_Jinkela_wire_795)
    );

    and_ii _667_ (
        .a(_268_),
        .b(_267_),
        .c(new_net_701)
    );

    bfr new_Jinkela_buffer_629 (
        .din(new_Jinkela_wire_818),
        .dout(new_Jinkela_wire_819)
    );

    or_bi _668_ (
        .a(new_Jinkela_wire_1338),
        .b(new_Jinkela_wire_1466),
        .c(_269_)
    );

    bfr new_Jinkela_buffer_614 (
        .din(new_Jinkela_wire_795),
        .dout(new_Jinkela_wire_796)
    );

    or_bi _669_ (
        .a(new_Jinkela_wire_837),
        .b(new_Jinkela_wire_1435),
        .c(_270_)
    );

    bfr new_Jinkela_buffer_650 (
        .din(new_Jinkela_wire_847),
        .dout(new_Jinkela_wire_848)
    );

    and_bi _670_ (
        .a(new_Jinkela_wire_838),
        .b(new_Jinkela_wire_1434),
        .c(_271_)
    );

    bfr new_Jinkela_buffer_615 (
        .din(new_Jinkela_wire_796),
        .dout(new_Jinkela_wire_797)
    );

    and_bi _671_ (
        .a(_270_),
        .b(_271_),
        .c(new_net_713)
    );

    bfr new_Jinkela_buffer_630 (
        .din(new_Jinkela_wire_819),
        .dout(new_Jinkela_wire_820)
    );

    or_bi _672_ (
        .a(new_Jinkela_wire_1441),
        .b(new_Jinkela_wire_1465),
        .c(_272_)
    );

    bfr new_Jinkela_buffer_616 (
        .din(new_Jinkela_wire_797),
        .dout(new_Jinkela_wire_798)
    );

    or_bi _673_ (
        .a(new_Jinkela_wire_276),
        .b(new_Jinkela_wire_1614),
        .c(_273_)
    );

    and_bi _674_ (
        .a(new_Jinkela_wire_275),
        .b(new_Jinkela_wire_1613),
        .c(_274_)
    );

    spl4L new_Jinkela_splitter_82 (
        .a(new_Jinkela_wire_945),
        .d(new_Jinkela_wire_946),
        .e(new_Jinkela_wire_947),
        .b(new_Jinkela_wire_948),
        .c(new_Jinkela_wire_949)
    );

    bfr new_Jinkela_buffer_617 (
        .din(new_Jinkela_wire_798),
        .dout(new_Jinkela_wire_799)
    );

    and_bi _675_ (
        .a(_273_),
        .b(_274_),
        .c(new_net_711)
    );

    bfr new_Jinkela_buffer_631 (
        .din(new_Jinkela_wire_820),
        .dout(new_Jinkela_wire_821)
    );

    or_bb _676_ (
        .a(new_Jinkela_wire_1255),
        .b(new_Jinkela_wire_1422),
        .c(_275_)
    );

    bfr new_Jinkela_buffer_618 (
        .din(new_Jinkela_wire_799),
        .dout(new_Jinkela_wire_800)
    );

    or_bb _677_ (
        .a(new_Jinkela_wire_1309),
        .b(new_Jinkela_wire_1226),
        .c(_276_)
    );

    bfr new_Jinkela_buffer_651 (
        .din(new_Jinkela_wire_848),
        .dout(new_Jinkela_wire_849)
    );

    and_bi _678_ (
        .a(new_Jinkela_wire_1520),
        .b(new_Jinkela_wire_32),
        .c(_277_)
    );

    bfr new_Jinkela_buffer_619 (
        .din(new_Jinkela_wire_800),
        .dout(new_Jinkela_wire_801)
    );

    and_bi _679_ (
        .a(new_Jinkela_wire_33),
        .b(new_Jinkela_wire_1519),
        .c(_278_)
    );

    bfr new_Jinkela_buffer_632 (
        .din(new_Jinkela_wire_821),
        .dout(new_Jinkela_wire_822)
    );

    and_ii _680_ (
        .a(_278_),
        .b(_277_),
        .c(new_net_695)
    );

    bfr new_Jinkela_buffer_620 (
        .din(new_Jinkela_wire_801),
        .dout(new_Jinkela_wire_802)
    );

    or_bb _681_ (
        .a(new_Jinkela_wire_1306),
        .b(new_Jinkela_wire_1206),
        .c(_279_)
    );

    spl4L new_Jinkela_splitter_79 (
        .a(new_Jinkela_wire_910),
        .d(new_Jinkela_wire_911),
        .e(new_Jinkela_wire_912),
        .b(new_Jinkela_wire_913),
        .c(new_Jinkela_wire_914)
    );

    and_bi _682_ (
        .a(new_Jinkela_wire_1166),
        .b(new_Jinkela_wire_628),
        .c(_280_)
    );

    spl2 new_Jinkela_splitter_68 (
        .a(new_Jinkela_wire_802),
        .b(new_Jinkela_wire_803),
        .c(new_Jinkela_wire_804)
    );

    and_bi _683_ (
        .a(new_Jinkela_wire_627),
        .b(new_Jinkela_wire_1165),
        .c(_281_)
    );

    bfr new_Jinkela_buffer_633 (
        .din(new_Jinkela_wire_822),
        .dout(new_Jinkela_wire_823)
    );

    and_ii _684_ (
        .a(_281_),
        .b(_280_),
        .c(new_net_705)
    );

    bfr new_Jinkela_buffer_194 (
        .din(new_Jinkela_wire_255),
        .dout(new_Jinkela_wire_256)
    );

    bfr new_Jinkela_buffer_177 (
        .din(new_Jinkela_wire_230),
        .dout(new_Jinkela_wire_231)
    );

    spl2 new_Jinkela_splitter_33 (
        .a(N45),
        .b(new_Jinkela_wire_383),
        .c(new_Jinkela_wire_385)
    );

    bfr new_Jinkela_buffer_178 (
        .din(new_Jinkela_wire_231),
        .dout(new_Jinkela_wire_232)
    );

    bfr new_Jinkela_buffer_195 (
        .din(new_Jinkela_wire_256),
        .dout(new_Jinkela_wire_257)
    );

    bfr new_Jinkela_buffer_179 (
        .din(new_Jinkela_wire_232),
        .dout(new_Jinkela_wire_233)
    );

    bfr new_Jinkela_buffer_216 (
        .din(new_Jinkela_wire_285),
        .dout(new_Jinkela_wire_286)
    );

    bfr new_Jinkela_buffer_180 (
        .din(new_Jinkela_wire_233),
        .dout(new_Jinkela_wire_234)
    );

    bfr new_Jinkela_buffer_196 (
        .din(new_Jinkela_wire_257),
        .dout(new_Jinkela_wire_258)
    );

    bfr new_Jinkela_buffer_181 (
        .din(new_Jinkela_wire_234),
        .dout(new_Jinkela_wire_235)
    );

    bfr new_Jinkela_buffer_182 (
        .din(new_Jinkela_wire_235),
        .dout(new_Jinkela_wire_236)
    );

    bfr new_Jinkela_buffer_197 (
        .din(new_Jinkela_wire_258),
        .dout(new_Jinkela_wire_259)
    );

    bfr new_Jinkela_buffer_183 (
        .din(new_Jinkela_wire_236),
        .dout(new_Jinkela_wire_237)
    );

    bfr new_Jinkela_buffer_217 (
        .din(new_Jinkela_wire_286),
        .dout(new_Jinkela_wire_287)
    );

    bfr new_Jinkela_buffer_184 (
        .din(new_Jinkela_wire_237),
        .dout(new_Jinkela_wire_238)
    );

    bfr new_Jinkela_buffer_198 (
        .din(new_Jinkela_wire_259),
        .dout(new_Jinkela_wire_260)
    );

    bfr new_Jinkela_buffer_185 (
        .din(new_Jinkela_wire_238),
        .dout(new_Jinkela_wire_239)
    );

    bfr new_Jinkela_buffer_242 (
        .din(new_Jinkela_wire_314),
        .dout(new_Jinkela_wire_315)
    );

    spl4L new_Jinkela_splitter_28 (
        .a(new_Jinkela_wire_316),
        .d(new_Jinkela_wire_317),
        .e(new_Jinkela_wire_318),
        .b(new_Jinkela_wire_319),
        .c(new_Jinkela_wire_320)
    );

    bfr new_Jinkela_buffer_186 (
        .din(new_Jinkela_wire_239),
        .dout(new_Jinkela_wire_240)
    );

    bfr new_Jinkela_buffer_199 (
        .din(new_Jinkela_wire_260),
        .dout(new_Jinkela_wire_261)
    );

    spl2 new_Jinkela_splitter_20 (
        .a(new_Jinkela_wire_240),
        .b(new_Jinkela_wire_241),
        .c(new_Jinkela_wire_242)
    );

    bfr new_Jinkela_buffer_200 (
        .din(new_Jinkela_wire_261),
        .dout(new_Jinkela_wire_262)
    );

    bfr new_Jinkela_buffer_218 (
        .din(new_Jinkela_wire_287),
        .dout(new_Jinkela_wire_288)
    );

    bfr new_Jinkela_buffer_243 (
        .din(new_Jinkela_wire_320),
        .dout(new_Jinkela_wire_321)
    );

    bfr new_Jinkela_buffer_201 (
        .din(new_Jinkela_wire_262),
        .dout(new_Jinkela_wire_263)
    );

    bfr new_Jinkela_buffer_219 (
        .din(new_Jinkela_wire_288),
        .dout(new_Jinkela_wire_289)
    );

    bfr new_Jinkela_buffer_202 (
        .din(new_Jinkela_wire_263),
        .dout(new_Jinkela_wire_264)
    );

    bfr new_Jinkela_buffer_203 (
        .din(new_Jinkela_wire_264),
        .dout(new_Jinkela_wire_265)
    );

    bfr new_Jinkela_buffer_220 (
        .din(new_Jinkela_wire_289),
        .dout(new_Jinkela_wire_290)
    );

    bfr new_Jinkela_buffer_204 (
        .din(new_Jinkela_wire_265),
        .dout(new_Jinkela_wire_266)
    );

    bfr new_Jinkela_buffer_269 (
        .din(new_Jinkela_wire_349),
        .dout(new_Jinkela_wire_350)
    );

    bfr new_Jinkela_buffer_205 (
        .din(new_Jinkela_wire_266),
        .dout(new_Jinkela_wire_267)
    );

    bfr new_Jinkela_buffer_221 (
        .din(new_Jinkela_wire_290),
        .dout(new_Jinkela_wire_291)
    );

    bfr new_Jinkela_buffer_206 (
        .din(new_Jinkela_wire_267),
        .dout(new_Jinkela_wire_268)
    );

    bfr new_Jinkela_buffer_244 (
        .din(new_Jinkela_wire_321),
        .dout(new_Jinkela_wire_322)
    );

    bfr new_Jinkela_buffer_207 (
        .din(new_Jinkela_wire_268),
        .dout(new_Jinkela_wire_269)
    );

    bfr new_Jinkela_buffer_222 (
        .din(new_Jinkela_wire_291),
        .dout(new_Jinkela_wire_292)
    );

    bfr new_Jinkela_buffer_208 (
        .din(new_Jinkela_wire_269),
        .dout(new_Jinkela_wire_270)
    );

    spl4L new_Jinkela_splitter_34 (
        .a(new_Jinkela_wire_385),
        .d(new_Jinkela_wire_386),
        .e(new_Jinkela_wire_387),
        .b(new_Jinkela_wire_388),
        .c(new_Jinkela_wire_389)
    );

    bfr new_Jinkela_buffer_322 (
        .din(N132),
        .dout(new_Jinkela_wire_418)
    );

    bfr new_Jinkela_buffer_209 (
        .din(new_Jinkela_wire_270),
        .dout(new_Jinkela_wire_271)
    );

    inv _475_ (
        .din(new_Jinkela_wire_1612),
        .dout(_087_)
    );

    or_bi _476_ (
        .a(new_Jinkela_wire_1652),
        .b(new_Jinkela_wire_1231),
        .c(_088_)
    );

    and_bi _477_ (
        .a(new_Jinkela_wire_564),
        .b(new_Jinkela_wire_211),
        .c(_089_)
    );

    and_bi _478_ (
        .a(new_Jinkela_wire_209),
        .b(new_Jinkela_wire_565),
        .c(_090_)
    );

    or_bb _479_ (
        .a(_090_),
        .b(_089_),
        .c(_091_)
    );

    or_ii _480_ (
        .a(new_Jinkela_wire_1051),
        .b(new_Jinkela_wire_1095),
        .c(_092_)
    );

    or_bi _481_ (
        .a(new_Jinkela_wire_178),
        .b(new_Jinkela_wire_281),
        .c(_093_)
    );

    and_bi _482_ (
        .a(new_Jinkela_wire_177),
        .b(new_Jinkela_wire_278),
        .c(_094_)
    );

    and_bi _483_ (
        .a(_093_),
        .b(_094_),
        .c(_095_)
    );

    and_bi _484_ (
        .a(new_Jinkela_wire_1639),
        .b(new_Jinkela_wire_1409),
        .c(_096_)
    );

    and_bi _485_ (
        .a(new_Jinkela_wire_1408),
        .b(new_Jinkela_wire_1638),
        .c(_097_)
    );

    or_bb _486_ (
        .a(_097_),
        .b(_096_),
        .c(_098_)
    );

    or_bb _487_ (
        .a(new_Jinkela_wire_1495),
        .b(new_Jinkela_wire_1440),
        .c(_099_)
    );

    and_bb _488_ (
        .a(new_Jinkela_wire_1494),
        .b(new_Jinkela_wire_1439),
        .c(_100_)
    );

    and_bi _489_ (
        .a(_099_),
        .b(_100_),
        .c(_101_)
    );

    or_bb _490_ (
        .a(new_Jinkela_wire_247),
        .b(new_Jinkela_wire_775),
        .c(_102_)
    );

    and_bb _491_ (
        .a(new_Jinkela_wire_248),
        .b(new_Jinkela_wire_776),
        .c(_103_)
    );

    and_bi _492_ (
        .a(_102_),
        .b(_103_),
        .c(_104_)
    );

    or_bi _493_ (
        .a(new_Jinkela_wire_458),
        .b(new_Jinkela_wire_633),
        .c(_105_)
    );

    and_bi _494_ (
        .a(new_Jinkela_wire_460),
        .b(new_Jinkela_wire_632),
        .c(_106_)
    );

    or_bi _495_ (
        .a(_106_),
        .b(_105_),
        .c(_107_)
    );

    or_bi _496_ (
        .a(new_Jinkela_wire_1387),
        .b(new_Jinkela_wire_1389),
        .c(_108_)
    );

    and_bi _497_ (
        .a(new_Jinkela_wire_1386),
        .b(new_Jinkela_wire_1388),
        .c(_109_)
    );

    and_bi _498_ (
        .a(_108_),
        .b(_109_),
        .c(_110_)
    );

    or_bb _499_ (
        .a(new_Jinkela_wire_1334),
        .b(new_Jinkela_wire_1675),
        .c(_111_)
    );

    and_bb _500_ (
        .a(new_Jinkela_wire_1333),
        .b(new_Jinkela_wire_1673),
        .c(_112_)
    );

    and_bi _501_ (
        .a(_111_),
        .b(_112_),
        .c(_113_)
    );

    and_bi _502_ (
        .a(new_Jinkela_wire_1377),
        .b(new_Jinkela_wire_1159),
        .c(_114_)
    );

    and_bi _503_ (
        .a(new_Jinkela_wire_1158),
        .b(new_Jinkela_wire_1376),
        .c(_115_)
    );

    or_bb _504_ (
        .a(_115_),
        .b(_114_),
        .c(_116_)
    );

    and_bi _505_ (
        .a(new_Jinkela_wire_1058),
        .b(new_Jinkela_wire_843),
        .c(_117_)
    );

    and_bi _506_ (
        .a(new_Jinkela_wire_840),
        .b(new_Jinkela_wire_1062),
        .c(_118_)
    );

    or_bb _507_ (
        .a(_118_),
        .b(_117_),
        .c(_119_)
    );

    or_ii _508_ (
        .a(new_Jinkela_wire_768),
        .b(new_Jinkela_wire_1049),
        .c(_120_)
    );

    or_bi _509_ (
        .a(new_Jinkela_wire_530),
        .b(new_Jinkela_wire_736),
        .c(_121_)
    );

    and_bi _510_ (
        .a(new_Jinkela_wire_526),
        .b(new_Jinkela_wire_735),
        .c(_122_)
    );

    and_bi _511_ (
        .a(_121_),
        .b(_122_),
        .c(_123_)
    );

    and_bi _512_ (
        .a(new_Jinkela_wire_1693),
        .b(new_Jinkela_wire_1286),
        .c(_124_)
    );

    and_bi _513_ (
        .a(new_Jinkela_wire_1285),
        .b(new_Jinkela_wire_1692),
        .c(_125_)
    );

    or_bb _514_ (
        .a(_125_),
        .b(_124_),
        .c(_126_)
    );

    or_bb _515_ (
        .a(new_Jinkela_wire_1315),
        .b(new_Jinkela_wire_1171),
        .c(_127_)
    );

    and_bb _516_ (
        .a(new_Jinkela_wire_1314),
        .b(new_Jinkela_wire_1170),
        .c(_128_)
    );

    bfr new_Jinkela_buffer_400 (
        .din(new_Jinkela_wire_517),
        .dout(new_Jinkela_wire_518)
    );

    bfr new_Jinkela_buffer_401 (
        .din(new_Jinkela_wire_518),
        .dout(new_Jinkela_wire_519)
    );

    bfr new_Jinkela_buffer_415 (
        .din(new_Jinkela_wire_540),
        .dout(new_Jinkela_wire_541)
    );

    bfr new_Jinkela_buffer_402 (
        .din(new_Jinkela_wire_519),
        .dout(new_Jinkela_wire_520)
    );

    bfr new_Jinkela_buffer_436 (
        .din(new_Jinkela_wire_569),
        .dout(new_Jinkela_wire_570)
    );

    bfr new_Jinkela_buffer_403 (
        .din(new_Jinkela_wire_520),
        .dout(new_Jinkela_wire_521)
    );

    bfr new_Jinkela_buffer_416 (
        .din(new_Jinkela_wire_541),
        .dout(new_Jinkela_wire_542)
    );

    bfr new_Jinkela_buffer_404 (
        .din(new_Jinkela_wire_521),
        .dout(new_Jinkela_wire_522)
    );

    bfr new_Jinkela_buffer_460 (
        .din(new_Jinkela_wire_601),
        .dout(new_Jinkela_wire_602)
    );

    bfr new_Jinkela_buffer_485 (
        .din(new_Jinkela_wire_629),
        .dout(new_Jinkela_wire_630)
    );

    spl2 new_Jinkela_splitter_44 (
        .a(new_Jinkela_wire_522),
        .b(new_Jinkela_wire_523),
        .c(new_Jinkela_wire_524)
    );

    bfr new_Jinkela_buffer_437 (
        .din(new_Jinkela_wire_570),
        .dout(new_Jinkela_wire_571)
    );

    bfr new_Jinkela_buffer_417 (
        .din(new_Jinkela_wire_542),
        .dout(new_Jinkela_wire_543)
    );

    bfr new_Jinkela_buffer_418 (
        .din(new_Jinkela_wire_543),
        .dout(new_Jinkela_wire_544)
    );

    spl2 new_Jinkela_splitter_60 (
        .a(N41),
        .b(new_Jinkela_wire_697),
        .c(new_Jinkela_wire_699)
    );

    bfr new_Jinkela_buffer_486 (
        .din(new_Jinkela_wire_635),
        .dout(new_Jinkela_wire_636)
    );

    bfr new_Jinkela_buffer_419 (
        .din(new_Jinkela_wire_544),
        .dout(new_Jinkela_wire_545)
    );

    bfr new_Jinkela_buffer_438 (
        .din(new_Jinkela_wire_571),
        .dout(new_Jinkela_wire_572)
    );

    bfr new_Jinkela_buffer_420 (
        .din(new_Jinkela_wire_545),
        .dout(new_Jinkela_wire_546)
    );

    bfr new_Jinkela_buffer_461 (
        .din(new_Jinkela_wire_602),
        .dout(new_Jinkela_wire_603)
    );

    bfr new_Jinkela_buffer_421 (
        .din(new_Jinkela_wire_546),
        .dout(new_Jinkela_wire_547)
    );

    bfr new_Jinkela_buffer_439 (
        .din(new_Jinkela_wire_572),
        .dout(new_Jinkela_wire_573)
    );

    bfr new_Jinkela_buffer_422 (
        .din(new_Jinkela_wire_547),
        .dout(new_Jinkela_wire_548)
    );

    bfr new_Jinkela_buffer_423 (
        .din(new_Jinkela_wire_548),
        .dout(new_Jinkela_wire_549)
    );

    bfr new_Jinkela_buffer_440 (
        .din(new_Jinkela_wire_573),
        .dout(new_Jinkela_wire_574)
    );

    bfr new_Jinkela_buffer_424 (
        .din(new_Jinkela_wire_549),
        .dout(new_Jinkela_wire_550)
    );

    bfr new_Jinkela_buffer_462 (
        .din(new_Jinkela_wire_603),
        .dout(new_Jinkela_wire_604)
    );

    bfr new_Jinkela_buffer_425 (
        .din(new_Jinkela_wire_550),
        .dout(new_Jinkela_wire_551)
    );

    bfr new_Jinkela_buffer_441 (
        .din(new_Jinkela_wire_574),
        .dout(new_Jinkela_wire_575)
    );

    bfr new_Jinkela_buffer_426 (
        .din(new_Jinkela_wire_551),
        .dout(new_Jinkela_wire_552)
    );

    spl4L new_Jinkela_splitter_61 (
        .a(new_Jinkela_wire_699),
        .d(new_Jinkela_wire_700),
        .e(new_Jinkela_wire_701),
        .b(new_Jinkela_wire_702),
        .c(new_Jinkela_wire_703)
    );

    bfr new_Jinkela_buffer_427 (
        .din(new_Jinkela_wire_552),
        .dout(new_Jinkela_wire_553)
    );

    bfr new_Jinkela_buffer_442 (
        .din(new_Jinkela_wire_575),
        .dout(new_Jinkela_wire_576)
    );

    bfr new_Jinkela_buffer_428 (
        .din(new_Jinkela_wire_553),
        .dout(new_Jinkela_wire_554)
    );

    bfr new_Jinkela_buffer_463 (
        .din(new_Jinkela_wire_604),
        .dout(new_Jinkela_wire_605)
    );

    bfr new_Jinkela_buffer_429 (
        .din(new_Jinkela_wire_554),
        .dout(new_Jinkela_wire_555)
    );

    bfr new_Jinkela_buffer_443 (
        .din(new_Jinkela_wire_576),
        .dout(new_Jinkela_wire_577)
    );

    bfr new_Jinkela_buffer_430 (
        .din(new_Jinkela_wire_555),
        .dout(new_Jinkela_wire_556)
    );

    spl4L new_Jinkela_splitter_58 (
        .a(new_Jinkela_wire_665),
        .d(new_Jinkela_wire_666),
        .e(new_Jinkela_wire_667),
        .b(new_Jinkela_wire_668),
        .c(new_Jinkela_wire_669)
    );

    bfr new_Jinkela_buffer_431 (
        .din(new_Jinkela_wire_556),
        .dout(new_Jinkela_wire_557)
    );

    bfr new_Jinkela_buffer_444 (
        .din(new_Jinkela_wire_577),
        .dout(new_Jinkela_wire_578)
    );

    spl2 new_Jinkela_splitter_47 (
        .a(new_Jinkela_wire_557),
        .b(new_Jinkela_wire_558),
        .c(new_Jinkela_wire_559)
    );

    bfr new_Jinkela_buffer_1 (
        .din(new_Jinkela_wire_6),
        .dout(new_Jinkela_wire_7)
    );

    bfr new_Jinkela_buffer_26 (
        .din(new_Jinkela_wire_34),
        .dout(new_Jinkela_wire_35)
    );

    bfr new_Jinkela_buffer_78 (
        .din(N134),
        .dout(new_Jinkela_wire_102)
    );

    bfr new_Jinkela_buffer_27 (
        .din(new_Jinkela_wire_40),
        .dout(new_Jinkela_wire_41)
    );

    bfr new_Jinkela_buffer_2 (
        .din(new_Jinkela_wire_7),
        .dout(new_Jinkela_wire_8)
    );

    bfr new_Jinkela_buffer_3 (
        .din(new_Jinkela_wire_8),
        .dout(new_Jinkela_wire_9)
    );

    bfr new_Jinkela_buffer_79 (
        .din(new_Jinkela_wire_102),
        .dout(new_Jinkela_wire_103)
    );

    bfr new_Jinkela_buffer_4 (
        .din(new_Jinkela_wire_9),
        .dout(new_Jinkela_wire_10)
    );

    spl4L new_Jinkela_splitter_7 (
        .a(new_Jinkela_wire_70),
        .d(new_Jinkela_wire_71),
        .e(new_Jinkela_wire_72),
        .b(new_Jinkela_wire_73),
        .c(new_Jinkela_wire_74)
    );

    bfr new_Jinkela_buffer_5 (
        .din(new_Jinkela_wire_10),
        .dout(new_Jinkela_wire_11)
    );

    bfr new_Jinkela_buffer_53 (
        .din(new_Jinkela_wire_74),
        .dout(new_Jinkela_wire_75)
    );

    spl2 new_Jinkela_splitter_12 (
        .a(N77),
        .b(new_Jinkela_wire_139),
        .c(new_Jinkela_wire_141)
    );

    bfr new_Jinkela_buffer_6 (
        .din(new_Jinkela_wire_11),
        .dout(new_Jinkela_wire_12)
    );

    bfr new_Jinkela_buffer_28 (
        .din(new_Jinkela_wire_41),
        .dout(new_Jinkela_wire_42)
    );

    bfr new_Jinkela_buffer_7 (
        .din(new_Jinkela_wire_12),
        .dout(new_Jinkela_wire_13)
    );

    bfr new_Jinkela_buffer_8 (
        .din(new_Jinkela_wire_13),
        .dout(new_Jinkela_wire_14)
    );

    bfr new_Jinkela_buffer_29 (
        .din(new_Jinkela_wire_42),
        .dout(new_Jinkela_wire_43)
    );

    bfr new_Jinkela_buffer_9 (
        .din(new_Jinkela_wire_14),
        .dout(new_Jinkela_wire_15)
    );

    spl2 new_Jinkela_splitter_9 (
        .a(N57),
        .b(new_Jinkela_wire_104),
        .c(new_Jinkela_wire_106)
    );

    bfr new_Jinkela_buffer_52 (
        .din(new_Jinkela_wire_68),
        .dout(new_Jinkela_wire_69)
    );

    bfr new_Jinkela_buffer_10 (
        .din(new_Jinkela_wire_15),
        .dout(new_Jinkela_wire_16)
    );

    bfr new_Jinkela_buffer_30 (
        .din(new_Jinkela_wire_43),
        .dout(new_Jinkela_wire_44)
    );

    bfr new_Jinkela_buffer_11 (
        .din(new_Jinkela_wire_16),
        .dout(new_Jinkela_wire_17)
    );

    bfr new_Jinkela_buffer_12 (
        .din(new_Jinkela_wire_17),
        .dout(new_Jinkela_wire_18)
    );

    bfr new_Jinkela_buffer_31 (
        .din(new_Jinkela_wire_44),
        .dout(new_Jinkela_wire_45)
    );

    bfr new_Jinkela_buffer_13 (
        .din(new_Jinkela_wire_18),
        .dout(new_Jinkela_wire_19)
    );

    spl4L new_Jinkela_splitter_13 (
        .a(new_Jinkela_wire_141),
        .d(new_Jinkela_wire_142),
        .e(new_Jinkela_wire_143),
        .b(new_Jinkela_wire_144),
        .c(new_Jinkela_wire_145)
    );

    spl4L new_Jinkela_splitter_10 (
        .a(new_Jinkela_wire_106),
        .d(new_Jinkela_wire_107),
        .e(new_Jinkela_wire_108),
        .b(new_Jinkela_wire_109),
        .c(new_Jinkela_wire_110)
    );

    bfr new_Jinkela_buffer_14 (
        .din(new_Jinkela_wire_19),
        .dout(new_Jinkela_wire_20)
    );

    bfr new_Jinkela_buffer_32 (
        .din(new_Jinkela_wire_45),
        .dout(new_Jinkela_wire_46)
    );

    bfr new_Jinkela_buffer_15 (
        .din(new_Jinkela_wire_20),
        .dout(new_Jinkela_wire_21)
    );

    bfr new_Jinkela_buffer_54 (
        .din(new_Jinkela_wire_75),
        .dout(new_Jinkela_wire_76)
    );

    bfr new_Jinkela_buffer_33 (
        .din(new_Jinkela_wire_46),
        .dout(new_Jinkela_wire_47)
    );

    bfr new_Jinkela_buffer_16 (
        .din(new_Jinkela_wire_21),
        .dout(new_Jinkela_wire_22)
    );

    bfr new_Jinkela_buffer_17 (
        .din(new_Jinkela_wire_22),
        .dout(new_Jinkela_wire_23)
    );

    bfr new_Jinkela_buffer_18 (
        .din(new_Jinkela_wire_23),
        .dout(new_Jinkela_wire_24)
    );

    bfr new_Jinkela_buffer_34 (
        .din(new_Jinkela_wire_47),
        .dout(new_Jinkela_wire_48)
    );

    bfr new_Jinkela_buffer_19 (
        .din(new_Jinkela_wire_24),
        .dout(new_Jinkela_wire_25)
    );

    bfr new_Jinkela_buffer_522 (
        .din(new_Jinkela_wire_679),
        .dout(new_Jinkela_wire_680)
    );

    bfr new_Jinkela_buffer_55 (
        .din(new_Jinkela_wire_76),
        .dout(new_Jinkela_wire_77)
    );

    bfr new_Jinkela_buffer_20 (
        .din(new_Jinkela_wire_25),
        .dout(new_Jinkela_wire_26)
    );

    bfr new_Jinkela_buffer_35 (
        .din(new_Jinkela_wire_48),
        .dout(new_Jinkela_wire_49)
    );

    bfr new_Jinkela_buffer_21 (
        .din(new_Jinkela_wire_26),
        .dout(new_Jinkela_wire_27)
    );

    bfr new_Jinkela_buffer_841 (
        .din(new_Jinkela_wire_1104),
        .dout(new_Jinkela_wire_1105)
    );

    bfr new_Jinkela_buffer_820 (
        .din(new_Jinkela_wire_1075),
        .dout(new_Jinkela_wire_1076)
    );

    spl2 new_Jinkela_splitter_101 (
        .a(_020_),
        .b(new_Jinkela_wire_1139),
        .c(new_Jinkela_wire_1140)
    );

    bfr new_Jinkela_buffer_821 (
        .din(new_Jinkela_wire_1076),
        .dout(new_Jinkela_wire_1077)
    );

    bfr new_Jinkela_buffer_842 (
        .din(new_Jinkela_wire_1105),
        .dout(new_Jinkela_wire_1106)
    );

    bfr new_Jinkela_buffer_822 (
        .din(new_Jinkela_wire_1077),
        .dout(new_Jinkela_wire_1078)
    );

    spl2 new_Jinkela_splitter_102 (
        .a(_166_),
        .b(new_Jinkela_wire_1141),
        .c(new_Jinkela_wire_1142)
    );

    bfr new_Jinkela_buffer_868 (
        .din(new_Jinkela_wire_1137),
        .dout(new_Jinkela_wire_1138)
    );

    bfr new_Jinkela_buffer_823 (
        .din(new_Jinkela_wire_1078),
        .dout(new_Jinkela_wire_1079)
    );

    bfr new_Jinkela_buffer_843 (
        .din(new_Jinkela_wire_1106),
        .dout(new_Jinkela_wire_1107)
    );

    bfr new_Jinkela_buffer_824 (
        .din(new_Jinkela_wire_1079),
        .dout(new_Jinkela_wire_1080)
    );

    spl2 new_Jinkela_splitter_106 (
        .a(_250_),
        .b(new_Jinkela_wire_1150),
        .c(new_Jinkela_wire_1151)
    );

    bfr new_Jinkela_buffer_825 (
        .din(new_Jinkela_wire_1080),
        .dout(new_Jinkela_wire_1081)
    );

    bfr new_Jinkela_buffer_844 (
        .din(new_Jinkela_wire_1107),
        .dout(new_Jinkela_wire_1108)
    );

    bfr new_Jinkela_buffer_826 (
        .din(new_Jinkela_wire_1081),
        .dout(new_Jinkela_wire_1082)
    );

    bfr new_Jinkela_buffer_827 (
        .din(new_Jinkela_wire_1082),
        .dout(new_Jinkela_wire_1083)
    );

    bfr new_Jinkela_buffer_845 (
        .din(new_Jinkela_wire_1108),
        .dout(new_Jinkela_wire_1109)
    );

    bfr new_Jinkela_buffer_828 (
        .din(new_Jinkela_wire_1083),
        .dout(new_Jinkela_wire_1084)
    );

    spl2 new_Jinkela_splitter_103 (
        .a(_305_),
        .b(new_Jinkela_wire_1143),
        .c(new_Jinkela_wire_1144)
    );

    bfr new_Jinkela_buffer_829 (
        .din(new_Jinkela_wire_1084),
        .dout(new_Jinkela_wire_1085)
    );

    bfr new_Jinkela_buffer_846 (
        .din(new_Jinkela_wire_1109),
        .dout(new_Jinkela_wire_1110)
    );

    bfr new_Jinkela_buffer_830 (
        .din(new_Jinkela_wire_1085),
        .dout(new_Jinkela_wire_1086)
    );

    spl3L new_Jinkela_splitter_104 (
        .a(_004_),
        .d(new_Jinkela_wire_1145),
        .b(new_Jinkela_wire_1146),
        .c(new_Jinkela_wire_1147)
    );

    bfr new_Jinkela_buffer_831 (
        .din(new_Jinkela_wire_1086),
        .dout(new_Jinkela_wire_1087)
    );

    bfr new_Jinkela_buffer_847 (
        .din(new_Jinkela_wire_1110),
        .dout(new_Jinkela_wire_1111)
    );

    bfr new_Jinkela_buffer_832 (
        .din(new_Jinkela_wire_1087),
        .dout(new_Jinkela_wire_1088)
    );

    spl2 new_Jinkela_splitter_107 (
        .a(_137_),
        .b(new_Jinkela_wire_1152),
        .c(new_Jinkela_wire_1153)
    );

    bfr new_Jinkela_buffer_833 (
        .din(new_Jinkela_wire_1088),
        .dout(new_Jinkela_wire_1089)
    );

    bfr new_Jinkela_buffer_848 (
        .din(new_Jinkela_wire_1111),
        .dout(new_Jinkela_wire_1112)
    );

    spl2 new_Jinkela_splitter_95 (
        .a(new_Jinkela_wire_1089),
        .b(new_Jinkela_wire_1090),
        .c(new_Jinkela_wire_1091)
    );

    bfr new_Jinkela_buffer_849 (
        .din(new_Jinkela_wire_1112),
        .dout(new_Jinkela_wire_1113)
    );

    spl2 new_Jinkela_splitter_109 (
        .a(_101_),
        .b(new_Jinkela_wire_1158),
        .c(new_Jinkela_wire_1159)
    );

    spl2 new_Jinkela_splitter_105 (
        .a(new_Jinkela_wire_1147),
        .b(new_Jinkela_wire_1148),
        .c(new_Jinkela_wire_1149)
    );

    bfr new_Jinkela_buffer_850 (
        .din(new_Jinkela_wire_1113),
        .dout(new_Jinkela_wire_1114)
    );

    bfr new_Jinkela_buffer_851 (
        .din(new_Jinkela_wire_1114),
        .dout(new_Jinkela_wire_1115)
    );

    spl2 new_Jinkela_splitter_108 (
        .a(_345_),
        .b(new_Jinkela_wire_1154),
        .c(new_Jinkela_wire_1155)
    );

    bfr new_Jinkela_buffer_869 (
        .din(new_net_691),
        .dout(new_Jinkela_wire_1156)
    );

    bfr new_Jinkela_buffer_852 (
        .din(new_Jinkela_wire_1115),
        .dout(new_Jinkela_wire_1116)
    );

    bfr new_Jinkela_buffer_870 (
        .din(new_net_703),
        .dout(new_Jinkela_wire_1157)
    );

    bfr new_Jinkela_buffer_853 (
        .din(new_Jinkela_wire_1116),
        .dout(new_Jinkela_wire_1117)
    );

    bfr new_Jinkela_buffer_871 (
        .din(new_net_699),
        .dout(new_Jinkela_wire_1160)
    );

    bfr new_Jinkela_buffer_854 (
        .din(new_Jinkela_wire_1117),
        .dout(new_Jinkela_wire_1118)
    );

    bfr new_Jinkela_buffer_223 (
        .din(new_Jinkela_wire_292),
        .dout(new_Jinkela_wire_293)
    );

    bfr new_Jinkela_buffer_1059 (
        .din(_175_),
        .dout(new_Jinkela_wire_1681)
    );

    bfr new_Jinkela_buffer_939 (
        .din(new_Jinkela_wire_1349),
        .dout(new_Jinkela_wire_1350)
    );

    bfr new_Jinkela_buffer_210 (
        .din(new_Jinkela_wire_271),
        .dout(new_Jinkela_wire_272)
    );

    spl4L new_Jinkela_splitter_249 (
        .a(_357_),
        .d(new_Jinkela_wire_1673),
        .e(new_Jinkela_wire_1674),
        .b(new_Jinkela_wire_1675),
        .c(new_Jinkela_wire_1676)
    );

    bfr new_Jinkela_buffer_245 (
        .din(new_Jinkela_wire_322),
        .dout(new_Jinkela_wire_323)
    );

    spl2 new_Jinkela_splitter_161 (
        .a(_044_),
        .b(new_Jinkela_wire_1370),
        .c(new_Jinkela_wire_1371)
    );

    spl2 new_Jinkela_splitter_250 (
        .a(_157_),
        .b(new_Jinkela_wire_1677),
        .c(new_Jinkela_wire_1678)
    );

    bfr new_Jinkela_buffer_211 (
        .din(new_Jinkela_wire_272),
        .dout(new_Jinkela_wire_273)
    );

    spl2 new_Jinkela_splitter_159 (
        .a(new_Jinkela_wire_1365),
        .b(new_Jinkela_wire_1366),
        .c(new_Jinkela_wire_1367)
    );

    bfr new_Jinkela_buffer_940 (
        .din(new_Jinkela_wire_1350),
        .dout(new_Jinkela_wire_1351)
    );

    bfr new_Jinkela_buffer_224 (
        .din(new_Jinkela_wire_293),
        .dout(new_Jinkela_wire_294)
    );

    spl2 new_Jinkela_splitter_251 (
        .a(_080_),
        .b(new_Jinkela_wire_1679),
        .c(new_Jinkela_wire_1680)
    );

    bfr new_Jinkela_buffer_1060 (
        .din(new_Jinkela_wire_1681),
        .dout(new_Jinkela_wire_1682)
    );

    bfr new_Jinkela_buffer_212 (
        .din(new_Jinkela_wire_273),
        .dout(new_Jinkela_wire_274)
    );

    spl2 new_Jinkela_splitter_253 (
        .a(_186_),
        .b(new_Jinkela_wire_1686),
        .c(new_Jinkela_wire_1687)
    );

    bfr new_Jinkela_buffer_1061 (
        .din(_163_),
        .dout(new_Jinkela_wire_1683)
    );

    bfr new_Jinkela_buffer_941 (
        .din(new_Jinkela_wire_1351),
        .dout(new_Jinkela_wire_1352)
    );

    spl2 new_Jinkela_splitter_257 (
        .a(_051_),
        .b(new_Jinkela_wire_1694),
        .c(new_Jinkela_wire_1695)
    );

    spl2 new_Jinkela_splitter_162 (
        .a(_136_),
        .b(new_Jinkela_wire_1372),
        .c(new_Jinkela_wire_1373)
    );

    spl2 new_Jinkela_splitter_23 (
        .a(new_Jinkela_wire_274),
        .b(new_Jinkela_wire_275),
        .c(new_Jinkela_wire_276)
    );

    spl2 new_Jinkela_splitter_163 (
        .a(_142_),
        .b(new_Jinkela_wire_1374),
        .c(new_Jinkela_wire_1375)
    );

    spl2 new_Jinkela_splitter_254 (
        .a(_001_),
        .b(new_Jinkela_wire_1688),
        .c(new_Jinkela_wire_1689)
    );

    spl2 new_Jinkela_splitter_252 (
        .a(new_Jinkela_wire_1683),
        .b(new_Jinkela_wire_1684),
        .c(new_Jinkela_wire_1685)
    );

    bfr new_Jinkela_buffer_942 (
        .din(new_Jinkela_wire_1352),
        .dout(new_Jinkela_wire_1353)
    );

    bfr new_Jinkela_buffer_246 (
        .din(new_Jinkela_wire_323),
        .dout(new_Jinkela_wire_324)
    );

    bfr new_Jinkela_buffer_225 (
        .din(new_Jinkela_wire_294),
        .dout(new_Jinkela_wire_295)
    );

    spl2 new_Jinkela_splitter_255 (
        .a(_154_),
        .b(new_Jinkela_wire_1690),
        .c(new_Jinkela_wire_1691)
    );

    bfr new_Jinkela_buffer_943 (
        .din(new_Jinkela_wire_1353),
        .dout(new_Jinkela_wire_1354)
    );

    bfr new_Jinkela_buffer_226 (
        .din(new_Jinkela_wire_295),
        .dout(new_Jinkela_wire_296)
    );

    bfr new_Jinkela_buffer_951 (
        .din(_336_),
        .dout(new_Jinkela_wire_1380)
    );

    bfr new_Jinkela_buffer_270 (
        .din(new_Jinkela_wire_355),
        .dout(new_Jinkela_wire_356)
    );

    spl2 new_Jinkela_splitter_164 (
        .a(_113_),
        .b(new_Jinkela_wire_1376),
        .c(new_Jinkela_wire_1377)
    );

    bfr new_Jinkela_buffer_944 (
        .din(new_Jinkela_wire_1354),
        .dout(new_Jinkela_wire_1355)
    );

    bfr new_Jinkela_buffer_295 (
        .din(new_Jinkela_wire_383),
        .dout(new_Jinkela_wire_384)
    );

    spl2 new_Jinkela_splitter_256 (
        .a(_123_),
        .b(new_Jinkela_wire_1692),
        .c(new_Jinkela_wire_1693)
    );

    bfr new_Jinkela_buffer_227 (
        .din(new_Jinkela_wire_296),
        .dout(new_Jinkela_wire_297)
    );

    spl2 new_Jinkela_splitter_258 (
        .a(new_Jinkela_wire_1696),
        .b(new_Jinkela_wire_1697),
        .c(new_Jinkela_wire_1698)
    );

    bfr new_Jinkela_buffer_247 (
        .din(new_Jinkela_wire_324),
        .dout(new_Jinkela_wire_325)
    );

    bfr new_Jinkela_buffer_1062 (
        .din(_129_),
        .dout(new_Jinkela_wire_1696)
    );

    spl2 new_Jinkela_splitter_260 (
        .a(_221_),
        .b(new_Jinkela_wire_1701),
        .c(new_Jinkela_wire_1702)
    );

    bfr new_Jinkela_buffer_945 (
        .din(new_Jinkela_wire_1355),
        .dout(new_Jinkela_wire_1356)
    );

    bfr new_Jinkela_buffer_228 (
        .din(new_Jinkela_wire_297),
        .dout(new_Jinkela_wire_298)
    );

    spl2 new_Jinkela_splitter_259 (
        .a(_330_),
        .b(new_Jinkela_wire_1699),
        .c(new_Jinkela_wire_1700)
    );

    spl2 new_Jinkela_splitter_165 (
        .a(_078_),
        .b(new_Jinkela_wire_1378),
        .c(new_Jinkela_wire_1379)
    );

    bfr new_Jinkela_buffer_323 (
        .din(new_Jinkela_wire_418),
        .dout(new_Jinkela_wire_419)
    );

    spl2 new_Jinkela_splitter_168 (
        .a(_107_),
        .b(new_Jinkela_wire_1388),
        .c(new_Jinkela_wire_1389)
    );

    bfr new_Jinkela_buffer_946 (
        .din(new_Jinkela_wire_1356),
        .dout(new_Jinkela_wire_1357)
    );

    bfr new_Jinkela_buffer_296 (
        .din(new_Jinkela_wire_389),
        .dout(new_Jinkela_wire_390)
    );

    bfr new_Jinkela_buffer_229 (
        .din(new_Jinkela_wire_298),
        .dout(new_Jinkela_wire_299)
    );

    spl2 new_Jinkela_splitter_261 (
        .a(_211_),
        .b(new_Jinkela_wire_1703),
        .c(new_Jinkela_wire_1704)
    );

    spl4L new_Jinkela_splitter_169 (
        .a(_244_),
        .d(new_Jinkela_wire_1390),
        .e(new_Jinkela_wire_1391),
        .b(new_Jinkela_wire_1392),
        .c(new_Jinkela_wire_1393)
    );

    bfr new_Jinkela_buffer_248 (
        .din(new_Jinkela_wire_325),
        .dout(new_Jinkela_wire_326)
    );

    spl2 new_Jinkela_splitter_262 (
        .a(_035_),
        .b(new_Jinkela_wire_1705),
        .c(new_Jinkela_wire_1706)
    );

    bfr new_Jinkela_buffer_947 (
        .din(new_Jinkela_wire_1357),
        .dout(new_Jinkela_wire_1358)
    );

    bfr new_Jinkela_buffer_230 (
        .din(new_Jinkela_wire_299),
        .dout(new_Jinkela_wire_300)
    );

    spl2 new_Jinkela_splitter_264 (
        .a(_007_),
        .b(new_Jinkela_wire_1709),
        .c(new_Jinkela_wire_1710)
    );

    spl2 new_Jinkela_splitter_167 (
        .a(_104_),
        .b(new_Jinkela_wire_1386),
        .c(new_Jinkela_wire_1387)
    );

    bfr new_Jinkela_buffer_271 (
        .din(new_Jinkela_wire_356),
        .dout(new_Jinkela_wire_357)
    );

    bfr new_Jinkela_buffer_952 (
        .din(new_Jinkela_wire_1380),
        .dout(new_Jinkela_wire_1381)
    );

    spl2 new_Jinkela_splitter_263 (
        .a(_176_),
        .b(new_Jinkela_wire_1707),
        .c(new_Jinkela_wire_1708)
    );

    bfr new_Jinkela_buffer_948 (
        .din(new_Jinkela_wire_1358),
        .dout(new_Jinkela_wire_1359)
    );

    bfr new_Jinkela_buffer_231 (
        .din(new_Jinkela_wire_300),
        .dout(new_Jinkela_wire_301)
    );

    bfr new_Jinkela_buffer_249 (
        .din(new_Jinkela_wire_326),
        .dout(new_Jinkela_wire_327)
    );

    bfr new_Jinkela_buffer_949 (
        .din(new_Jinkela_wire_1359),
        .dout(new_Jinkela_wire_1360)
    );

    bfr new_Jinkela_buffer_232 (
        .din(new_Jinkela_wire_301),
        .dout(new_Jinkela_wire_302)
    );

    bfr new_Jinkela_buffer_953 (
        .din(new_Jinkela_wire_1381),
        .dout(new_Jinkela_wire_1382)
    );

    spl4L new_Jinkela_splitter_158 (
        .a(new_Jinkela_wire_1360),
        .d(new_Jinkela_wire_1361),
        .e(new_Jinkela_wire_1362),
        .b(new_Jinkela_wire_1363),
        .c(new_Jinkela_wire_1364)
    );

    bfr new_Jinkela_buffer_233 (
        .din(new_Jinkela_wire_302),
        .dout(new_Jinkela_wire_303)
    );

    bfr new_Jinkela_buffer_960 (
        .din(_092_),
        .dout(new_Jinkela_wire_1407)
    );

    bfr new_Jinkela_buffer_250 (
        .din(new_Jinkela_wire_327),
        .dout(new_Jinkela_wire_328)
    );

    bfr new_Jinkela_buffer_954 (
        .din(new_Jinkela_wire_1382),
        .dout(new_Jinkela_wire_1383)
    );

    bfr new_Jinkela_buffer_234 (
        .din(new_Jinkela_wire_303),
        .dout(new_Jinkela_wire_304)
    );

    bfr new_Jinkela_buffer_956 (
        .din(_151_),
        .dout(new_Jinkela_wire_1395)
    );

    bfr new_Jinkela_buffer_272 (
        .din(new_Jinkela_wire_357),
        .dout(new_Jinkela_wire_358)
    );

    bfr new_Jinkela_buffer_955 (
        .din(_241_),
        .dout(new_Jinkela_wire_1394)
    );

    bfr new_Jinkela_buffer_235 (
        .din(new_Jinkela_wire_304),
        .dout(new_Jinkela_wire_305)
    );

    spl2 new_Jinkela_splitter_166 (
        .a(new_Jinkela_wire_1383),
        .b(new_Jinkela_wire_1384),
        .c(new_Jinkela_wire_1385)
    );

    bfr new_Jinkela_buffer_251 (
        .din(new_Jinkela_wire_328),
        .dout(new_Jinkela_wire_329)
    );

    spl2 new_Jinkela_splitter_171 (
        .a(_318_),
        .b(new_Jinkela_wire_1401),
        .c(new_Jinkela_wire_1402)
    );

    spl2 new_Jinkela_splitter_172 (
        .a(_309_),
        .b(new_Jinkela_wire_1403),
        .c(new_Jinkela_wire_1404)
    );

    bfr new_Jinkela_buffer_236 (
        .din(new_Jinkela_wire_305),
        .dout(new_Jinkela_wire_306)
    );

    bfr new_Jinkela_buffer_957 (
        .din(new_Jinkela_wire_1395),
        .dout(new_Jinkela_wire_1396)
    );

    bfr new_Jinkela_buffer_237 (
        .din(new_Jinkela_wire_306),
        .dout(new_Jinkela_wire_307)
    );

    bfr new_Jinkela_buffer_252 (
        .din(new_Jinkela_wire_329),
        .dout(new_Jinkela_wire_330)
    );

    bfr new_Jinkela_buffer_958 (
        .din(new_Jinkela_wire_1396),
        .dout(new_Jinkela_wire_1397)
    );

    bfr new_Jinkela_buffer_238 (
        .din(new_Jinkela_wire_307),
        .dout(new_Jinkela_wire_308)
    );

    spl2 new_Jinkela_splitter_173 (
        .a(_026_),
        .b(new_Jinkela_wire_1405),
        .c(new_Jinkela_wire_1406)
    );

    bfr new_Jinkela_buffer_273 (
        .din(new_Jinkela_wire_358),
        .dout(new_Jinkela_wire_359)
    );

    bfr new_Jinkela_buffer_959 (
        .din(new_Jinkela_wire_1397),
        .dout(new_Jinkela_wire_1398)
    );

    bfr new_Jinkela_buffer_239 (
        .din(new_Jinkela_wire_308),
        .dout(new_Jinkela_wire_309)
    );

    spl4L new_Jinkela_splitter_178 (
        .a(_226_),
        .d(new_Jinkela_wire_1423),
        .e(new_Jinkela_wire_1424),
        .b(new_Jinkela_wire_1425),
        .c(new_Jinkela_wire_1426)
    );

    spl2 new_Jinkela_splitter_174 (
        .a(new_Jinkela_wire_1407),
        .b(new_Jinkela_wire_1408),
        .c(new_Jinkela_wire_1409)
    );

    bfr new_Jinkela_buffer_115 (
        .din(new_Jinkela_wire_152),
        .dout(new_Jinkela_wire_153)
    );

    bfr new_Jinkela_buffer_253 (
        .din(new_Jinkela_wire_330),
        .dout(new_Jinkela_wire_331)
    );

    spl2 new_Jinkela_splitter_170 (
        .a(new_Jinkela_wire_1398),
        .b(new_Jinkela_wire_1399),
        .c(new_Jinkela_wire_1400)
    );

    spl2 new_Jinkela_splitter_26 (
        .a(new_Jinkela_wire_309),
        .b(new_Jinkela_wire_310),
        .c(new_Jinkela_wire_311)
    );

    spl2 new_Jinkela_splitter_176 (
        .a(_224_),
        .b(new_Jinkela_wire_1412),
        .c(new_Jinkela_wire_1413)
    );

    bfr new_Jinkela_buffer_254 (
        .din(new_Jinkela_wire_331),
        .dout(new_Jinkela_wire_332)
    );

    spl2 new_Jinkela_splitter_175 (
        .a(_333_),
        .b(new_Jinkela_wire_1410),
        .c(new_Jinkela_wire_1411)
    );

    bfr new_Jinkela_buffer_324 (
        .din(N135),
        .dout(new_Jinkela_wire_420)
    );

    spl2 new_Jinkela_splitter_177 (
        .a(_146_),
        .b(new_Jinkela_wire_1414),
        .c(new_Jinkela_wire_1415)
    );

    spl2 new_Jinkela_splitter_36 (
        .a(N61),
        .b(new_Jinkela_wire_422),
        .c(new_Jinkela_wire_424)
    );

    bfr new_Jinkela_buffer_274 (
        .din(new_Jinkela_wire_359),
        .dout(new_Jinkela_wire_360)
    );

    and_bi _685_ (
        .a(new_Jinkela_wire_1275),
        .b(new_Jinkela_wire_1307),
        .c(_282_)
    );

    and_bi _686_ (
        .a(new_Jinkela_wire_1311),
        .b(new_Jinkela_wire_696),
        .c(_283_)
    );

    and_bi _687_ (
        .a(new_Jinkela_wire_695),
        .b(new_Jinkela_wire_1310),
        .c(_284_)
    );

    or_bb _688_ (
        .a(_284_),
        .b(_283_),
        .c(new_net_697)
    );

    and_bi _689_ (
        .a(new_Jinkela_wire_1491),
        .b(new_Jinkela_wire_1161),
        .c(_285_)
    );

    and_bi _690_ (
        .a(new_Jinkela_wire_1469),
        .b(new_Jinkela_wire_1046),
        .c(_286_)
    );

    and_bi _691_ (
        .a(new_Jinkela_wire_1045),
        .b(new_Jinkela_wire_1468),
        .c(_287_)
    );

    or_bb _692_ (
        .a(_287_),
        .b(_286_),
        .c(N727)
    );

    or_bb _693_ (
        .a(new_Jinkela_wire_1571),
        .b(new_Jinkela_wire_1707),
        .c(_288_)
    );

    or_bb _694_ (
        .a(new_Jinkela_wire_1178),
        .b(new_Jinkela_wire_1552),
        .c(_289_)
    );

    or_bb _695_ (
        .a(new_Jinkela_wire_1302),
        .b(new_Jinkela_wire_1610),
        .c(_290_)
    );

    and_bi _696_ (
        .a(new_Jinkela_wire_137),
        .b(new_Jinkela_wire_1616),
        .c(_291_)
    );

    and_bi _697_ (
        .a(new_Jinkela_wire_1615),
        .b(new_Jinkela_wire_138),
        .c(_292_)
    );

    and_ii _698_ (
        .a(_292_),
        .b(_291_),
        .c(N738)
    );

    or_bi _699_ (
        .a(new_Jinkela_wire_1308),
        .b(new_Jinkela_wire_1464),
        .c(_293_)
    );

    and_bi _700_ (
        .a(new_Jinkela_wire_381),
        .b(new_Jinkela_wire_1317),
        .c(_294_)
    );

    and_bi _701_ (
        .a(new_Jinkela_wire_1316),
        .b(new_Jinkela_wire_382),
        .c(_295_)
    );

    and_ii _702_ (
        .a(_295_),
        .b(_294_),
        .c(new_net_699)
    );

    or_bi _703_ (
        .a(new_Jinkela_wire_1301),
        .b(new_Jinkela_wire_1493),
        .c(_296_)
    );

    and_bi _704_ (
        .a(new_Jinkela_wire_456),
        .b(new_Jinkela_wire_1473),
        .c(_297_)
    );

    and_bi _705_ (
        .a(new_Jinkela_wire_1472),
        .b(new_Jinkela_wire_455),
        .c(_298_)
    );

    and_ii _706_ (
        .a(_298_),
        .b(_297_),
        .c(N739)
    );

    and_bi _707_ (
        .a(new_Jinkela_wire_1272),
        .b(new_Jinkela_wire_1392),
        .c(_299_)
    );

    and_bi _708_ (
        .a(new_Jinkela_wire_1659),
        .b(new_Jinkela_wire_101),
        .c(_300_)
    );

    and_bi _709_ (
        .a(new_Jinkela_wire_100),
        .b(new_Jinkela_wire_1658),
        .c(_301_)
    );

    or_bb _710_ (
        .a(_301_),
        .b(_300_),
        .c(new_net_685)
    );

    or_bb _711_ (
        .a(new_Jinkela_wire_1391),
        .b(new_Jinkela_wire_1227),
        .c(_302_)
    );

    and_bi _712_ (
        .a(new_Jinkela_wire_1369),
        .b(new_Jinkela_wire_1129),
        .c(_303_)
    );

    and_bi _713_ (
        .a(new_Jinkela_wire_1128),
        .b(new_Jinkela_wire_1368),
        .c(_304_)
    );

    and_ii _714_ (
        .a(_304_),
        .b(_303_),
        .c(new_net_689)
    );

    or_bb _715_ (
        .a(new_Jinkela_wire_1390),
        .b(new_Jinkela_wire_1203),
        .c(_305_)
    );

    and_bi _716_ (
        .a(new_Jinkela_wire_1144),
        .b(new_Jinkela_wire_907),
        .c(_306_)
    );

    and_bi _717_ (
        .a(new_Jinkela_wire_906),
        .b(new_Jinkela_wire_1143),
        .c(_307_)
    );

    and_ii _718_ (
        .a(_307_),
        .b(_306_),
        .c(new_net_703)
    );

    or_bb _719_ (
        .a(new_Jinkela_wire_1177),
        .b(new_Jinkela_wire_1185),
        .c(_308_)
    );

    or_bi _720_ (
        .a(new_Jinkela_wire_1321),
        .b(new_Jinkela_wire_1363),
        .c(_309_)
    );

    and_bi _721_ (
        .a(new_Jinkela_wire_1404),
        .b(new_Jinkela_wire_1091),
        .c(_310_)
    );

    and_bi _722_ (
        .a(new_Jinkela_wire_1090),
        .b(new_Jinkela_wire_1403),
        .c(_311_)
    );

    and_ii _723_ (
        .a(_311_),
        .b(_310_),
        .c(N733)
    );

    or_bi _724_ (
        .a(new_Jinkela_wire_1423),
        .b(new_Jinkela_wire_1362),
        .c(_312_)
    );

    and_bi _725_ (
        .a(new_Jinkela_wire_1283),
        .b(new_Jinkela_wire_559),
        .c(_313_)
    );

    and_bi _726_ (
        .a(new_Jinkela_wire_558),
        .b(new_Jinkela_wire_1282),
        .c(_314_)
    );

    bfr new_Jinkela_buffer_80 (
        .din(new_Jinkela_wire_104),
        .dout(new_Jinkela_wire_105)
    );

    bfr new_Jinkela_buffer_652 (
        .din(new_Jinkela_wire_849),
        .dout(new_Jinkela_wire_850)
    );

    bfr new_Jinkela_buffer_961 (
        .din(new_Jinkela_wire_1415),
        .dout(new_Jinkela_wire_1416)
    );

    and_bi _517_ (
        .a(_127_),
        .b(_128_),
        .c(_129_)
    );

    bfr new_Jinkela_buffer_22 (
        .din(new_Jinkela_wire_27),
        .dout(new_Jinkela_wire_28)
    );

    bfr new_Jinkela_buffer_634 (
        .din(new_Jinkela_wire_823),
        .dout(new_Jinkela_wire_824)
    );

    or_bb _518_ (
        .a(new_Jinkela_wire_806),
        .b(new_Jinkela_wire_947),
        .c(_130_)
    );

    bfr new_Jinkela_buffer_968 (
        .din(_088_),
        .dout(new_Jinkela_wire_1427)
    );

    bfr new_Jinkela_buffer_36 (
        .din(new_Jinkela_wire_49),
        .dout(new_Jinkela_wire_50)
    );

    bfr new_Jinkela_buffer_701 (
        .din(new_Jinkela_wire_914),
        .dout(new_Jinkela_wire_915)
    );

    spl2 new_Jinkela_splitter_180 (
        .a(_189_),
        .b(new_Jinkela_wire_1432),
        .c(new_Jinkela_wire_1433)
    );

    and_bb _519_ (
        .a(new_Jinkela_wire_808),
        .b(new_Jinkela_wire_948),
        .c(_131_)
    );

    bfr new_Jinkela_buffer_970 (
        .din(new_net_685),
        .dout(new_Jinkela_wire_1431)
    );

    bfr new_Jinkela_buffer_23 (
        .din(new_Jinkela_wire_28),
        .dout(new_Jinkela_wire_29)
    );

    bfr new_Jinkela_buffer_635 (
        .din(new_Jinkela_wire_824),
        .dout(new_Jinkela_wire_825)
    );

    bfr new_Jinkela_buffer_962 (
        .din(new_Jinkela_wire_1416),
        .dout(new_Jinkela_wire_1417)
    );

    and_bi _520_ (
        .a(_130_),
        .b(_131_),
        .c(_132_)
    );

    bfr new_Jinkela_buffer_56 (
        .din(new_Jinkela_wire_77),
        .dout(new_Jinkela_wire_78)
    );

    bfr new_Jinkela_buffer_653 (
        .din(new_Jinkela_wire_850),
        .dout(new_Jinkela_wire_851)
    );

    or_bi _521_ (
        .a(new_Jinkela_wire_495),
        .b(new_Jinkela_wire_37),
        .c(_133_)
    );

    bfr new_Jinkela_buffer_24 (
        .din(new_Jinkela_wire_29),
        .dout(new_Jinkela_wire_30)
    );

    bfr new_Jinkela_buffer_636 (
        .din(new_Jinkela_wire_825),
        .dout(new_Jinkela_wire_826)
    );

    bfr new_Jinkela_buffer_963 (
        .din(new_Jinkela_wire_1417),
        .dout(new_Jinkela_wire_1418)
    );

    and_bi _522_ (
        .a(new_Jinkela_wire_494),
        .b(new_Jinkela_wire_35),
        .c(_134_)
    );

    bfr new_Jinkela_buffer_37 (
        .din(new_Jinkela_wire_50),
        .dout(new_Jinkela_wire_51)
    );

    bfr new_Jinkela_buffer_676 (
        .din(new_Jinkela_wire_881),
        .dout(new_Jinkela_wire_882)
    );

    or_bi _523_ (
        .a(_134_),
        .b(_133_),
        .c(_135_)
    );

    bfr new_Jinkela_buffer_969 (
        .din(new_Jinkela_wire_1427),
        .dout(new_Jinkela_wire_1428)
    );

    bfr new_Jinkela_buffer_25 (
        .din(new_Jinkela_wire_30),
        .dout(new_Jinkela_wire_31)
    );

    bfr new_Jinkela_buffer_637 (
        .din(new_Jinkela_wire_826),
        .dout(new_Jinkela_wire_827)
    );

    bfr new_Jinkela_buffer_964 (
        .din(new_Jinkela_wire_1418),
        .dout(new_Jinkela_wire_1419)
    );

    or_bi _524_ (
        .a(new_Jinkela_wire_1304),
        .b(new_Jinkela_wire_1446),
        .c(_136_)
    );

    spl2 new_Jinkela_splitter_15 (
        .a(N17),
        .b(new_Jinkela_wire_173),
        .c(new_Jinkela_wire_175)
    );

    bfr new_Jinkela_buffer_654 (
        .din(new_Jinkela_wire_851),
        .dout(new_Jinkela_wire_852)
    );

    spl2 new_Jinkela_splitter_181 (
        .a(_269_),
        .b(new_Jinkela_wire_1434),
        .c(new_Jinkela_wire_1435)
    );

    and_bi _525_ (
        .a(new_Jinkela_wire_1303),
        .b(new_Jinkela_wire_1445),
        .c(_137_)
    );

    spl2 new_Jinkela_splitter_184 (
        .a(_135_),
        .b(new_Jinkela_wire_1445),
        .c(new_Jinkela_wire_1446)
    );

    spl2 new_Jinkela_splitter_2 (
        .a(new_Jinkela_wire_31),
        .b(new_Jinkela_wire_32),
        .c(new_Jinkela_wire_33)
    );

    bfr new_Jinkela_buffer_638 (
        .din(new_Jinkela_wire_827),
        .dout(new_Jinkela_wire_828)
    );

    bfr new_Jinkela_buffer_965 (
        .din(new_Jinkela_wire_1419),
        .dout(new_Jinkela_wire_1420)
    );

    and_bi _526_ (
        .a(new_Jinkela_wire_1373),
        .b(new_Jinkela_wire_1153),
        .c(_138_)
    );

    bfr new_Jinkela_buffer_57 (
        .din(new_Jinkela_wire_78),
        .dout(new_Jinkela_wire_79)
    );

    spl2 new_Jinkela_splitter_84 (
        .a(N9),
        .b(new_Jinkela_wire_977),
        .c(new_Jinkela_wire_979)
    );

    spl2 new_Jinkela_splitter_179 (
        .a(new_Jinkela_wire_1428),
        .b(new_Jinkela_wire_1429),
        .c(new_Jinkela_wire_1430)
    );

    or_bb _527_ (
        .a(new_Jinkela_wire_1279),
        .b(new_Jinkela_wire_1149),
        .c(_139_)
    );

    bfr new_Jinkela_buffer_38 (
        .din(new_Jinkela_wire_51),
        .dout(new_Jinkela_wire_52)
    );

    bfr new_Jinkela_buffer_639 (
        .din(new_Jinkela_wire_828),
        .dout(new_Jinkela_wire_829)
    );

    bfr new_Jinkela_buffer_966 (
        .din(new_Jinkela_wire_1420),
        .dout(new_Jinkela_wire_1421)
    );

    or_bi _528_ (
        .a(new_Jinkela_wire_1152),
        .b(new_Jinkela_wire_1372),
        .c(_140_)
    );

    bfr new_Jinkela_buffer_39 (
        .din(new_Jinkela_wire_52),
        .dout(new_Jinkela_wire_53)
    );

    bfr new_Jinkela_buffer_655 (
        .din(new_Jinkela_wire_852),
        .dout(new_Jinkela_wire_853)
    );

    and_bi _529_ (
        .a(new_Jinkela_wire_1148),
        .b(new_Jinkela_wire_1511),
        .c(_141_)
    );

    bfr new_Jinkela_buffer_971 (
        .din(_091_),
        .dout(new_Jinkela_wire_1436)
    );

    bfr new_Jinkela_buffer_81 (
        .din(new_Jinkela_wire_110),
        .dout(new_Jinkela_wire_111)
    );

    bfr new_Jinkela_buffer_640 (
        .din(new_Jinkela_wire_829),
        .dout(new_Jinkela_wire_830)
    );

    bfr new_Jinkela_buffer_967 (
        .din(new_Jinkela_wire_1421),
        .dout(new_Jinkela_wire_1422)
    );

    and_bi _530_ (
        .a(_139_),
        .b(_141_),
        .c(_142_)
    );

    bfr new_Jinkela_buffer_40 (
        .din(new_Jinkela_wire_53),
        .dout(new_Jinkela_wire_54)
    );

    bfr new_Jinkela_buffer_677 (
        .din(new_Jinkela_wire_882),
        .dout(new_Jinkela_wire_883)
    );

    spl4L new_Jinkela_splitter_183 (
        .a(_253_),
        .d(new_Jinkela_wire_1441),
        .e(new_Jinkela_wire_1442),
        .b(new_Jinkela_wire_1443),
        .c(new_Jinkela_wire_1444)
    );

    and_bi _531_ (
        .a(new_Jinkela_wire_1375),
        .b(new_Jinkela_wire_1698),
        .c(_143_)
    );

    bfr new_Jinkela_buffer_58 (
        .din(new_Jinkela_wire_79),
        .dout(new_Jinkela_wire_80)
    );

    bfr new_Jinkela_buffer_641 (
        .din(new_Jinkela_wire_830),
        .dout(new_Jinkela_wire_831)
    );

    and_bi _532_ (
        .a(new_Jinkela_wire_1697),
        .b(new_Jinkela_wire_1374),
        .c(_144_)
    );

    bfr new_Jinkela_buffer_41 (
        .din(new_Jinkela_wire_54),
        .dout(new_Jinkela_wire_55)
    );

    bfr new_Jinkela_buffer_656 (
        .din(new_Jinkela_wire_853),
        .dout(new_Jinkela_wire_854)
    );

    bfr new_Jinkela_buffer_972 (
        .din(new_Jinkela_wire_1436),
        .dout(new_Jinkela_wire_1437)
    );

    or_bb _533_ (
        .a(_144_),
        .b(_143_),
        .c(_145_)
    );

    spl2 new_Jinkela_splitter_18 (
        .a(N49),
        .b(new_Jinkela_wire_208),
        .c(new_Jinkela_wire_210)
    );

    bfr new_Jinkela_buffer_642 (
        .din(new_Jinkela_wire_831),
        .dout(new_Jinkela_wire_832)
    );

    or_bi _534_ (
        .a(new_Jinkela_wire_1237),
        .b(new_Jinkela_wire_1346),
        .c(_146_)
    );

    bfr new_Jinkela_buffer_108 (
        .din(new_Jinkela_wire_145),
        .dout(new_Jinkela_wire_146)
    );

    spl2 new_Jinkela_splitter_185 (
        .a(new_Jinkela_wire_1447),
        .b(new_Jinkela_wire_1448),
        .c(new_Jinkela_wire_1449)
    );

    bfr new_Jinkela_buffer_42 (
        .din(new_Jinkela_wire_55),
        .dout(new_Jinkela_wire_56)
    );

    bfr new_Jinkela_buffer_973 (
        .din(new_Jinkela_wire_1437),
        .dout(new_Jinkela_wire_1438)
    );

    or_bb _535_ (
        .a(new_Jinkela_wire_1414),
        .b(new_Jinkela_wire_1430),
        .c(_147_)
    );

    bfr new_Jinkela_buffer_700 (
        .din(new_Jinkela_wire_908),
        .dout(new_Jinkela_wire_909)
    );

    bfr new_Jinkela_buffer_59 (
        .din(new_Jinkela_wire_80),
        .dout(new_Jinkela_wire_81)
    );

    bfr new_Jinkela_buffer_643 (
        .din(new_Jinkela_wire_832),
        .dout(new_Jinkela_wire_833)
    );

    or_bi _536_ (
        .a(new_Jinkela_wire_1348),
        .b(new_Jinkela_wire_1238),
        .c(_148_)
    );

    bfr new_Jinkela_buffer_974 (
        .din(_060_),
        .dout(new_Jinkela_wire_1447)
    );

    bfr new_Jinkela_buffer_43 (
        .din(new_Jinkela_wire_56),
        .dout(new_Jinkela_wire_57)
    );

    bfr new_Jinkela_buffer_657 (
        .din(new_Jinkela_wire_854),
        .dout(new_Jinkela_wire_855)
    );

    spl2 new_Jinkela_splitter_182 (
        .a(new_Jinkela_wire_1438),
        .b(new_Jinkela_wire_1439),
        .c(new_Jinkela_wire_1440)
    );

    or_bb _537_ (
        .a(new_Jinkela_wire_1572),
        .b(new_Jinkela_wire_1429),
        .c(_149_)
    );

    spl4L new_Jinkela_splitter_16 (
        .a(new_Jinkela_wire_175),
        .d(new_Jinkela_wire_176),
        .e(new_Jinkela_wire_177),
        .b(new_Jinkela_wire_178),
        .c(new_Jinkela_wire_179)
    );

    bfr new_Jinkela_buffer_644 (
        .din(new_Jinkela_wire_833),
        .dout(new_Jinkela_wire_834)
    );

    spl4L new_Jinkela_splitter_186 (
        .a(_085_),
        .d(new_Jinkela_wire_1450),
        .e(new_Jinkela_wire_1451),
        .b(new_Jinkela_wire_1452),
        .c(new_Jinkela_wire_1453)
    );

    and_bb _538_ (
        .a(new_Jinkela_wire_1207),
        .b(new_Jinkela_wire_1558),
        .c(_150_)
    );

    bfr new_Jinkela_buffer_44 (
        .din(new_Jinkela_wire_57),
        .dout(new_Jinkela_wire_58)
    );

    bfr new_Jinkela_buffer_678 (
        .din(new_Jinkela_wire_883),
        .dout(new_Jinkela_wire_884)
    );

    spl2 new_Jinkela_splitter_188 (
        .a(_285_),
        .b(new_Jinkela_wire_1468),
        .c(new_Jinkela_wire_1469)
    );

    or_ii _539_ (
        .a(new_Jinkela_wire_419),
        .b(new_Jinkela_wire_1050),
        .c(_151_)
    );

    bfr new_Jinkela_buffer_60 (
        .din(new_Jinkela_wire_81),
        .dout(new_Jinkela_wire_82)
    );

    bfr new_Jinkela_buffer_645 (
        .din(new_Jinkela_wire_834),
        .dout(new_Jinkela_wire_835)
    );

    bfr new_Jinkela_buffer_975 (
        .din(new_Jinkela_wire_1453),
        .dout(new_Jinkela_wire_1454)
    );

    or_bi _540_ (
        .a(new_Jinkela_wire_427),
        .b(new_Jinkela_wire_384),
        .c(_152_)
    );

    bfr new_Jinkela_buffer_45 (
        .din(new_Jinkela_wire_58),
        .dout(new_Jinkela_wire_59)
    );

    bfr new_Jinkela_buffer_658 (
        .din(new_Jinkela_wire_855),
        .dout(new_Jinkela_wire_856)
    );

    and_bi _541_ (
        .a(new_Jinkela_wire_425),
        .b(new_Jinkela_wire_388),
        .c(_153_)
    );

    bfr new_Jinkela_buffer_976 (
        .din(new_Jinkela_wire_1454),
        .dout(new_Jinkela_wire_1455)
    );

    bfr new_Jinkela_buffer_82 (
        .din(new_Jinkela_wire_111),
        .dout(new_Jinkela_wire_112)
    );

    bfr new_Jinkela_buffer_646 (
        .din(new_Jinkela_wire_835),
        .dout(new_Jinkela_wire_836)
    );

    spl2 new_Jinkela_splitter_190 (
        .a(_296_),
        .b(new_Jinkela_wire_1472),
        .c(new_Jinkela_wire_1473)
    );

    or_bi _542_ (
        .a(_153_),
        .b(_152_),
        .c(_154_)
    );

    bfr new_Jinkela_buffer_46 (
        .din(new_Jinkela_wire_59),
        .dout(new_Jinkela_wire_60)
    );

    or_bi _543_ (
        .a(new_Jinkela_wire_912),
        .b(new_Jinkela_wire_1016),
        .c(_155_)
    );

    bfr new_Jinkela_buffer_61 (
        .din(new_Jinkela_wire_82),
        .dout(new_Jinkela_wire_83)
    );

    spl2 new_Jinkela_splitter_71 (
        .a(new_Jinkela_wire_836),
        .b(new_Jinkela_wire_837),
        .c(new_Jinkela_wire_838)
    );

    spl3L new_Jinkela_splitter_191 (
        .a(_169_),
        .d(new_Jinkela_wire_1474),
        .b(new_Jinkela_wire_1475),
        .c(new_Jinkela_wire_1476)
    );

    and_bi _544_ (
        .a(new_Jinkela_wire_909),
        .b(new_Jinkela_wire_1017),
        .c(_156_)
    );

    bfr new_Jinkela_buffer_977 (
        .din(new_Jinkela_wire_1455),
        .dout(new_Jinkela_wire_1456)
    );

    bfr new_Jinkela_buffer_47 (
        .din(new_Jinkela_wire_60),
        .dout(new_Jinkela_wire_61)
    );

    bfr new_Jinkela_buffer_679 (
        .din(new_Jinkela_wire_884),
        .dout(new_Jinkela_wire_885)
    );

    or_bi _545_ (
        .a(_156_),
        .b(_155_),
        .c(_157_)
    );

    bfr new_Jinkela_buffer_994 (
        .din(new_net_689),
        .dout(new_Jinkela_wire_1498)
    );

    bfr new_Jinkela_buffer_659 (
        .din(new_Jinkela_wire_856),
        .dout(new_Jinkela_wire_857)
    );

    spl2 new_Jinkela_splitter_195 (
        .a(_098_),
        .b(new_Jinkela_wire_1494),
        .c(new_Jinkela_wire_1495)
    );

    or_bi _546_ (
        .a(new_Jinkela_wire_1691),
        .b(new_Jinkela_wire_1678),
        .c(_158_)
    );

    bfr new_Jinkela_buffer_107 (
        .din(new_Jinkela_wire_139),
        .dout(new_Jinkela_wire_140)
    );

    bfr new_Jinkela_buffer_978 (
        .din(new_Jinkela_wire_1456),
        .dout(new_Jinkela_wire_1457)
    );

    bfr new_Jinkela_buffer_48 (
        .din(new_Jinkela_wire_61),
        .dout(new_Jinkela_wire_62)
    );

    bfr new_Jinkela_buffer_660 (
        .din(new_Jinkela_wire_857),
        .dout(new_Jinkela_wire_858)
    );

    and_bi _547_ (
        .a(new_Jinkela_wire_1690),
        .b(new_Jinkela_wire_1677),
        .c(_159_)
    );

    bfr new_Jinkela_buffer_62 (
        .din(new_Jinkela_wire_83),
        .dout(new_Jinkela_wire_84)
    );

    or_bi _548_ (
        .a(_159_),
        .b(_158_),
        .c(_160_)
    );

    bfr new_Jinkela_buffer_727 (
        .din(new_Jinkela_wire_943),
        .dout(new_Jinkela_wire_944)
    );

    bfr new_Jinkela_buffer_979 (
        .din(new_Jinkela_wire_1457),
        .dout(new_Jinkela_wire_1458)
    );

    bfr new_Jinkela_buffer_49 (
        .din(new_Jinkela_wire_62),
        .dout(new_Jinkela_wire_63)
    );

    bfr new_Jinkela_buffer_661 (
        .din(new_Jinkela_wire_858),
        .dout(new_Jinkela_wire_859)
    );

    or_bi _549_ (
        .a(new_Jinkela_wire_1400),
        .b(new_Jinkela_wire_1620),
        .c(_161_)
    );

    bfr new_Jinkela_buffer_83 (
        .din(new_Jinkela_wire_112),
        .dout(new_Jinkela_wire_113)
    );

    bfr new_Jinkela_buffer_680 (
        .din(new_Jinkela_wire_885),
        .dout(new_Jinkela_wire_886)
    );

    spl2 new_Jinkela_splitter_189 (
        .a(_183_),
        .b(new_Jinkela_wire_1470),
        .c(new_Jinkela_wire_1471)
    );

    and_bi _550_ (
        .a(new_Jinkela_wire_1399),
        .b(new_Jinkela_wire_1619),
        .c(_162_)
    );

    bfr new_Jinkela_buffer_50 (
        .din(new_Jinkela_wire_63),
        .dout(new_Jinkela_wire_64)
    );

    bfr new_Jinkela_buffer_662 (
        .din(new_Jinkela_wire_859),
        .dout(new_Jinkela_wire_860)
    );

    bfr new_Jinkela_buffer_986 (
        .din(new_Jinkela_wire_1477),
        .dout(new_Jinkela_wire_1478)
    );

    and_bi _551_ (
        .a(_161_),
        .b(_162_),
        .c(_163_)
    );

    bfr new_Jinkela_buffer_980 (
        .din(new_Jinkela_wire_1458),
        .dout(new_Jinkela_wire_1459)
    );

    bfr new_Jinkela_buffer_63 (
        .din(new_Jinkela_wire_84),
        .dout(new_Jinkela_wire_85)
    );

    bfr new_Jinkela_buffer_702 (
        .din(new_Jinkela_wire_915),
        .dout(new_Jinkela_wire_916)
    );

    or_bb _552_ (
        .a(new_Jinkela_wire_1278),
        .b(new_Jinkela_wire_1336),
        .c(_164_)
    );

    bfr new_Jinkela_buffer_996 (
        .din(new_net_709),
        .dout(new_Jinkela_wire_1500)
    );

    bfr new_Jinkela_buffer_51 (
        .din(new_Jinkela_wire_64),
        .dout(new_Jinkela_wire_65)
    );

    bfr new_Jinkela_buffer_663 (
        .din(new_Jinkela_wire_860),
        .dout(new_Jinkela_wire_861)
    );

    bfr new_Jinkela_buffer_985 (
        .din(new_Jinkela_wire_1476),
        .dout(new_Jinkela_wire_1477)
    );

    and_bi _553_ (
        .a(new_Jinkela_wire_1337),
        .b(new_Jinkela_wire_1510),
        .c(_165_)
    );

    bfr new_Jinkela_buffer_981 (
        .din(new_Jinkela_wire_1459),
        .dout(new_Jinkela_wire_1460)
    );

    bfr new_Jinkela_buffer_681 (
        .din(new_Jinkela_wire_886),
        .dout(new_Jinkela_wire_887)
    );

    and_bi _554_ (
        .a(_164_),
        .b(_165_),
        .c(_166_)
    );

    spl2 new_Jinkela_splitter_5 (
        .a(new_Jinkela_wire_65),
        .b(new_Jinkela_wire_66),
        .c(new_Jinkela_wire_67)
    );

    bfr new_Jinkela_buffer_664 (
        .din(new_Jinkela_wire_861),
        .dout(new_Jinkela_wire_862)
    );

    and_bi _555_ (
        .a(new_Jinkela_wire_1142),
        .b(new_Jinkela_wire_1685),
        .c(_167_)
    );

    bfr new_Jinkela_buffer_982 (
        .din(new_Jinkela_wire_1460),
        .dout(new_Jinkela_wire_1461)
    );

    bfr new_Jinkela_buffer_84 (
        .din(new_Jinkela_wire_113),
        .dout(new_Jinkela_wire_114)
    );

    spl4L new_Jinkela_splitter_85 (
        .a(new_Jinkela_wire_979),
        .d(new_Jinkela_wire_980),
        .e(new_Jinkela_wire_981),
        .b(new_Jinkela_wire_982),
        .c(new_Jinkela_wire_983)
    );

    and_bi _556_ (
        .a(new_Jinkela_wire_1684),
        .b(new_Jinkela_wire_1141),
        .c(_168_)
    );

    spl2 new_Jinkela_splitter_87 (
        .a(N13),
        .b(new_Jinkela_wire_1012),
        .c(new_Jinkela_wire_1014)
    );

    spl2 new_Jinkela_splitter_196 (
        .a(_205_),
        .b(new_Jinkela_wire_1496),
        .c(new_Jinkela_wire_1497)
    );

    bfr new_Jinkela_buffer_64 (
        .din(new_Jinkela_wire_85),
        .dout(new_Jinkela_wire_86)
    );

    bfr new_Jinkela_buffer_665 (
        .din(new_Jinkela_wire_862),
        .dout(new_Jinkela_wire_863)
    );

    bfr new_Jinkela_buffer_995 (
        .din(new_net_705),
        .dout(new_Jinkela_wire_1499)
    );

    or_bb _557_ (
        .a(_168_),
        .b(_167_),
        .c(_169_)
    );

    bfr new_Jinkela_buffer_983 (
        .din(new_Jinkela_wire_1461),
        .dout(new_Jinkela_wire_1462)
    );

    bfr new_Jinkela_buffer_65 (
        .din(new_Jinkela_wire_86),
        .dout(new_Jinkela_wire_87)
    );

    bfr new_Jinkela_buffer_682 (
        .din(new_Jinkela_wire_887),
        .dout(new_Jinkela_wire_888)
    );

    or_bb _558_ (
        .a(new_Jinkela_wire_1481),
        .b(_150_),
        .c(_170_)
    );

    spl2 new_Jinkela_splitter_111 (
        .a(_279_),
        .b(new_Jinkela_wire_1165),
        .c(new_Jinkela_wire_1166)
    );

    spl2 new_Jinkela_splitter_119 (
        .a(_234_),
        .b(new_Jinkela_wire_1192),
        .c(new_Jinkela_wire_1193)
    );

    bfr new_Jinkela_buffer_855 (
        .din(new_Jinkela_wire_1118),
        .dout(new_Jinkela_wire_1119)
    );

    spl4L new_Jinkela_splitter_110 (
        .a(_217_),
        .d(new_Jinkela_wire_1161),
        .e(new_Jinkela_wire_1162),
        .b(new_Jinkela_wire_1163),
        .c(new_Jinkela_wire_1164)
    );

    bfr new_Jinkela_buffer_856 (
        .din(new_Jinkela_wire_1119),
        .dout(new_Jinkela_wire_1120)
    );

    spl2 new_Jinkela_splitter_113 (
        .a(_339_),
        .b(new_Jinkela_wire_1172),
        .c(new_Jinkela_wire_1173)
    );

    bfr new_Jinkela_buffer_857 (
        .din(new_Jinkela_wire_1120),
        .dout(new_Jinkela_wire_1121)
    );

    bfr new_Jinkela_buffer_858 (
        .din(new_Jinkela_wire_1121),
        .dout(new_Jinkela_wire_1122)
    );

    bfr new_Jinkela_buffer_872 (
        .din(_119_),
        .dout(new_Jinkela_wire_1167)
    );

    bfr new_Jinkela_buffer_859 (
        .din(new_Jinkela_wire_1122),
        .dout(new_Jinkela_wire_1123)
    );

    bfr new_Jinkela_buffer_873 (
        .din(new_Jinkela_wire_1167),
        .dout(new_Jinkela_wire_1168)
    );

    bfr new_Jinkela_buffer_860 (
        .din(new_Jinkela_wire_1123),
        .dout(new_Jinkela_wire_1124)
    );

    spl2 new_Jinkela_splitter_114 (
        .a(_029_),
        .b(new_Jinkela_wire_1174),
        .c(new_Jinkela_wire_1175)
    );

    bfr new_Jinkela_buffer_861 (
        .din(new_Jinkela_wire_1124),
        .dout(new_Jinkela_wire_1125)
    );

    bfr new_Jinkela_buffer_874 (
        .din(new_Jinkela_wire_1168),
        .dout(new_Jinkela_wire_1169)
    );

    bfr new_Jinkela_buffer_862 (
        .din(new_Jinkela_wire_1125),
        .dout(new_Jinkela_wire_1126)
    );

    bfr new_Jinkela_buffer_875 (
        .din(new_net_701),
        .dout(new_Jinkela_wire_1176)
    );

    bfr new_Jinkela_buffer_876 (
        .din(_087_),
        .dout(new_Jinkela_wire_1179)
    );

    bfr new_Jinkela_buffer_863 (
        .din(new_Jinkela_wire_1126),
        .dout(new_Jinkela_wire_1127)
    );

    spl2 new_Jinkela_splitter_112 (
        .a(new_Jinkela_wire_1169),
        .b(new_Jinkela_wire_1170),
        .c(new_Jinkela_wire_1171)
    );

    spl2 new_Jinkela_splitter_98 (
        .a(new_Jinkela_wire_1127),
        .b(new_Jinkela_wire_1128),
        .c(new_Jinkela_wire_1129)
    );

    spl2 new_Jinkela_splitter_115 (
        .a(_288_),
        .b(new_Jinkela_wire_1177),
        .c(new_Jinkela_wire_1178)
    );

    spl2 new_Jinkela_splitter_121 (
        .a(_149_),
        .b(new_Jinkela_wire_1207),
        .c(new_Jinkela_wire_1208)
    );

    spl3L new_Jinkela_splitter_117 (
        .a(_041_),
        .d(new_Jinkela_wire_1187),
        .b(new_Jinkela_wire_1188),
        .c(new_Jinkela_wire_1189)
    );

    bfr new_Jinkela_buffer_878 (
        .din(new_Jinkela_wire_1180),
        .dout(new_Jinkela_wire_1181)
    );

    bfr new_Jinkela_buffer_877 (
        .din(new_Jinkela_wire_1179),
        .dout(new_Jinkela_wire_1180)
    );

    spl2 new_Jinkela_splitter_118 (
        .a(new_Jinkela_wire_1189),
        .b(new_Jinkela_wire_1190),
        .c(new_Jinkela_wire_1191)
    );

    bfr new_Jinkela_buffer_879 (
        .din(new_Jinkela_wire_1181),
        .dout(new_Jinkela_wire_1182)
    );

    bfr new_Jinkela_buffer_882 (
        .din(new_Jinkela_wire_1193),
        .dout(new_Jinkela_wire_1194)
    );

    bfr new_Jinkela_buffer_880 (
        .din(new_Jinkela_wire_1182),
        .dout(new_Jinkela_wire_1183)
    );

    bfr new_Jinkela_buffer_896 (
        .din(_195_),
        .dout(new_Jinkela_wire_1214)
    );

    bfr new_Jinkela_buffer_881 (
        .din(new_Jinkela_wire_1183),
        .dout(new_Jinkela_wire_1184)
    );

    bfr new_Jinkela_buffer_885 (
        .din(new_Jinkela_wire_1196),
        .dout(new_Jinkela_wire_1197)
    );

    bfr new_Jinkela_buffer_883 (
        .din(new_Jinkela_wire_1194),
        .dout(new_Jinkela_wire_1195)
    );

    spl2 new_Jinkela_splitter_116 (
        .a(new_Jinkela_wire_1184),
        .b(new_Jinkela_wire_1185),
        .c(new_Jinkela_wire_1186)
    );

    spl2 new_Jinkela_splitter_124 (
        .a(_008_),
        .b(new_Jinkela_wire_1231),
        .c(new_Jinkela_wire_1232)
    );

    bfr new_Jinkela_buffer_884 (
        .din(new_Jinkela_wire_1195),
        .dout(new_Jinkela_wire_1196)
    );

    bfr new_Jinkela_buffer_892 (
        .din(new_Jinkela_wire_1209),
        .dout(new_Jinkela_wire_1210)
    );

    bfr new_Jinkela_buffer_891 (
        .din(new_Jinkela_wire_1208),
        .dout(new_Jinkela_wire_1209)
    );

    bfr new_Jinkela_buffer_886 (
        .din(new_Jinkela_wire_1197),
        .dout(new_Jinkela_wire_1198)
    );

    spl2 new_Jinkela_splitter_125 (
        .a(_230_),
        .b(new_Jinkela_wire_1233),
        .c(new_Jinkela_wire_1234)
    );

    bfr new_Jinkela_buffer_906 (
        .din(new_net_693),
        .dout(new_Jinkela_wire_1230)
    );

    spl2 new_Jinkela_splitter_122 (
        .a(new_Jinkela_wire_1214),
        .b(new_Jinkela_wire_1215),
        .c(new_Jinkela_wire_1216)
    );

    bfr new_Jinkela_buffer_464 (
        .din(new_Jinkela_wire_605),
        .dout(new_Jinkela_wire_606)
    );

    bfr new_Jinkela_buffer_445 (
        .din(new_Jinkela_wire_578),
        .dout(new_Jinkela_wire_579)
    );

    bfr new_Jinkela_buffer_512 (
        .din(new_Jinkela_wire_669),
        .dout(new_Jinkela_wire_670)
    );

    bfr new_Jinkela_buffer_446 (
        .din(new_Jinkela_wire_579),
        .dout(new_Jinkela_wire_580)
    );

    bfr new_Jinkela_buffer_465 (
        .din(new_Jinkela_wire_606),
        .dout(new_Jinkela_wire_607)
    );

    bfr new_Jinkela_buffer_447 (
        .din(new_Jinkela_wire_580),
        .dout(new_Jinkela_wire_581)
    );

    bfr new_Jinkela_buffer_487 (
        .din(new_Jinkela_wire_636),
        .dout(new_Jinkela_wire_637)
    );

    bfr new_Jinkela_buffer_448 (
        .din(new_Jinkela_wire_581),
        .dout(new_Jinkela_wire_582)
    );

    bfr new_Jinkela_buffer_466 (
        .din(new_Jinkela_wire_607),
        .dout(new_Jinkela_wire_608)
    );

    bfr new_Jinkela_buffer_449 (
        .din(new_Jinkela_wire_582),
        .dout(new_Jinkela_wire_583)
    );

    spl2 new_Jinkela_splitter_63 (
        .a(N5),
        .b(new_Jinkela_wire_732),
        .c(new_Jinkela_wire_734)
    );

    bfr new_Jinkela_buffer_450 (
        .din(new_Jinkela_wire_583),
        .dout(new_Jinkela_wire_584)
    );

    bfr new_Jinkela_buffer_467 (
        .din(new_Jinkela_wire_608),
        .dout(new_Jinkela_wire_609)
    );

    bfr new_Jinkela_buffer_451 (
        .din(new_Jinkela_wire_584),
        .dout(new_Jinkela_wire_585)
    );

    bfr new_Jinkela_buffer_488 (
        .din(new_Jinkela_wire_637),
        .dout(new_Jinkela_wire_638)
    );

    bfr new_Jinkela_buffer_452 (
        .din(new_Jinkela_wire_585),
        .dout(new_Jinkela_wire_586)
    );

    bfr new_Jinkela_buffer_468 (
        .din(new_Jinkela_wire_609),
        .dout(new_Jinkela_wire_610)
    );

    bfr new_Jinkela_buffer_453 (
        .din(new_Jinkela_wire_586),
        .dout(new_Jinkela_wire_587)
    );

    bfr new_Jinkela_buffer_511 (
        .din(new_Jinkela_wire_663),
        .dout(new_Jinkela_wire_664)
    );

    bfr new_Jinkela_buffer_454 (
        .din(new_Jinkela_wire_587),
        .dout(new_Jinkela_wire_588)
    );

    bfr new_Jinkela_buffer_469 (
        .din(new_Jinkela_wire_610),
        .dout(new_Jinkela_wire_611)
    );

    bfr new_Jinkela_buffer_455 (
        .din(new_Jinkela_wire_588),
        .dout(new_Jinkela_wire_589)
    );

    bfr new_Jinkela_buffer_489 (
        .din(new_Jinkela_wire_638),
        .dout(new_Jinkela_wire_639)
    );

    bfr new_Jinkela_buffer_456 (
        .din(new_Jinkela_wire_589),
        .dout(new_Jinkela_wire_590)
    );

    bfr new_Jinkela_buffer_470 (
        .din(new_Jinkela_wire_611),
        .dout(new_Jinkela_wire_612)
    );

    bfr new_Jinkela_buffer_457 (
        .din(new_Jinkela_wire_590),
        .dout(new_Jinkela_wire_591)
    );

    bfr new_Jinkela_buffer_458 (
        .din(new_Jinkela_wire_591),
        .dout(new_Jinkela_wire_592)
    );

    bfr new_Jinkela_buffer_471 (
        .din(new_Jinkela_wire_612),
        .dout(new_Jinkela_wire_613)
    );

    spl2 new_Jinkela_splitter_50 (
        .a(new_Jinkela_wire_592),
        .b(new_Jinkela_wire_593),
        .c(new_Jinkela_wire_594)
    );

    bfr new_Jinkela_buffer_472 (
        .din(new_Jinkela_wire_613),
        .dout(new_Jinkela_wire_614)
    );

    bfr new_Jinkela_buffer_490 (
        .din(new_Jinkela_wire_639),
        .dout(new_Jinkela_wire_640)
    );

    bfr new_Jinkela_buffer_537 (
        .din(new_Jinkela_wire_697),
        .dout(new_Jinkela_wire_698)
    );

    bfr new_Jinkela_buffer_473 (
        .din(new_Jinkela_wire_614),
        .dout(new_Jinkela_wire_615)
    );

    bfr new_Jinkela_buffer_491 (
        .din(new_Jinkela_wire_640),
        .dout(new_Jinkela_wire_641)
    );

    bfr new_Jinkela_buffer_474 (
        .din(new_Jinkela_wire_615),
        .dout(new_Jinkela_wire_616)
    );

    bfr new_Jinkela_buffer_513 (
        .din(new_Jinkela_wire_670),
        .dout(new_Jinkela_wire_671)
    );

    bfr new_Jinkela_buffer_475 (
        .din(new_Jinkela_wire_616),
        .dout(new_Jinkela_wire_617)
    );

    bfr new_Jinkela_buffer_492 (
        .din(new_Jinkela_wire_641),
        .dout(new_Jinkela_wire_642)
    );

    bfr new_Jinkela_buffer_476 (
        .din(new_Jinkela_wire_617),
        .dout(new_Jinkela_wire_618)
    );

    spl4L new_Jinkela_splitter_64 (
        .a(new_Jinkela_wire_734),
        .d(new_Jinkela_wire_735),
        .e(new_Jinkela_wire_736),
        .b(new_Jinkela_wire_737),
        .c(new_Jinkela_wire_738)
    );

    bfr new_Jinkela_buffer_591 (
        .din(N130),
        .dout(new_Jinkela_wire_767)
    );

    bfr new_Jinkela_buffer_477 (
        .din(new_Jinkela_wire_618),
        .dout(new_Jinkela_wire_619)
    );

    bfr new_Jinkela_buffer_666 (
        .din(new_Jinkela_wire_863),
        .dout(new_Jinkela_wire_864)
    );

    bfr new_Jinkela_buffer_703 (
        .din(new_Jinkela_wire_916),
        .dout(new_Jinkela_wire_917)
    );

    bfr new_Jinkela_buffer_667 (
        .din(new_Jinkela_wire_864),
        .dout(new_Jinkela_wire_865)
    );

    bfr new_Jinkela_buffer_683 (
        .din(new_Jinkela_wire_888),
        .dout(new_Jinkela_wire_889)
    );

    bfr new_Jinkela_buffer_668 (
        .din(new_Jinkela_wire_865),
        .dout(new_Jinkela_wire_866)
    );

    bfr new_Jinkela_buffer_669 (
        .din(new_Jinkela_wire_866),
        .dout(new_Jinkela_wire_867)
    );

    bfr new_Jinkela_buffer_684 (
        .din(new_Jinkela_wire_889),
        .dout(new_Jinkela_wire_890)
    );

    bfr new_Jinkela_buffer_670 (
        .din(new_Jinkela_wire_867),
        .dout(new_Jinkela_wire_868)
    );

    bfr new_Jinkela_buffer_704 (
        .din(new_Jinkela_wire_917),
        .dout(new_Jinkela_wire_918)
    );

    bfr new_Jinkela_buffer_671 (
        .din(new_Jinkela_wire_868),
        .dout(new_Jinkela_wire_869)
    );

    bfr new_Jinkela_buffer_685 (
        .din(new_Jinkela_wire_890),
        .dout(new_Jinkela_wire_891)
    );

    bfr new_Jinkela_buffer_672 (
        .din(new_Jinkela_wire_869),
        .dout(new_Jinkela_wire_870)
    );

    bfr new_Jinkela_buffer_728 (
        .din(new_Jinkela_wire_949),
        .dout(new_Jinkela_wire_950)
    );

    bfr new_Jinkela_buffer_753 (
        .din(new_Jinkela_wire_977),
        .dout(new_Jinkela_wire_978)
    );

    bfr new_Jinkela_buffer_673 (
        .din(new_Jinkela_wire_870),
        .dout(new_Jinkela_wire_871)
    );

    bfr new_Jinkela_buffer_686 (
        .din(new_Jinkela_wire_891),
        .dout(new_Jinkela_wire_892)
    );

    spl2 new_Jinkela_splitter_74 (
        .a(new_Jinkela_wire_871),
        .b(new_Jinkela_wire_872),
        .c(new_Jinkela_wire_873)
    );

    bfr new_Jinkela_buffer_687 (
        .din(new_Jinkela_wire_892),
        .dout(new_Jinkela_wire_893)
    );

    bfr new_Jinkela_buffer_705 (
        .din(new_Jinkela_wire_918),
        .dout(new_Jinkela_wire_919)
    );

    spl4L new_Jinkela_splitter_88 (
        .a(new_Jinkela_wire_1014),
        .d(new_Jinkela_wire_1015),
        .e(new_Jinkela_wire_1016),
        .b(new_Jinkela_wire_1017),
        .c(new_Jinkela_wire_1018)
    );

    bfr new_Jinkela_buffer_688 (
        .din(new_Jinkela_wire_893),
        .dout(new_Jinkela_wire_894)
    );

    bfr new_Jinkela_buffer_706 (
        .din(new_Jinkela_wire_919),
        .dout(new_Jinkela_wire_920)
    );

    bfr new_Jinkela_buffer_689 (
        .din(new_Jinkela_wire_894),
        .dout(new_Jinkela_wire_895)
    );

    bfr new_Jinkela_buffer_729 (
        .din(new_Jinkela_wire_950),
        .dout(new_Jinkela_wire_951)
    );

    bfr new_Jinkela_buffer_690 (
        .din(new_Jinkela_wire_895),
        .dout(new_Jinkela_wire_896)
    );

    bfr new_Jinkela_buffer_707 (
        .din(new_Jinkela_wire_920),
        .dout(new_Jinkela_wire_921)
    );

    bfr new_Jinkela_buffer_691 (
        .din(new_Jinkela_wire_896),
        .dout(new_Jinkela_wire_897)
    );

    spl2 new_Jinkela_splitter_90 (
        .a(N137),
        .b(new_Jinkela_wire_1047),
        .c(new_Jinkela_wire_1052)
    );

    bfr new_Jinkela_buffer_692 (
        .din(new_Jinkela_wire_897),
        .dout(new_Jinkela_wire_898)
    );

    bfr new_Jinkela_buffer_708 (
        .din(new_Jinkela_wire_921),
        .dout(new_Jinkela_wire_922)
    );

    bfr new_Jinkela_buffer_693 (
        .din(new_Jinkela_wire_898),
        .dout(new_Jinkela_wire_899)
    );

    bfr new_Jinkela_buffer_730 (
        .din(new_Jinkela_wire_951),
        .dout(new_Jinkela_wire_952)
    );

    bfr new_Jinkela_buffer_694 (
        .din(new_Jinkela_wire_899),
        .dout(new_Jinkela_wire_900)
    );

    bfr new_Jinkela_buffer_709 (
        .din(new_Jinkela_wire_922),
        .dout(new_Jinkela_wire_923)
    );

    bfr new_Jinkela_buffer_695 (
        .din(new_Jinkela_wire_900),
        .dout(new_Jinkela_wire_901)
    );

    bfr new_Jinkela_buffer_754 (
        .din(new_Jinkela_wire_983),
        .dout(new_Jinkela_wire_984)
    );

    bfr new_Jinkela_buffer_696 (
        .din(new_Jinkela_wire_901),
        .dout(new_Jinkela_wire_902)
    );

    bfr new_Jinkela_buffer_710 (
        .din(new_Jinkela_wire_923),
        .dout(new_Jinkela_wire_924)
    );

    bfr new_Jinkela_buffer_697 (
        .din(new_Jinkela_wire_902),
        .dout(new_Jinkela_wire_903)
    );

    bfr new_Jinkela_buffer_731 (
        .din(new_Jinkela_wire_952),
        .dout(new_Jinkela_wire_953)
    );

    bfr new_Jinkela_buffer_698 (
        .din(new_Jinkela_wire_903),
        .dout(new_Jinkela_wire_904)
    );

    bfr new_Jinkela_buffer_711 (
        .din(new_Jinkela_wire_924),
        .dout(new_Jinkela_wire_925)
    );

    bfr new_Jinkela_buffer_255 (
        .din(new_Jinkela_wire_332),
        .dout(new_Jinkela_wire_333)
    );

    spl2 new_Jinkela_splitter_39 (
        .a(N85),
        .b(new_Jinkela_wire_457),
        .c(new_Jinkela_wire_459)
    );

    bfr new_Jinkela_buffer_325 (
        .din(new_Jinkela_wire_420),
        .dout(new_Jinkela_wire_421)
    );

    bfr new_Jinkela_buffer_256 (
        .din(new_Jinkela_wire_333),
        .dout(new_Jinkela_wire_334)
    );

    bfr new_Jinkela_buffer_275 (
        .din(new_Jinkela_wire_360),
        .dout(new_Jinkela_wire_361)
    );

    bfr new_Jinkela_buffer_257 (
        .din(new_Jinkela_wire_334),
        .dout(new_Jinkela_wire_335)
    );

    bfr new_Jinkela_buffer_297 (
        .din(new_Jinkela_wire_390),
        .dout(new_Jinkela_wire_391)
    );

    bfr new_Jinkela_buffer_258 (
        .din(new_Jinkela_wire_335),
        .dout(new_Jinkela_wire_336)
    );

    bfr new_Jinkela_buffer_276 (
        .din(new_Jinkela_wire_361),
        .dout(new_Jinkela_wire_362)
    );

    bfr new_Jinkela_buffer_259 (
        .din(new_Jinkela_wire_336),
        .dout(new_Jinkela_wire_337)
    );

    bfr new_Jinkela_buffer_326 (
        .din(new_Jinkela_wire_422),
        .dout(new_Jinkela_wire_423)
    );

    bfr new_Jinkela_buffer_260 (
        .din(new_Jinkela_wire_337),
        .dout(new_Jinkela_wire_338)
    );

    bfr new_Jinkela_buffer_277 (
        .din(new_Jinkela_wire_362),
        .dout(new_Jinkela_wire_363)
    );

    bfr new_Jinkela_buffer_261 (
        .din(new_Jinkela_wire_338),
        .dout(new_Jinkela_wire_339)
    );

    bfr new_Jinkela_buffer_298 (
        .din(new_Jinkela_wire_391),
        .dout(new_Jinkela_wire_392)
    );

    bfr new_Jinkela_buffer_262 (
        .din(new_Jinkela_wire_339),
        .dout(new_Jinkela_wire_340)
    );

    bfr new_Jinkela_buffer_278 (
        .din(new_Jinkela_wire_363),
        .dout(new_Jinkela_wire_364)
    );

    bfr new_Jinkela_buffer_263 (
        .din(new_Jinkela_wire_340),
        .dout(new_Jinkela_wire_341)
    );

    spl2 new_Jinkela_splitter_42 (
        .a(N117),
        .b(new_Jinkela_wire_491),
        .c(new_Jinkela_wire_493)
    );

    bfr new_Jinkela_buffer_264 (
        .din(new_Jinkela_wire_341),
        .dout(new_Jinkela_wire_342)
    );

    bfr new_Jinkela_buffer_279 (
        .din(new_Jinkela_wire_364),
        .dout(new_Jinkela_wire_365)
    );

    bfr new_Jinkela_buffer_265 (
        .din(new_Jinkela_wire_342),
        .dout(new_Jinkela_wire_343)
    );

    bfr new_Jinkela_buffer_299 (
        .din(new_Jinkela_wire_392),
        .dout(new_Jinkela_wire_393)
    );

    bfr new_Jinkela_buffer_266 (
        .din(new_Jinkela_wire_343),
        .dout(new_Jinkela_wire_344)
    );

    bfr new_Jinkela_buffer_280 (
        .din(new_Jinkela_wire_365),
        .dout(new_Jinkela_wire_366)
    );

    bfr new_Jinkela_buffer_267 (
        .din(new_Jinkela_wire_344),
        .dout(new_Jinkela_wire_345)
    );

    spl4L new_Jinkela_splitter_37 (
        .a(new_Jinkela_wire_424),
        .d(new_Jinkela_wire_425),
        .e(new_Jinkela_wire_426),
        .b(new_Jinkela_wire_427),
        .c(new_Jinkela_wire_428)
    );

    bfr new_Jinkela_buffer_268 (
        .din(new_Jinkela_wire_345),
        .dout(new_Jinkela_wire_346)
    );

    bfr new_Jinkela_buffer_281 (
        .din(new_Jinkela_wire_366),
        .dout(new_Jinkela_wire_367)
    );

    spl2 new_Jinkela_splitter_29 (
        .a(new_Jinkela_wire_346),
        .b(new_Jinkela_wire_347),
        .c(new_Jinkela_wire_348)
    );

    bfr new_Jinkela_buffer_282 (
        .din(new_Jinkela_wire_367),
        .dout(new_Jinkela_wire_368)
    );

    bfr new_Jinkela_buffer_300 (
        .din(new_Jinkela_wire_393),
        .dout(new_Jinkela_wire_394)
    );

    spl4L new_Jinkela_splitter_40 (
        .a(new_Jinkela_wire_459),
        .d(new_Jinkela_wire_460),
        .e(new_Jinkela_wire_461),
        .b(new_Jinkela_wire_462),
        .c(new_Jinkela_wire_463)
    );

    bfr new_Jinkela_buffer_283 (
        .din(new_Jinkela_wire_368),
        .dout(new_Jinkela_wire_369)
    );

    bfr new_Jinkela_buffer_301 (
        .din(new_Jinkela_wire_394),
        .dout(new_Jinkela_wire_395)
    );

    bfr new_Jinkela_buffer_284 (
        .din(new_Jinkela_wire_369),
        .dout(new_Jinkela_wire_370)
    );

    bfr new_Jinkela_buffer_285 (
        .din(new_Jinkela_wire_370),
        .dout(new_Jinkela_wire_371)
    );

    bfr new_Jinkela_buffer_302 (
        .din(new_Jinkela_wire_395),
        .dout(new_Jinkela_wire_396)
    );

    bfr new_Jinkela_buffer_286 (
        .din(new_Jinkela_wire_371),
        .dout(new_Jinkela_wire_372)
    );

    bfr new_Jinkela_buffer_327 (
        .din(new_Jinkela_wire_428),
        .dout(new_Jinkela_wire_429)
    );

    bfr new_Jinkela_buffer_287 (
        .din(new_Jinkela_wire_372),
        .dout(new_Jinkela_wire_373)
    );

    bfr new_Jinkela_buffer_303 (
        .din(new_Jinkela_wire_396),
        .dout(new_Jinkela_wire_397)
    );

    and_ii _727_ (
        .a(_314_),
        .b(_313_),
        .c(N729)
    );

    bfr new_Jinkela_buffer_984 (
        .din(new_Jinkela_wire_1462),
        .dout(new_Jinkela_wire_1463)
    );

    or_bb _728_ (
        .a(new_Jinkela_wire_1320),
        .b(new_Jinkela_wire_1607),
        .c(_315_)
    );

    spl2 new_Jinkela_splitter_200 (
        .a(_194_),
        .b(new_Jinkela_wire_1512),
        .c(new_Jinkela_wire_1513)
    );

    bfr new_Jinkela_buffer_987 (
        .din(new_Jinkela_wire_1478),
        .dout(new_Jinkela_wire_1479)
    );

    and_bi _729_ (
        .a(new_Jinkela_wire_731),
        .b(new_Jinkela_wire_1670),
        .c(_316_)
    );

    spl4L new_Jinkela_splitter_187 (
        .a(new_Jinkela_wire_1463),
        .d(new_Jinkela_wire_1464),
        .e(new_Jinkela_wire_1465),
        .b(new_Jinkela_wire_1466),
        .c(new_Jinkela_wire_1467)
    );

    and_bi _730_ (
        .a(new_Jinkela_wire_1669),
        .b(new_Jinkela_wire_730),
        .c(_317_)
    );

    and_ii _731_ (
        .a(_317_),
        .b(_316_),
        .c(N734)
    );

    bfr new_Jinkela_buffer_988 (
        .din(new_Jinkela_wire_1479),
        .dout(new_Jinkela_wire_1480)
    );

    or_bb _732_ (
        .a(new_Jinkela_wire_1425),
        .b(new_Jinkela_wire_1609),
        .c(_318_)
    );

    and_bi _733_ (
        .a(new_Jinkela_wire_348),
        .b(new_Jinkela_wire_1402),
        .c(_319_)
    );

    bfr new_Jinkela_buffer_989 (
        .din(new_Jinkela_wire_1482),
        .dout(new_Jinkela_wire_1483)
    );

    spl2 new_Jinkela_splitter_198 (
        .a(_171_),
        .b(new_Jinkela_wire_1503),
        .c(new_Jinkela_wire_1504)
    );

    and_bi _734_ (
        .a(new_Jinkela_wire_1401),
        .b(new_Jinkela_wire_347),
        .c(_320_)
    );

    spl2 new_Jinkela_splitter_192 (
        .a(new_Jinkela_wire_1480),
        .b(new_Jinkela_wire_1481),
        .c(new_Jinkela_wire_1482)
    );

    spl2 new_Jinkela_splitter_197 (
        .a(_066_),
        .b(new_Jinkela_wire_1501),
        .c(new_Jinkela_wire_1502)
    );

    and_ii _735_ (
        .a(_320_),
        .b(_319_),
        .c(N730)
    );

    or_bi _736_ (
        .a(new_Jinkela_wire_1319),
        .b(new_Jinkela_wire_1490),
        .c(_321_)
    );

    spl2 new_Jinkela_splitter_199 (
        .a(_140_),
        .b(new_Jinkela_wire_1510),
        .c(new_Jinkela_wire_1511)
    );

    bfr new_Jinkela_buffer_997 (
        .din(new_Jinkela_wire_1504),
        .dout(new_Jinkela_wire_1505)
    );

    and_bi _737_ (
        .a(new_Jinkela_wire_1635),
        .b(new_Jinkela_wire_417),
        .c(_322_)
    );

    spl2 new_Jinkela_splitter_193 (
        .a(new_Jinkela_wire_1483),
        .b(new_Jinkela_wire_1484),
        .c(new_Jinkela_wire_1485)
    );

    and_bi _738_ (
        .a(new_Jinkela_wire_416),
        .b(new_Jinkela_wire_1634),
        .c(_323_)
    );

    bfr new_Jinkela_buffer_990 (
        .din(new_Jinkela_wire_1485),
        .dout(new_Jinkela_wire_1486)
    );

    and_ii _739_ (
        .a(_323_),
        .b(_322_),
        .c(N735)
    );

    spl2 new_Jinkela_splitter_203 (
        .a(_017_),
        .b(new_Jinkela_wire_1521),
        .c(new_Jinkela_wire_1522)
    );

    or_bi _740_ (
        .a(new_Jinkela_wire_1299),
        .b(new_Jinkela_wire_1253),
        .c(_324_)
    );

    bfr new_Jinkela_buffer_998 (
        .din(new_Jinkela_wire_1505),
        .dout(new_Jinkela_wire_1506)
    );

    and_bi _741_ (
        .a(new_Jinkela_wire_1666),
        .b(new_Jinkela_wire_242),
        .c(_325_)
    );

    bfr new_Jinkela_buffer_991 (
        .din(new_Jinkela_wire_1486),
        .dout(new_Jinkela_wire_1487)
    );

    and_bi _742_ (
        .a(new_Jinkela_wire_241),
        .b(new_Jinkela_wire_1665),
        .c(_326_)
    );

    and_ii _743_ (
        .a(_326_),
        .b(_325_),
        .c(N736)
    );

    bfr new_Jinkela_buffer_992 (
        .din(new_Jinkela_wire_1487),
        .dout(new_Jinkela_wire_1488)
    );

    or_bi _744_ (
        .a(new_Jinkela_wire_1300),
        .b(new_Jinkela_wire_1361),
        .c(_327_)
    );

    bfr new_Jinkela_buffer_1002 (
        .din(_179_),
        .dout(new_Jinkela_wire_1514)
    );

    bfr new_Jinkela_buffer_999 (
        .din(new_Jinkela_wire_1506),
        .dout(new_Jinkela_wire_1507)
    );

    and_bi _745_ (
        .a(new_Jinkela_wire_1524),
        .b(new_Jinkela_wire_873),
        .c(_328_)
    );

    bfr new_Jinkela_buffer_993 (
        .din(new_Jinkela_wire_1488),
        .dout(new_Jinkela_wire_1489)
    );

    and_bi _746_ (
        .a(new_Jinkela_wire_872),
        .b(new_Jinkela_wire_1523),
        .c(_329_)
    );

    and_ii _747_ (
        .a(_329_),
        .b(_328_),
        .c(N737)
    );

    spl4L new_Jinkela_splitter_194 (
        .a(new_Jinkela_wire_1489),
        .d(new_Jinkela_wire_1490),
        .e(new_Jinkela_wire_1491),
        .b(new_Jinkela_wire_1492),
        .c(new_Jinkela_wire_1493)
    );

    and_bi _748_ (
        .a(new_Jinkela_wire_1492),
        .b(new_Jinkela_wire_1424),
        .c(_330_)
    );

    bfr new_Jinkela_buffer_1003 (
        .din(new_Jinkela_wire_1514),
        .dout(new_Jinkela_wire_1515)
    );

    and_bi _749_ (
        .a(new_Jinkela_wire_1700),
        .b(new_Jinkela_wire_942),
        .c(_331_)
    );

    spl2 new_Jinkela_splitter_202 (
        .a(_276_),
        .b(new_Jinkela_wire_1519),
        .c(new_Jinkela_wire_1520)
    );

    bfr new_Jinkela_buffer_1000 (
        .din(new_Jinkela_wire_1507),
        .dout(new_Jinkela_wire_1508)
    );

    and_bi _750_ (
        .a(new_Jinkela_wire_941),
        .b(new_Jinkela_wire_1699),
        .c(_332_)
    );

    bfr new_Jinkela_buffer_1001 (
        .din(new_Jinkela_wire_1508),
        .dout(new_Jinkela_wire_1509)
    );

    or_bb _751_ (
        .a(_332_),
        .b(_331_),
        .c(N731)
    );

    or_bi _752_ (
        .a(new_Jinkela_wire_1318),
        .b(new_Jinkela_wire_1252),
        .c(_333_)
    );

    bfr new_Jinkela_buffer_1004 (
        .din(new_Jinkela_wire_1515),
        .dout(new_Jinkela_wire_1516)
    );

    and_bi _753_ (
        .a(new_Jinkela_wire_1411),
        .b(new_Jinkela_wire_594),
        .c(_334_)
    );

    and_bi _754_ (
        .a(new_Jinkela_wire_593),
        .b(new_Jinkela_wire_1410),
        .c(_335_)
    );

    spl2 new_Jinkela_splitter_204 (
        .a(_327_),
        .b(new_Jinkela_wire_1523),
        .c(new_Jinkela_wire_1524)
    );

    spl2 new_Jinkela_splitter_201 (
        .a(new_Jinkela_wire_1516),
        .b(new_Jinkela_wire_1517),
        .c(new_Jinkela_wire_1518)
    );

    and_ii _755_ (
        .a(_335_),
        .b(_334_),
        .c(N732)
    );

    spl2 new_Jinkela_splitter_206 (
        .a(_216_),
        .b(new_Jinkela_wire_1530),
        .c(new_Jinkela_wire_1531)
    );

    spl2 new_Jinkela_splitter_205 (
        .a(_348_),
        .b(new_Jinkela_wire_1528),
        .c(new_Jinkela_wire_1529)
    );

    bfr new_Jinkela_buffer_1006 (
        .din(new_Jinkela_wire_1525),
        .dout(new_Jinkela_wire_1526)
    );

    bfr new_Jinkela_buffer_1005 (
        .din(_237_),
        .dout(new_Jinkela_wire_1525)
    );

    spl2 new_Jinkela_splitter_208 (
        .a(_014_),
        .b(new_Jinkela_wire_1534),
        .c(new_Jinkela_wire_1535)
    );

    bfr new_Jinkela_buffer_1007 (
        .din(new_Jinkela_wire_1526),
        .dout(new_Jinkela_wire_1527)
    );

    spl2 new_Jinkela_splitter_207 (
        .a(_057_),
        .b(new_Jinkela_wire_1532),
        .c(new_Jinkela_wire_1533)
    );

    bfr new_Jinkela_buffer_1008 (
        .din(new_net_713),
        .dout(new_Jinkela_wire_1540)
    );

    spl2 new_Jinkela_splitter_209 (
        .a(_023_),
        .b(new_Jinkela_wire_1536),
        .c(new_Jinkela_wire_1537)
    );

    spl2 new_Jinkela_splitter_210 (
        .a(_213_),
        .b(new_Jinkela_wire_1538),
        .c(new_Jinkela_wire_1539)
    );

    bfr new_Jinkela_buffer_1012 (
        .din(_225_),
        .dout(new_Jinkela_wire_1546)
    );

    bfr new_Jinkela_buffer_1009 (
        .din(_198_),
        .dout(new_Jinkela_wire_1541)
    );

    or_bi _408_ (
        .a(_019_),
        .b(_018_),
        .c(_020_)
    );

    spl2 new_Jinkela_splitter_213 (
        .a(_242_),
        .b(new_Jinkela_wire_1554),
        .c(new_Jinkela_wire_1555)
    );

    bfr new_Jinkela_buffer_1010 (
        .din(new_Jinkela_wire_1541),
        .dout(new_Jinkela_wire_1542)
    );

    bfr new_Jinkela_buffer_493 (
        .din(new_Jinkela_wire_642),
        .dout(new_Jinkela_wire_643)
    );

    bfr new_Jinkela_buffer_133 (
        .din(new_Jinkela_wire_173),
        .dout(new_Jinkela_wire_174)
    );

    bfr new_Jinkela_buffer_66 (
        .din(new_Jinkela_wire_87),
        .dout(new_Jinkela_wire_88)
    );

    bfr new_Jinkela_buffer_478 (
        .din(new_Jinkela_wire_619),
        .dout(new_Jinkela_wire_620)
    );

    bfr new_Jinkela_buffer_85 (
        .din(new_Jinkela_wire_114),
        .dout(new_Jinkela_wire_115)
    );

    bfr new_Jinkela_buffer_514 (
        .din(new_Jinkela_wire_671),
        .dout(new_Jinkela_wire_672)
    );

    bfr new_Jinkela_buffer_67 (
        .din(new_Jinkela_wire_88),
        .dout(new_Jinkela_wire_89)
    );

    bfr new_Jinkela_buffer_479 (
        .din(new_Jinkela_wire_620),
        .dout(new_Jinkela_wire_621)
    );

    spl2 new_Jinkela_splitter_21 (
        .a(N93),
        .b(new_Jinkela_wire_243),
        .c(new_Jinkela_wire_245)
    );

    bfr new_Jinkela_buffer_494 (
        .din(new_Jinkela_wire_643),
        .dout(new_Jinkela_wire_644)
    );

    bfr new_Jinkela_buffer_134 (
        .din(new_Jinkela_wire_179),
        .dout(new_Jinkela_wire_180)
    );

    bfr new_Jinkela_buffer_68 (
        .din(new_Jinkela_wire_89),
        .dout(new_Jinkela_wire_90)
    );

    bfr new_Jinkela_buffer_480 (
        .din(new_Jinkela_wire_621),
        .dout(new_Jinkela_wire_622)
    );

    bfr new_Jinkela_buffer_86 (
        .din(new_Jinkela_wire_115),
        .dout(new_Jinkela_wire_116)
    );

    bfr new_Jinkela_buffer_69 (
        .din(new_Jinkela_wire_90),
        .dout(new_Jinkela_wire_91)
    );

    bfr new_Jinkela_buffer_481 (
        .din(new_Jinkela_wire_622),
        .dout(new_Jinkela_wire_623)
    );

    bfr new_Jinkela_buffer_109 (
        .din(new_Jinkela_wire_146),
        .dout(new_Jinkela_wire_147)
    );

    bfr new_Jinkela_buffer_495 (
        .din(new_Jinkela_wire_644),
        .dout(new_Jinkela_wire_645)
    );

    bfr new_Jinkela_buffer_70 (
        .din(new_Jinkela_wire_91),
        .dout(new_Jinkela_wire_92)
    );

    bfr new_Jinkela_buffer_482 (
        .din(new_Jinkela_wire_623),
        .dout(new_Jinkela_wire_624)
    );

    bfr new_Jinkela_buffer_87 (
        .din(new_Jinkela_wire_116),
        .dout(new_Jinkela_wire_117)
    );

    bfr new_Jinkela_buffer_515 (
        .din(new_Jinkela_wire_672),
        .dout(new_Jinkela_wire_673)
    );

    bfr new_Jinkela_buffer_71 (
        .din(new_Jinkela_wire_92),
        .dout(new_Jinkela_wire_93)
    );

    bfr new_Jinkela_buffer_483 (
        .din(new_Jinkela_wire_624),
        .dout(new_Jinkela_wire_625)
    );

    bfr new_Jinkela_buffer_496 (
        .din(new_Jinkela_wire_645),
        .dout(new_Jinkela_wire_646)
    );

    bfr new_Jinkela_buffer_72 (
        .din(new_Jinkela_wire_93),
        .dout(new_Jinkela_wire_94)
    );

    bfr new_Jinkela_buffer_484 (
        .din(new_Jinkela_wire_625),
        .dout(new_Jinkela_wire_626)
    );

    bfr new_Jinkela_buffer_88 (
        .din(new_Jinkela_wire_117),
        .dout(new_Jinkela_wire_118)
    );

    bfr new_Jinkela_buffer_538 (
        .din(new_Jinkela_wire_703),
        .dout(new_Jinkela_wire_704)
    );

    bfr new_Jinkela_buffer_564 (
        .din(new_Jinkela_wire_732),
        .dout(new_Jinkela_wire_733)
    );

    bfr new_Jinkela_buffer_73 (
        .din(new_Jinkela_wire_94),
        .dout(new_Jinkela_wire_95)
    );

    spl2 new_Jinkela_splitter_53 (
        .a(new_Jinkela_wire_626),
        .b(new_Jinkela_wire_627),
        .c(new_Jinkela_wire_628)
    );

    bfr new_Jinkela_buffer_110 (
        .din(new_Jinkela_wire_147),
        .dout(new_Jinkela_wire_148)
    );

    bfr new_Jinkela_buffer_516 (
        .din(new_Jinkela_wire_673),
        .dout(new_Jinkela_wire_674)
    );

    or_bi _387_ (
        .a(new_Jinkela_wire_599),
        .b(new_Jinkela_wire_3),
        .c(_361_)
    );

    bfr new_Jinkela_buffer_74 (
        .din(new_Jinkela_wire_95),
        .dout(new_Jinkela_wire_96)
    );

    bfr new_Jinkela_buffer_497 (
        .din(new_Jinkela_wire_646),
        .dout(new_Jinkela_wire_647)
    );

    or_bi _365_ (
        .a(_338_),
        .b(_337_),
        .c(_339_)
    );

    bfr new_Jinkela_buffer_89 (
        .din(new_Jinkela_wire_118),
        .dout(new_Jinkela_wire_119)
    );

    bfr new_Jinkela_buffer_498 (
        .din(new_Jinkela_wire_647),
        .dout(new_Jinkela_wire_648)
    );

    or_bi _363_ (
        .a(new_Jinkela_wire_108),
        .b(new_Jinkela_wire_698),
        .c(_337_)
    );

    bfr new_Jinkela_buffer_75 (
        .din(new_Jinkela_wire_96),
        .dout(new_Jinkela_wire_97)
    );

    bfr new_Jinkela_buffer_593 (
        .din(N133),
        .dout(new_Jinkela_wire_769)
    );

    and_bi _364_ (
        .a(new_Jinkela_wire_105),
        .b(new_Jinkela_wire_702),
        .c(_338_)
    );

    bfr new_Jinkela_buffer_499 (
        .din(new_Jinkela_wire_648),
        .dout(new_Jinkela_wire_649)
    );

    or_ii _362_ (
        .a(new_Jinkela_wire_313),
        .b(new_Jinkela_wire_1056),
        .c(_336_)
    );

    or_bi _366_ (
        .a(new_Jinkela_wire_319),
        .b(new_Jinkela_wire_982),
        .c(_340_)
    );

    bfr new_Jinkela_buffer_76 (
        .din(new_Jinkela_wire_97),
        .dout(new_Jinkela_wire_98)
    );

    bfr new_Jinkela_buffer_517 (
        .din(new_Jinkela_wire_674),
        .dout(new_Jinkela_wire_675)
    );

    and_bi _370_ (
        .a(new_Jinkela_wire_1172),
        .b(new_Jinkela_wire_1591),
        .c(_344_)
    );

    bfr new_Jinkela_buffer_90 (
        .din(new_Jinkela_wire_119),
        .dout(new_Jinkela_wire_120)
    );

    bfr new_Jinkela_buffer_500 (
        .din(new_Jinkela_wire_649),
        .dout(new_Jinkela_wire_650)
    );

    or_bi _369_ (
        .a(new_Jinkela_wire_1173),
        .b(new_Jinkela_wire_1592),
        .c(_343_)
    );

    bfr new_Jinkela_buffer_77 (
        .din(new_Jinkela_wire_98),
        .dout(new_Jinkela_wire_99)
    );

    bfr new_Jinkela_buffer_539 (
        .din(new_Jinkela_wire_704),
        .dout(new_Jinkela_wire_705)
    );

    and_bi _367_ (
        .a(new_Jinkela_wire_318),
        .b(new_Jinkela_wire_981),
        .c(_341_)
    );

    bfr new_Jinkela_buffer_111 (
        .din(new_Jinkela_wire_148),
        .dout(new_Jinkela_wire_149)
    );

    bfr new_Jinkela_buffer_501 (
        .din(new_Jinkela_wire_650),
        .dout(new_Jinkela_wire_651)
    );

    spl2 new_Jinkela_splitter_8 (
        .a(new_Jinkela_wire_99),
        .b(new_Jinkela_wire_100),
        .c(new_Jinkela_wire_101)
    );

    bfr new_Jinkela_buffer_518 (
        .din(new_Jinkela_wire_675),
        .dout(new_Jinkela_wire_676)
    );

    and_bi _379_ (
        .a(new_Jinkela_wire_879),
        .b(new_Jinkela_wire_1099),
        .c(_353_)
    );

    or_bi _368_ (
        .a(_341_),
        .b(_340_),
        .c(_342_)
    );

    spl4L new_Jinkela_splitter_19 (
        .a(new_Jinkela_wire_210),
        .d(new_Jinkela_wire_211),
        .e(new_Jinkela_wire_212),
        .b(new_Jinkela_wire_213),
        .c(new_Jinkela_wire_214)
    );

    bfr new_Jinkela_buffer_502 (
        .din(new_Jinkela_wire_651),
        .dout(new_Jinkela_wire_652)
    );

    or_bi _371_ (
        .a(_344_),
        .b(_343_),
        .c(_345_)
    );

    bfr new_Jinkela_buffer_91 (
        .din(new_Jinkela_wire_120),
        .dout(new_Jinkela_wire_121)
    );

    bfr new_Jinkela_buffer_592 (
        .din(new_Jinkela_wire_767),
        .dout(new_Jinkela_wire_768)
    );

    or_bi _372_ (
        .a(new_Jinkela_wire_1385),
        .b(new_Jinkela_wire_1155),
        .c(_346_)
    );

    bfr new_Jinkela_buffer_92 (
        .din(new_Jinkela_wire_121),
        .dout(new_Jinkela_wire_122)
    );

    bfr new_Jinkela_buffer_503 (
        .din(new_Jinkela_wire_652),
        .dout(new_Jinkela_wire_653)
    );

    and_bi _373_ (
        .a(new_Jinkela_wire_1384),
        .b(new_Jinkela_wire_1154),
        .c(_347_)
    );

    bfr new_Jinkela_buffer_112 (
        .din(new_Jinkela_wire_149),
        .dout(new_Jinkela_wire_150)
    );

    bfr new_Jinkela_buffer_519 (
        .din(new_Jinkela_wire_676),
        .dout(new_Jinkela_wire_677)
    );

    and_bi _374_ (
        .a(_346_),
        .b(_347_),
        .c(_348_)
    );

    bfr new_Jinkela_buffer_93 (
        .din(new_Jinkela_wire_122),
        .dout(new_Jinkela_wire_123)
    );

    bfr new_Jinkela_buffer_504 (
        .din(new_Jinkela_wire_653),
        .dout(new_Jinkela_wire_654)
    );

    or_bb _375_ (
        .a(new_Jinkela_wire_140),
        .b(new_Jinkela_wire_72),
        .c(_349_)
    );

    bfr new_Jinkela_buffer_540 (
        .din(new_Jinkela_wire_705),
        .dout(new_Jinkela_wire_706)
    );

    bfr new_Jinkela_buffer_160 (
        .din(new_Jinkela_wire_208),
        .dout(new_Jinkela_wire_209)
    );

    and_bb _376_ (
        .a(new_Jinkela_wire_142),
        .b(new_Jinkela_wire_71),
        .c(_350_)
    );

    bfr new_Jinkela_buffer_94 (
        .din(new_Jinkela_wire_123),
        .dout(new_Jinkela_wire_124)
    );

    bfr new_Jinkela_buffer_505 (
        .din(new_Jinkela_wire_654),
        .dout(new_Jinkela_wire_655)
    );

    and_bi _377_ (
        .a(_349_),
        .b(_350_),
        .c(_351_)
    );

    bfr new_Jinkela_buffer_113 (
        .din(new_Jinkela_wire_150),
        .dout(new_Jinkela_wire_151)
    );

    bfr new_Jinkela_buffer_520 (
        .din(new_Jinkela_wire_677),
        .dout(new_Jinkela_wire_678)
    );

    or_bi _378_ (
        .a(new_Jinkela_wire_878),
        .b(new_Jinkela_wire_1100),
        .c(_352_)
    );

    bfr new_Jinkela_buffer_95 (
        .din(new_Jinkela_wire_124),
        .dout(new_Jinkela_wire_125)
    );

    bfr new_Jinkela_buffer_506 (
        .din(new_Jinkela_wire_655),
        .dout(new_Jinkela_wire_656)
    );

    or_bi _380_ (
        .a(_353_),
        .b(_352_),
        .c(_354_)
    );

    bfr new_Jinkela_buffer_135 (
        .din(new_Jinkela_wire_180),
        .dout(new_Jinkela_wire_181)
    );

    bfr new_Jinkela_buffer_565 (
        .din(new_Jinkela_wire_738),
        .dout(new_Jinkela_wire_739)
    );

    or_bi _381_ (
        .a(new_Jinkela_wire_1637),
        .b(new_Jinkela_wire_1292),
        .c(_355_)
    );

    bfr new_Jinkela_buffer_96 (
        .din(new_Jinkela_wire_125),
        .dout(new_Jinkela_wire_126)
    );

    bfr new_Jinkela_buffer_507 (
        .din(new_Jinkela_wire_656),
        .dout(new_Jinkela_wire_657)
    );

    and_bi _382_ (
        .a(new_Jinkela_wire_1636),
        .b(new_Jinkela_wire_1291),
        .c(_356_)
    );

    bfr new_Jinkela_buffer_114 (
        .din(new_Jinkela_wire_151),
        .dout(new_Jinkela_wire_152)
    );

    bfr new_Jinkela_buffer_521 (
        .din(new_Jinkela_wire_678),
        .dout(new_Jinkela_wire_679)
    );

    and_bi _383_ (
        .a(_355_),
        .b(_356_),
        .c(_357_)
    );

    bfr new_Jinkela_buffer_97 (
        .din(new_Jinkela_wire_126),
        .dout(new_Jinkela_wire_127)
    );

    bfr new_Jinkela_buffer_508 (
        .din(new_Jinkela_wire_657),
        .dout(new_Jinkela_wire_658)
    );

    or_bb _384_ (
        .a(new_Jinkela_wire_354),
        .b(new_Jinkela_wire_668),
        .c(_358_)
    );

    spl4L new_Jinkela_splitter_22 (
        .a(new_Jinkela_wire_245),
        .d(new_Jinkela_wire_246),
        .e(new_Jinkela_wire_247),
        .b(new_Jinkela_wire_248),
        .c(new_Jinkela_wire_249)
    );

    bfr new_Jinkela_buffer_541 (
        .din(new_Jinkela_wire_706),
        .dout(new_Jinkela_wire_707)
    );

    spl2 new_Jinkela_splitter_24 (
        .a(N1),
        .b(new_Jinkela_wire_277),
        .c(new_Jinkela_wire_279)
    );

    and_bb _385_ (
        .a(new_Jinkela_wire_350),
        .b(new_Jinkela_wire_667),
        .c(_359_)
    );

    bfr new_Jinkela_buffer_98 (
        .din(new_Jinkela_wire_127),
        .dout(new_Jinkela_wire_128)
    );

    bfr new_Jinkela_buffer_509 (
        .din(new_Jinkela_wire_658),
        .dout(new_Jinkela_wire_659)
    );

    and_bi _386_ (
        .a(_358_),
        .b(_359_),
        .c(_360_)
    );

endmodule
