module c3540(G1, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, G30, G31, G32, G33, G34, G35, G3519, G3520, G3521, G3522, G3523, G3524, G3525, G3526, G3527, G3528, G3529, G3530, G3531, G3532, G3533, G3534, G3535, G3536, G3537, G3538, G3539, G3540, G36, G37, G38, G39, G4, G40, G41, G42, G43, G44, G45, G46, G47, G48, G49, G5, G50, G6, G7, G8, G9);
	wire new_net_3102;
	wire new_net_2822;
	wire new_net_3367;
	wire new_net_2977;
	wire new_net_2390;
	wire new_net_2071;
	wire new_net_2151;
	wire new_net_1233;
	wire new_net_2112;
	wire new_net_2353;
	wire new_net_2048;
	wire new_net_2833;
	wire new_net_2537;
	wire new_net_1492;
	wire new_net_2081;
	wire new_net_2653;
	wire new_net_1360;
	wire new_net_3103;
	wire new_net_2406;
	wire new_net_3342;
	wire new_net_2624;
	wire new_net_2247;
	wire new_net_3247;
	wire new_net_2692;
	wire _0022_;
	wire _0064_;
	wire _0106_;
	wire _0148_;
	wire _0190_;
	wire _0232_;
	wire _0274_;
	wire _0316_;
	wire _0358_;
	wire _0400_;
	wire new_net_2226;
	wire new_net_2633;
	wire new_net_1538;
	wire new_net_3126;
	wire new_net_1005;
	wire new_net_1131;
	wire new_net_3245;
	wire new_net_3000;
	wire new_net_3037;
	wire new_net_2560;
	wire new_net_1188;
	wire new_net_153;
	wire new_net_192;
	wire new_net_297;
	wire new_net_489;
	wire new_net_648;
	wire new_net_684;
	wire new_net_753;
	wire new_net_1029;
	wire new_net_1059;
	wire new_net_1064;
	wire new_net_1760;
	wire new_net_1981;
	wire new_net_3251;
	wire new_net_2941;
	wire new_net_1181;
	wire new_net_2610;
	wire new_net_1660;
	wire new_net_1039;
	wire new_net_2023;
	wire new_net_2423;
	wire new_net_3257;
	wire new_net_3016;
	wire _0315_;
	wire new_net_2024;
	wire _0611_;
	wire _0149_;
	wire _0023_;
	wire _0065_;
	wire _0107_;
	wire _0191_;
	wire _0233_;
	wire _0275_;
	wire _0317_;
	wire _0359_;
	wire new_net_2322;
	wire new_net_2989;
	wire new_net_2190;
	wire new_net_2546;
	wire new_net_3388;
	wire new_net_3310;
	wire new_net_661;
	wire new_net_1779;
	wire new_net_1677;
	wire new_net_1389;
	wire new_net_3;
	wire new_net_134;
	wire new_net_227;
	wire new_net_596;
	wire new_net_701;
	wire new_net_872;
	wire new_net_941;
	wire new_net_1171;
	wire new_net_1536;
	wire new_net_1715;
	wire new_net_2596;
	wire new_net_3044;
	wire new_net_3272;
	wire new_net_3397;
	wire new_net_2784;
	wire new_net_1924;
	wire new_net_1849;
	wire new_net_1265;
	wire new_net_3068;
	wire new_net_3361;
	wire new_net_3285;
	wire new_net_3283;
	wire new_net_2858;
	wire new_net_3070;
	wire _0570_;
	wire _0150_;
	wire _0024_;
	wire _0066_;
	wire _0108_;
	wire _0192_;
	wire _0234_;
	wire _0276_;
	wire _0318_;
	wire _0360_;
	wire _0444_;
	wire _0159_;
	wire new_net_1420;
	wire new_net_1522;
	wire new_net_2078;
	wire new_net_3372;
	wire new_net_2217;
	wire _0176_;
	wire new_net_1290;
	wire new_net_916;
	wire new_net_1739;
	wire new_net_3418;
	wire new_net_1737;
	wire new_net_511;
	wire new_net_2838;
	wire _0485_;
	wire new_net_100;
	wire new_net_1497;
	wire new_net_2658;
	wire new_net_3116;
	wire new_net_154;
	wire new_net_298;
	wire new_net_490;
	wire new_net_754;
	wire new_net_1030;
	wire new_net_1767;
	wire new_net_2051;
	wire new_net_2137;
	wire new_net_2225;
	wire new_net_1445;
	wire new_net_3347;
	wire new_net_3207;
	wire _0526_;
	wire new_net_1048;
	wire new_net_3133;
	wire new_net_2374;
	wire new_net_1321;
	wire new_net_2477;
	wire new_net_756;
	wire new_net_3405;
	wire _0697_;
	wire _0193_;
	wire _0235_;
	wire _0277_;
	wire _0025_;
	wire _0067_;
	wire _0109_;
	wire _0151_;
	wire _0319_;
	wire _0361_;
	wire new_net_2020;
	wire new_net_2046;
	wire new_net_2994;
	wire new_net_2276;
	wire new_net_2616;
	wire new_net_2946;
	wire new_net_1352;
	wire new_net_2685;
	wire new_net_135;
	wire _0037_;
	wire new_net_597;
	wire new_net_702;
	wire new_net_804;
	wire _0322_;
	wire new_net_873;
	wire new_net_942;
	wire new_net_1719;
	wire new_net_1731;
	wire new_net_3080;
	wire new_net_2367;
	wire _0339_;
	wire new_net_2197;
	wire _0363_;
	wire new_net_2301;
	wire new_net_533;
	wire new_net_2551;
	wire _0356_;
	wire new_net_1747;
	wire _0530_;
	wire new_net_193;
	wire _0194_;
	wire _0236_;
	wire _0278_;
	wire _0026_;
	wire _0068_;
	wire _0110_;
	wire _0152_;
	wire _0320_;
	wire new_net_811;
	wire new_net_946;
	wire new_net_1383;
	wire new_net_2790;
	wire new_net_3179;
	wire _0404_;
	wire _0397_;
	wire new_net_818;
	wire new_net_1651;
	wire new_net_2601;
	wire new_net_3216;
	wire new_net_953;
	wire new_net_2315;
	wire _0421_;
	wire new_net_830;
	wire new_net_1196;
	wire new_net_1929;
	wire new_net_689;
	wire new_net_2313;
	wire new_net_1553;
	wire new_net_839;
	wire new_net_404;
	wire new_net_155;
	wire new_net_299;
	wire new_net_1013;
	wire new_net_1635;
	wire new_net_1859;
	wire new_net_1882;
	wire new_net_2317;
	wire new_net_2635;
	wire new_net_2651;
	wire new_net_696;
	wire new_net_846;
	wire new_net_1570;
	wire new_net_705;
	wire new_net_3379;
	wire new_net_2430;
	wire new_net_1568;
	wire new_net_3083;
	wire new_net_3238;
	wire new_net_712;
	wire new_net_3165;
	wire new_net_3203;
	wire new_net_2918;
	wire new_net_2582;
	wire _0489_;
	wire _0783_;
	wire new_net_102;
	wire _0657_;
	wire _0027_;
	wire _0069_;
	wire _0111_;
	wire _0195_;
	wire _0237_;
	wire _0279_;
	wire _0788_;
	wire new_net_2058;
	wire new_net_1914;
	wire new_net_2033;
	wire new_net_1439;
	wire new_net_3209;
	wire new_net_3352;
	wire new_net_3138;
	wire new_net_1868;
	wire new_net_136;
	wire new_net_580;
	wire new_net_598;
	wire new_net_703;
	wire new_net_805;
	wire new_net_943;
	wire new_net_997;
	wire new_net_1499;
	wire new_net_1681;
	wire new_net_1720;
	wire new_net_2482;
	wire new_net_2818;
	wire new_net_1412;
	wire new_net_3149;
	wire new_net_1793;
	wire new_net_1988;
	wire new_net_2491;
	wire new_net_2255;
	wire _0448_;
	wire _0742_;
	wire _0616_;
	wire _0028_;
	wire _0070_;
	wire _0112_;
	wire _0196_;
	wire _0238_;
	wire _0280_;
	wire _0154_;
	wire new_net_2539;
	wire new_net_2620;
	wire new_net_2770;
	wire new_net_3260;
	wire new_net_3338;
	wire new_net_2690;
	wire new_net_2298;
	wire new_net_2872;
	wire new_net_2087;
	wire new_net_2964;
	wire new_net_1757;
	wire new_net_156;
	wire new_net_300;
	wire new_net_48;
	wire new_net_405;
	wire new_net_840;
	wire new_net_1014;
	wire new_net_1208;
	wire new_net_1688;
	wire new_net_1865;
	wire new_net_2171;
	wire new_net_2202;
	wire new_net_2169;
	wire new_net_2556;
	wire _0095_;
	wire _0683_;
	wire new_net_1304;
	wire new_net_1505;
	wire new_net_1899;
	wire new_net_55;
	wire new_net_3099;
	wire new_net_2076;
	wire new_net_3184;
	wire new_net_1106;
	wire new_net_2174;
	wire new_net_1656;
	wire new_net_3221;
	wire new_net_2323;
	wire _0701_;
	wire _0575_;
	wire _0449_;
	wire _0743_;
	wire new_net_229;
	wire _0197_;
	wire _0239_;
	wire _0281_;
	wire _0029_;
	wire _0071_;
	wire new_net_494;
	wire new_net_1286;
	wire _0445_;
	wire new_net_2863;
	wire new_net_775;
	wire new_net_1065;
	wire new_net_3295;
	wire new_net_3199;
	wire _0177_;
	wire new_net_501;
	wire new_net_2462;
	wire new_net_1362;
	wire new_net_1672;
	wire new_net_2001;
	wire new_net_3058;
	wire new_net_3384;
	wire _0486_;
	wire new_net_1441;
	wire new_net_1943;
	wire new_net_3051;
	wire new_net_3301;
	wire new_net_137;
	wire new_net_581;
	wire new_net_599;
	wire new_net_704;
	wire new_net_890;
	wire new_net_944;
	wire new_net_998;
	wire new_net_520;
	wire new_net_1521;
	wire new_net_1573;
	wire new_net_2131;
	wire new_net_3120;
	wire new_net_2628;
	wire new_net_3170;
	wire new_net_2034;
	wire new_net_2224;
	wire new_net_2735;
	wire new_net_1317;
	wire new_net_2923;
	wire new_net_2062;
	wire new_net_2587;
	wire new_net_2695;
	wire _0527_;
	wire new_net_2634;
	wire new_net_3092;
	wire new_net_1109;
	wire new_net_1918;
	wire new_net_2446;
	wire new_net_1090;
	wire new_net_1682;
	wire _0534_;
	wire new_net_195;
	wire _0702_;
	wire _0198_;
	wire _0240_;
	wire _0282_;
	wire _0030_;
	wire _0072_;
	wire _0114_;
	wire _0156_;
	wire new_net_3145;
	wire new_net_2710;
	wire new_net_1348;
	wire new_net_3079;
	wire new_net_3334;
	wire new_net_1100;
	wire new_net_1692;
	wire new_net_2573;
	wire new_net_406;
	wire new_net_49;
	wire new_net_103;
	wire new_net_157;
	wire new_net_301;
	wire new_net_841;
	wire new_net_1015;
	wire new_net_1032;
	wire _0323_;
	wire new_net_1253;
	wire new_net_1173;
	wire new_net_2958;
	wire new_net_2929;
	wire new_net_2775;
	wire new_net_1201;
	wire new_net_2228;
	wire _0364_;
	wire new_net_1379;
	wire new_net_2879;
	wire _0357_;
	wire new_net_1083;
	wire _0493_;
	wire _0787_;
	wire _0661_;
	wire _0535_;
	wire _0199_;
	wire _0241_;
	wire _0157_;
	wire _0031_;
	wire _0381_;
	wire _0073_;
	wire new_net_1950;
	wire new_net_2091;
	wire new_net_2469;
	wire new_net_2096;
	wire _0405_;
	wire new_net_822;
	wire new_net_551;
	wire _0398_;
	wire _0422_;
	wire new_net_3009;
	wire new_net_2248;
	wire new_net_3191;
	wire new_net_2756;
	wire new_net_138;
	wire new_net_582;
	wire new_net_600;
	wire new_net_891;
	wire new_net_945;
	wire new_net_1210;
	wire new_net_1637;
	wire new_net_1671;
	wire new_net_1862;
	wire new_net_1945;
	wire _0724_;
	wire new_net_1280;
	wire new_net_3110;
	wire new_net_1527;
	wire _0765_;
	wire new_net_1435;
	wire _0452_;
	wire _0662_;
	wire _0620_;
	wire _0746_;
	wire _0494_;
	wire _0032_;
	wire _0074_;
	wire _0116_;
	wire _0158_;
	wire _0200_;
	wire new_net_999;
	wire new_net_1809;
	wire new_net_2006;
	wire new_net_2507;
	wire new_net_2526;
	wire new_net_2729;
	wire new_net_3056;
	wire new_net_3086;
	wire new_net_3306;
	wire new_net_1006;
	wire new_net_1311;
	wire new_net_1135;
	wire new_net_2340;
	wire new_net_2474;
	wire new_net_2925;
	wire new_net_3175;
	wire _0242_;
	wire new_net_3402;
	wire new_net_2740;
	wire new_net_403;
	wire new_net_2789;
	wire new_net_1852;
	wire new_net_230;
	wire new_net_302;
	wire new_net_50;
	wire new_net_104;
	wire new_net_158;
	wire new_net_407;
	wire new_net_1022;
	wire new_net_1033;
	wire new_net_1052;
	wire new_net_1823;
	wire new_net_2718;
	wire new_net_2347;
	wire _0283_;
	wire new_net_1870;
	wire new_net_3075;
	wire _0568_;
	wire new_net_3330;
	wire new_net_2643;
	wire new_net_1905;
	wire new_net_3328;
	wire new_net_1040;
	wire new_net_2715;
	wire new_net_3255;
	wire new_net_2117;
	wire _0705_;
	wire _0579_;
	wire _0453_;
	wire _0747_;
	wire _0621_;
	wire _0495_;
	wire _0789_;
	wire _0201_;
	wire _0243_;
	wire _0285_;
	wire new_net_1699;
	wire new_net_1938;
	wire new_net_3156;
	wire new_net_662;
	wire new_net_139;
	wire new_net_196;
	wire _0079_;
	wire new_net_601;
	wire new_net_652;
	wire new_net_892;
	wire new_net_1213;
	wire new_net_1884;
	wire new_net_2013;
	wire new_net_2232;
	wire new_net_2470;
	wire new_net_2884;
	wire new_net_3039;
	wire _0684_;
	wire new_net_2379;
	wire new_net_1619;
	wire new_net_3270;
	wire new_net_1206;
	wire new_net_2101;
	wire new_net_2281;
	wire new_net_1340;
	wire new_net_2814;
	wire new_net_1398;
	wire new_net_3354;
	wire new_net_2352;
	wire _0706_;
	wire _0580_;
	wire _0137_;
	wire _0454_;
	wire _0748_;
	wire _0034_;
	wire _0076_;
	wire _0118_;
	wire _0160_;
	wire _0202_;
	wire new_net_1795;
	wire new_net_2427;
	wire new_net_3014;
	wire _0446_;
	wire new_net_3196;
	wire new_net_2761;
	wire new_net_3228;
	wire new_net_1150;
	wire new_net_1799;
	wire new_net_2649;
	wire _0463_;
	wire new_net_3025;
	wire new_net_512;
	wire new_net_3115;
	wire _0487_;
	wire new_net_101;
	wire new_net_408;
	wire new_net_51;
	wire new_net_159;
	wire new_net_231;
	wire new_net_303;
	wire new_net_876;
	wire new_net_1034;
	wire new_net_1053;
	wire new_net_1084;
	wire new_net_1193;
	wire new_net_1371;
	wire new_net_1429;
	wire new_net_1837;
	wire new_net_2057;
	wire new_net_2466;
	wire new_net_2059;
	wire new_net_2809;
	wire new_net_2030;
	wire _0528_;
	wire new_net_3033;
	wire new_net_2512;
	wire new_net_1580;
	wire new_net_1895;
	wire new_net_1978;
	wire new_net_1101;
	wire new_net_2930;
	wire new_net_2747;
	wire _0665_;
	wire _0539_;
	wire _0707_;
	wire _0581_;
	wire _0035_;
	wire _0077_;
	wire _0119_;
	wire _0161_;
	wire _0203_;
	wire _0245_;
	wire new_net_757;
	wire new_net_1583;
	wire new_net_1647;
	wire new_net_1402;
	wire new_net_2673;
	wire new_net_2794;
	wire new_net_1769;
	wire new_net_2568;
	wire new_net_2980;
	wire new_net_1097;
	wire new_net_1875;
	wire new_net_2905;
	wire new_net_197;
	wire new_net_653;
	wire new_net_893;
	wire new_net_2487;
	wire new_net_2497;
	wire new_net_2521;
	wire new_net_1770;
	wire new_net_2498;
	wire new_net_2533;
	wire new_net_2627;
	wire _0324_;
	wire new_net_1601;
	wire new_net_2258;
	wire new_net_1105;
	wire new_net_3161;
	wire new_net_2843;
	wire _0341_;
	wire new_net_1704;
	wire new_net_2262;
	wire new_net_2332;
	wire _0365_;
	wire new_net_1842;
	wire new_net_2165;
	wire new_net_2302;
	wire new_net_534;
	wire _0624_;
	wire _0498_;
	wire _0792_;
	wire new_net_1054;
	wire _0666_;
	wire _0540_;
	wire _0036_;
	wire _0078_;
	wire _0120_;
	wire _0162_;
	wire new_net_3274;
	wire _0382_;
	wire new_net_2704;
	wire new_net_947;
	wire _0406_;
	wire new_net_2891;
	wire new_net_1458;
	wire new_net_1951;
	wire new_net_2973;
	wire _0399_;
	wire new_net_819;
	wire new_net_2386;
	wire new_net_2067;
	wire new_net_2706;
	wire new_net_954;
	wire new_net_2889;
	wire new_net_2147;
	wire new_net_2860;
	wire _0423_;
	wire new_net_1725;
	wire _0708_;
	wire new_net_690;
	wire new_net_1276;
	wire new_net_160;
	wire new_net_232;
	wire new_net_304;
	wire new_net_409;
	wire new_net_808;
	wire new_net_877;
	wire new_net_1035;
	wire new_net_1334;
	wire new_net_1673;
	wire new_net_1689;
	wire new_net_1729;
	wire new_net_2318;
	wire _0725_;
	wire new_net_2827;
	wire new_net_2357;
	wire new_net_847;
	wire new_net_3021;
	wire _0749_;
	wire new_net_706;
	wire new_net_2431;
	wire new_net_3048;
	wire new_net_1431;
	wire new_net_854;
	wire new_net_2766;
	wire new_net_1830;
	wire new_net_2805;
	wire _0766_;
	wire new_net_713;
	wire new_net_3027;
	wire _0583_;
	wire _0457_;
	wire _0751_;
	wire _0625_;
	wire _0499_;
	wire _0793_;
	wire _0667_;
	wire _0541_;
	wire _0205_;
	wire _0247_;
	wire _0790_;
	wire new_net_1307;
	wire new_net_1365;
	wire new_net_3122;
	wire _0219_;
	wire new_net_1510;
	wire new_net_2016;
	wire new_net_3320;
	wire new_net_2517;
	wire new_net_198;
	wire new_net_654;
	wire new_net_759;
	wire new_net_894;
	wire new_net_1528;
	wire new_net_1540;
	wire new_net_1631;
	wire new_net_1792;
	wire new_net_1891;
	wire new_net_2041;
	wire new_net_2138;
	wire new_net_2937;
	wire new_net_2606;
	wire new_net_2935;
	wire _0284_;
	wire new_net_2752;
	wire _0569_;
	wire new_net_1961;
	wire new_net_1764;
	wire new_net_3411;
	wire new_net_2358;
	wire new_net_3321;
	wire _0710_;
	wire _0584_;
	wire _0458_;
	wire _0752_;
	wire _0626_;
	wire _0500_;
	wire _0794_;
	wire new_net_106;
	wire _0038_;
	wire _0080_;
	wire _0610_;
	wire new_net_1880;
	wire _0603_;
	wire new_net_1968;
	wire new_net_2292;
	wire new_net_2910;
	wire new_net_1608;
	wire new_net_1776;
	wire new_net_1997;
	wire new_net_2503;
	wire new_net_3420;
	wire new_net_2660;
	wire new_net_2127;
	wire _0644_;
	wire new_net_1711;
	wire new_net_2592;
	wire new_net_2168;
	wire new_net_3268;
	wire new_net_161;
	wire new_net_233;
	wire new_net_305;
	wire _0668_;
	wire new_net_809;
	wire new_net_878;
	wire new_net_1001;
	wire new_net_1036;
	wire new_net_1207;
	wire new_net_1639;
	wire new_net_1545;
	wire new_net_2780;
	wire new_net_2852;
	wire new_net_3357;
	wire _0685_;
	wire new_net_2450;
	wire new_net_1753;
	wire new_net_1952;
	wire new_net_3006;
	wire new_net_56;
	wire new_net_1394;
	wire new_net_3279;
	wire new_net_3004;
	wire _0121_;
	wire new_net_2932;
	wire new_net_2896;
	wire new_net_2823;
	wire new_net_3368;
	wire _0669_;
	wire _0543_;
	wire _0711_;
	wire new_net_141;
	wire _0585_;
	wire _0459_;
	wire _0753_;
	wire _0627_;
	wire _0165_;
	wire _0039_;
	wire new_net_1270;
	wire new_net_2072;
	wire new_net_2152;
	wire new_net_495;
	wire new_net_2113;
	wire _0447_;
	wire new_net_2459;
	wire new_net_776;
	wire new_net_2834;
	wire _0179_;
	wire new_net_2538;
	wire new_net_2082;
	wire new_net_2433;
	wire new_net_2654;
	wire _0464_;
	wire new_net_1425;
	wire new_net_1835;
	wire new_net_2407;
	wire new_net_3343;
	wire _0488_;
	wire new_net_199;
	wire new_net_655;
	wire new_net_760;
	wire new_net_895;
	wire new_net_1212;
	wire new_net_1798;
	wire new_net_1845;
	wire new_net_1892;
	wire new_net_1923;
	wire new_net_2028;
	wire new_net_2265;
	wire new_net_521;
	wire _0505_;
	wire new_net_1539;
	wire new_net_3127;
	wire _0529_;
	wire _0522_;
	wire new_net_1450;
	wire new_net_3246;
	wire new_net_3096;
	wire _0546_;
	wire _0628_;
	wire _0502_;
	wire _0796_;
	wire new_net_107;
	wire _0670_;
	wire _0544_;
	wire new_net_53;
	wire new_net_410;
	wire _0712_;
	wire _0586_;
	wire new_net_888;
	wire new_net_2561;
	wire _0563_;
	wire new_net_3252;
	wire new_net_1856;
	wire new_net_2942;
	wire new_net_2797;
	wire new_net_2611;
	wire new_net_3234;
	wire new_net_162;
	wire new_net_306;
	wire new_net_585;
	wire new_net_708;
	wire new_net_1002;
	wire new_net_1037;
	wire new_net_1886;
	wire new_net_2021;
	wire new_net_2025;
	wire _0040_;
	wire new_net_2363;
	wire _0325_;
	wire new_net_1299;
	wire new_net_1772;
	wire new_net_1940;
	wire new_net_2191;
	wire new_net_2326;
	wire _0342_;
	wire new_net_588;
	wire new_net_1205;
	wire new_net_2542;
	wire new_net_2547;
	wire new_net_1257;
	wire new_net_3389;
	wire new_net_3311;
	wire new_net_1780;
	wire _0366_;
	wire new_net_3426;
	wire new_net_1613;
	wire new_net_1678;
	wire _0587_;
	wire _0461_;
	wire _0755_;
	wire _0629_;
	wire _0503_;
	wire _0797_;
	wire _0671_;
	wire _0545_;
	wire _0713_;
	wire new_net_142;
	wire new_net_1260;
	wire new_net_1454;
	wire new_net_2063;
	wire new_net_2471;
	wire _0383_;
	wire new_net_1716;
	wire new_net_2597;
	wire new_net_3398;
	wire _0407_;
	wire new_net_823;
	wire new_net_2785;
	wire new_net_1925;
	wire new_net_2173;
	wire new_net_1330;
	wire new_net_1549;
	wire new_net_3286;
	wire new_net_3362;
	wire _0424_;
	wire new_net_3284;
	wire _0709_;
	wire new_net_200;
	wire new_net_497;
	wire new_net_656;
	wire new_net_692;
	wire new_net_896;
	wire new_net_1653;
	wire new_net_1724;
	wire new_net_1761;
	wire new_net_1958;
	wire new_net_2351;
	wire new_net_2859;
	wire new_net_3071;
	wire _0441_;
	wire new_net_1595;
	wire new_net_2398;
	wire new_net_2901;
	wire _0726_;
	wire new_net_3373;
	wire new_net_642;
	wire new_net_3393;
	wire new_net_3415;
	wire _0750_;
	wire new_net_2218;
	wire new_net_1740;
	wire new_net_2914;
	wire new_net_2578;
	wire new_net_1361;
	wire new_net_1738;
	wire _0714_;
	wire _0588_;
	wire _0462_;
	wire _0756_;
	wire new_net_234;
	wire new_net_411;
	wire _0630_;
	wire _0504_;
	wire _0672_;
	wire new_net_54;
	wire _0791_;
	wire new_net_1000;
	wire new_net_1838;
	wire new_net_2029;
	wire new_net_2162;
	wire new_net_3348;
	wire new_net_3030;
	wire new_net_2861;
	wire new_net_2031;
	wire _0220_;
	wire new_net_3134;
	wire new_net_2985;
	wire _0244_;
	wire new_net_1016;
	wire new_net_163;
	wire new_net_307;
	wire new_net_586;
	wire new_net_604;
	wire new_net_709;
	wire new_net_1038;
	wire new_net_1209;
	wire new_net_1502;
	wire new_net_1584;
	wire new_net_1771;
	wire new_net_1023;
	wire new_net_3406;
	wire new_net_1133;
	wire new_net_2277;
	wire new_net_1246;
	wire new_net_2452;
	wire new_net_1906;
	wire new_net_2949;
	wire new_net_2617;
	wire _0001_;
	wire _0043_;
	wire _0085_;
	wire _0127_;
	wire _0211_;
	wire _0253_;
	wire _0295_;
	wire _0169_;
	wire _0337_;
	wire _0379_;
	wire new_net_1666;
	wire new_net_2179;
	wire new_net_1141;
	wire new_net_1147;
	wire new_net_2686;
	wire new_net_2368;
	wire _0652_;
	wire new_net_2198;
	wire new_net_663;
	wire new_net_108;
	wire new_net_201;
	wire new_net_498;
	wire new_net_657;
	wire new_net_693;
	wire new_net_897;
	wire _0081_;
	wire new_net_1020;
	wire new_net_1158;
	wire new_net_1590;
	wire new_net_2552;
	wire new_net_1390;
	wire new_net_3316;
	wire new_net_3180;
	wire _0098_;
	wire new_net_1788;
	wire _0122_;
	wire new_net_1266;
	wire new_net_1652;
	wire new_net_3217;
	wire new_net_2316;
	wire _0002_;
	wire _0044_;
	wire _0086_;
	wire _0128_;
	wire _0212_;
	wire _0254_;
	wire _0296_;
	wire _0170_;
	wire _0338_;
	wire _0380_;
	wire _0139_;
	wire new_net_1554;
	wire new_net_3291;
	wire _0163_;
	wire new_net_1421;
	wire new_net_2052;
	wire new_net_2354;
	wire new_net_2720;
	wire new_net_3380;
	wire new_net_2288;
	wire _0180_;
	wire new_net_1291;
	wire new_net_918;
	wire new_net_1250;
	wire new_net_3297;
	wire new_net_513;
	wire new_net_3239;
	wire new_net_164;
	wire new_net_308;
	wire new_net_587;
	wire new_net_605;
	wire new_net_710;
	wire new_net_950;
	wire new_net_1183;
	wire new_net_1530;
	wire new_net_1797;
	wire new_net_1808;
	wire new_net_2583;
	wire new_net_2919;
	wire new_net_3204;
	wire new_net_3063;
	wire _0506_;
	wire new_net_1446;
	wire new_net_1915;
	wire new_net_2411;
	wire new_net_2998;
	wire new_net_3210;
	wire new_net_1947;
	wire new_net_1195;
	wire new_net_1322;
	wire new_net_1643;
	wire _0465_;
	wire _0759_;
	wire _0213_;
	wire _0255_;
	wire _0297_;
	wire _0045_;
	wire _0003_;
	wire _0087_;
	wire _0129_;
	wire _0171_;
	wire _0547_;
	wire new_net_758;
	wire new_net_3139;
	wire new_net_2483;
	wire new_net_2143;
	wire new_net_1765;
	wire new_net_2569;
	wire new_net_3150;
	wire new_net_1096;
	wire new_net_1869;
	wire new_net_109;
	wire new_net_202;
	wire new_net_898;
	wire new_net_1021;
	wire new_net_1077;
	wire new_net_1132;
	wire new_net_1211;
	wire new_net_1252;
	wire new_net_1353;
	wire new_net_1785;
	wire new_net_1934;
	wire new_net_2256;
	wire _0041_;
	wire new_net_2954;
	wire new_net_2771;
	wire new_net_3339;
	wire _0326_;
	wire new_net_2621;
	wire _0058_;
	wire new_net_2299;
	wire _0343_;
	wire new_net_2370;
	wire new_net_2873;
	wire new_net_2088;
	wire new_net_2965;
	wire _0367_;
	wire new_net_806;
	wire _0718_;
	wire _0214_;
	wire _0256_;
	wire _0298_;
	wire _0046_;
	wire _0004_;
	wire _0088_;
	wire _0130_;
	wire _0172_;
	wire _0340_;
	wire new_net_2166;
	wire new_net_3324;
	wire new_net_2307;
	wire new_net_2665;
	wire new_net_2967;
	wire _0384_;
	wire new_net_1384;
	wire new_net_948;
	wire new_net_2557;
	wire new_net_1506;
	wire _0408_;
	wire new_net_1900;
	wire new_net_3042;
	wire new_net_955;
	wire new_net_3185;
	wire new_net_165;
	wire new_net_309;
	wire new_net_606;
	wire new_net_691;
	wire new_net_711;
	wire new_net_831;
	wire new_net_951;
	wire new_net_1071;
	wire new_net_1176;
	wire new_net_1258;
	wire new_net_1556;
	wire new_net_1907;
	wire new_net_3222;
	wire new_net_2680;
	wire new_net_848;
	wire new_net_3296;
	wire new_net_707;
	wire new_net_2866;
	wire new_net_3200;
	wire new_net_2463;
	wire new_net_855;
	wire new_net_2002;
	wire _0551_;
	wire _0425_;
	wire _0215_;
	wire _0257_;
	wire _0299_;
	wire _0173_;
	wire _0005_;
	wire _0047_;
	wire _0089_;
	wire _0131_;
	wire new_net_1944;
	wire new_net_2978;
	wire new_net_3052;
	wire _0204_;
	wire new_net_2132;
	wire new_net_1574;
	wire new_net_3302;
	wire new_net_2629;
	wire new_net_3171;
	wire new_net_2736;
	wire new_net_1440;
	wire new_net_2924;
	wire new_net_2588;
	wire new_net_3093;
	wire new_net_2270;
	wire new_net_2696;
	wire new_net_1850;
	wire new_net_2447;
	wire new_net_110;
	wire new_net_236;
	wire new_net_812;
	wire new_net_881;
	wire new_net_2142;
	wire new_net_2253;
	wire new_net_2815;
	wire new_net_3010;
	wire new_net_1683;
	wire new_net_3022;
	wire _0262_;
	wire new_net_1954;
	wire new_net_3146;
	wire _0286_;
	wire new_net_2711;
	wire _0571_;
	wire new_net_2489;
	wire new_net_1413;
	wire new_net_3335;
	wire _0510_;
	wire _0678_;
	wire _0006_;
	wire _0048_;
	wire _0090_;
	wire _0132_;
	wire _0174_;
	wire _0216_;
	wire _0258_;
	wire _0300_;
	wire _0612_;
	wire new_net_1099;
	wire new_net_1775;
	wire new_net_2574;
	wire new_net_2869;
	wire new_net_2961;
	wire new_net_2959;
	wire new_net_2327;
	wire _0653_;
	wire new_net_2880;
	wire new_net_166;
	wire new_net_310;
	wire new_net_763;
	wire new_net_832;
	wire new_net_952;
	wire new_net_1633;
	wire new_net_1655;
	wire new_net_1763;
	wire new_net_2089;
	wire _0082_;
	wire new_net_2375;
	wire new_net_2092;
	wire new_net_2778;
	wire new_net_1262;
	wire new_net_3066;
	wire new_net_2097;
	wire new_net_2205;
	wire _0099_;
	wire new_net_57;
	wire _0123_;
	wire new_net_2522;
	wire _0469_;
	wire _0763_;
	wire _0637_;
	wire _0511_;
	wire _0217_;
	wire _0259_;
	wire _0301_;
	wire _0049_;
	wire _0007_;
	wire _0091_;
	wire _0140_;
	wire new_net_2757;
	wire new_net_3192;
	wire new_net_1836;
	wire new_net_3370;
	wire _0164_;
	wire new_net_496;
	wire new_net_1287;
	wire new_net_1345;
	wire new_net_2681;
	wire new_net_1733;
	wire new_net_1178;
	wire new_net_1561;
	wire new_net_3111;
	wire new_net_2990;
	wire _0466_;
	wire new_net_237;
	wire new_net_813;
	wire new_net_882;
	wire new_net_1177;
	wire new_net_1504;
	wire _0490_;
	wire new_net_1442;
	wire new_net_1885;
	wire new_net_2269;
	wire new_net_2422;
	wire new_net_2159;
	wire new_net_2508;
	wire new_net_2730;
	wire new_net_522;
	wire new_net_2007;
	wire new_net_3242;
	wire new_net_1576;
	wire new_net_2848;
	wire _0507_;
	wire new_net_3307;
	wire new_net_1318;
	wire new_net_1376;
	wire new_net_2668;
	wire _0531_;
	wire new_net_2475;
	wire new_net_2743;
	wire new_net_2926;
	wire new_net_3176;
	wire new_net_3403;
	wire new_net_2741;
	wire _0722_;
	wire _0596_;
	wire _0470_;
	wire _0764_;
	wire _0218_;
	wire _0260_;
	wire _0302_;
	wire _0050_;
	wire _0008_;
	wire _0092_;
	wire _0548_;
	wire new_net_880;
	wire new_net_1982;
	wire new_net_2895;
	wire new_net_889;
	wire new_net_1955;
	wire new_net_2348;
	wire new_net_1871;
	wire new_net_3076;
	wire new_net_1685;
	wire new_net_2564;
	wire new_net_1229;
	wire new_net_3331;
	wire new_net_143;
	wire new_net_2644;
	wire new_net_2453;
	wire new_net_3329;
	wire new_net_1349;
	wire new_net_1407;
	wire new_net_2716;
	wire new_net_2494;
	wire new_net_167;
	wire new_net_311;
	wire new_net_764;
	wire new_net_1165;
	wire new_net_1197;
	wire new_net_1259;
	wire new_net_1591;
	wire new_net_1705;
	wire new_net_1717;
	wire new_net_1806;
	wire new_net_2118;
	wire new_net_2492;
	wire _0042_;
	wire new_net_1098;
	wire new_net_3157;
	wire _0327_;
	wire new_net_1700;
	wire _0059_;
	wire new_net_1773;
	wire _0344_;
	wire new_net_589;
	wire new_net_727;
	wire new_net_2231;
	wire _0429_;
	wire _0723_;
	wire new_net_147;
	wire _0597_;
	wire _0261_;
	wire _0303_;
	wire _0009_;
	wire _0051_;
	wire _0093_;
	wire _0135_;
	wire _0368_;
	wire new_net_2700;
	wire new_net_2545;
	wire new_net_2969;
	wire new_net_3345;
	wire _0385_;
	wire new_net_2382;
	wire new_net_2885;
	wire new_net_2380;
	wire _0409_;
	wire new_net_824;
	wire new_net_1721;
	wire _0694_;
	wire new_net_2104;
	wire new_net_2333;
	wire new_net_2102;
	wire new_net_2282;
	wire new_net_238;
	wire _0426_;
	wire new_net_814;
	wire new_net_1041;
	wire new_net_1163;
	wire new_net_1216;
	wire new_net_1532;
	wire new_net_1541;
	wire new_net_1735;
	wire new_net_1778;
	wire new_net_2527;
	wire new_net_1860;
	wire new_net_3017;
	wire new_net_3045;
	wire new_net_2284;
	wire new_net_2428;
	wire new_net_3105;
	wire new_net_1281;
	wire new_net_1572;
	wire new_net_1833;
	wire new_net_2762;
	wire new_net_3229;
	wire new_net_3118;
	wire new_net_2156;
	wire _0682_;
	wire _0556_;
	wire new_net_59;
	wire _0430_;
	wire new_net_416;
	wire _0010_;
	wire _0052_;
	wire _0094_;
	wire _0136_;
	wire _0178_;
	wire new_net_1533;
	wire new_net_1436;
	wire new_net_1911;
	wire new_net_2995;
	wire new_net_2467;
	wire new_net_458;
	wire new_net_1056;
	wire new_net_3423;
	wire new_net_2060;
	wire new_net_1746;
	wire new_net_2412;
	wire _0222_;
	wire new_net_1312;
	wire new_net_2513;
	wire _0246_;
	wire new_net_1017;
	wire new_net_1820;
	wire new_net_168;
	wire new_net_312;
	wire new_net_1236;
	wire new_net_1592;
	wire new_net_1787;
	wire new_net_1896;
	wire new_net_2038;
	wire new_net_2108;
	wire new_net_2242;
	wire new_net_2252;
	wire new_net_2602;
	wire new_net_2748;
	wire new_net_2931;
	wire new_net_1024;
	wire new_net_1930;
	wire new_net_2591;
	wire new_net_412;
	wire new_net_2795;
	wire new_net_3325;
	wire _0287_;
	wire new_net_1242;
	wire _0572_;
	wire new_net_2981;
	wire _0304_;
	wire new_net_1876;
	wire _0767_;
	wire _0431_;
	wire _0641_;
	wire new_net_148;
	wire _0515_;
	wire _0557_;
	wire _0221_;
	wire _0305_;
	wire _0263_;
	wire _0011_;
	wire _0589_;
	wire new_net_2180;
	wire _0613_;
	wire new_net_2906;
	wire new_net_2499;
	wire new_net_2324;
	wire new_net_1602;
	wire new_net_1142;
	wire new_net_3038;
	wire new_net_2844;
	wire new_net_3162;
	wire _0654_;
	wire new_net_1498;
	wire new_net_239;
	wire new_net_851;
	wire new_net_664;
	wire new_net_1007;
	wire new_net_1042;
	wire new_net_1094;
	wire new_net_1686;
	wire new_net_1726;
	wire new_net_1744;
	wire new_net_1175;
	wire new_net_1843;
	wire new_net_3353;
	wire _0083_;
	wire new_net_1501;
	wire new_net_2238;
	wire new_net_3275;
	wire new_net_1058;
	wire _0100_;
	wire new_net_2892;
	wire new_net_2819;
	wire new_net_2974;
	wire _0124_;
	wire new_net_2387;
	wire new_net_2068;
	wire new_net_2707;
	wire _0600_;
	wire _0474_;
	wire _0768_;
	wire _0642_;
	wire _0516_;
	wire new_net_417;
	wire _0054_;
	wire _0012_;
	wire _0096_;
	wire _0138_;
	wire new_net_1283;
	wire new_net_1341;
	wire _0141_;
	wire new_net_1730;
	wire new_net_2109;
	wire new_net_1825;
	wire new_net_1075;
	wire new_net_2287;
	wire new_net_2534;
	wire new_net_2800;
	wire new_net_2828;
	wire _0450_;
	wire new_net_1483;
	wire new_net_2432;
	wire new_net_2802;
	wire _0467_;
	wire new_net_169;
	wire new_net_205;
	wire new_net_313;
	wire new_net_502;
	wire new_net_514;
	wire new_net_697;
	wire new_net_1161;
	wire new_net_1223;
	wire _0491_;
	wire new_net_1831;
	wire new_net_2222;
	wire new_net_2806;
	wire new_net_1743;
	wire new_net_1372;
	wire new_net_3123;
	wire new_net_2271;
	wire new_net_3428;
	wire _0508_;
	wire new_net_1227;
	wire new_net_2035;
	wire new_net_1812;
	wire _0532_;
	wire new_net_3034;
	wire _0433_;
	wire _0727_;
	wire _0601_;
	wire _0475_;
	wire _0769_;
	wire _0643_;
	wire _0181_;
	wire _0055_;
	wire _0013_;
	wire _0097_;
	wire _0549_;
	wire new_net_678;
	wire new_net_1853;
	wire new_net_2343;
	wire new_net_2640;
	wire new_net_2938;
	wire new_net_1403;
	wire new_net_2607;
	wire new_net_2936;
	wire new_net_2753;
	wire new_net_1986;
	wire new_net_1693;
	wire new_net_3412;
	wire new_net_1989;
	wire new_net_2359;
	wire new_net_591;
	wire new_net_609;
	wire new_net_714;
	wire new_net_852;
	wire new_net_1008;
	wire new_net_1179;
	wire new_net_1657;
	wire new_net_1727;
	wire new_net_1800;
	wire new_net_2135;
	wire new_net_2148;
	wire new_net_2455;
	wire new_net_2986;
	wire new_net_1969;
	wire _0328_;
	wire new_net_2293;
	wire new_net_2911;
	wire new_net_1609;
	wire new_net_2504;
	wire new_net_1275;
	wire _0345_;
	wire _0686_;
	wire _0560_;
	wire new_net_61;
	wire _0434_;
	wire _0728_;
	wire _0369_;
	wire _0602_;
	wire _0182_;
	wire _0014_;
	wire _0056_;
	wire new_net_807;
	wire new_net_1712;
	wire new_net_2593;
	wire new_net_2849;
	wire new_net_3269;
	wire new_net_3394;
	wire new_net_2781;
	wire new_net_2853;
	wire _0386_;
	wire new_net_607;
	wire new_net_3213;
	wire new_net_3431;
	wire new_net_949;
	wire new_net_3358;
	wire new_net_2851;
	wire _0410_;
	wire new_net_1620;
	wire new_net_1754;
	wire new_net_3280;
	wire _0695_;
	wire new_net_2249;
	wire new_net_2243;
	wire new_net_149;
	wire new_net_170;
	wire new_net_206;
	wire new_net_314;
	wire _0427_;
	wire new_net_503;
	wire new_net_698;
	wire new_net_902;
	wire new_net_1463;
	wire new_net_1277;
	wire new_net_1519;
	wire new_net_2394;
	wire new_net_2824;
	wire new_net_2392;
	wire new_net_3369;
	wire new_net_2073;
	wire _0736_;
	wire new_net_2153;
	wire new_net_2206;
	wire new_net_2114;
	wire new_net_849;
	wire new_net_1734;
	wire new_net_777;
	wire new_net_2835;
	wire new_net_1122;
	wire new_net_1432;
	wire new_net_1861;
	wire new_net_1494;
	wire new_net_2655;
	wire _0645_;
	wire _0519_;
	wire _0687_;
	wire _0561_;
	wire _0435_;
	wire _0729_;
	wire _0183_;
	wire _0225_;
	wire _0267_;
	wire _0057_;
	wire _0770_;
	wire new_net_1118;
	wire new_net_3084;
	wire new_net_3344;
	wire _0206_;
	wire new_net_1308;
	wire new_net_1366;
	wire new_net_3287;
	wire new_net_0;
	wire new_net_3130;
	wire new_net_1189;
	wire new_net_3128;
	wire _0223_;
	wire new_net_418;
	wire new_net_7;
	wire new_net_9;
	wire new_net_523;
	wire new_net_592;
	wire new_net_610;
	wire new_net_715;
	wire new_net_853;
	wire new_net_1009;
	wire new_net_1117;
	wire new_net_1919;
	wire new_net_2350;
	wire new_net_3097;
	wire new_net_2562;
	wire new_net_1983;
	wire _0264_;
	wire new_net_2485;
	wire new_net_1762;
	wire _0288_;
	wire new_net_1857;
	wire new_net_2565;
	wire _0573_;
	wire new_net_1962;
	wire new_net_2943;
	wire new_net_2798;
	wire new_net_2612;
	wire new_net_1662;
	wire _0604_;
	wire _0478_;
	wire _0772_;
	wire _0646_;
	wire _0520_;
	wire _0688_;
	wire _0562_;
	wire _0142_;
	wire _0184_;
	wire _0226_;
	wire _0590_;
	wire _0614_;
	wire new_net_649;
	wire new_net_2364;
	wire new_net_3261;
	wire _0631_;
	wire new_net_3363;
	wire new_net_3265;
	wire new_net_2192;
	wire new_net_2548;
	wire new_net_3390;
	wire _0655_;
	wire new_net_1783;
	wire new_net_2543;
	wire new_net_315;
	wire new_net_114;
	wire new_net_150;
	wire new_net_171;
	wire new_net_207;
	wire new_net_504;
	wire new_net_885;
	wire new_net_903;
	wire new_net_1091;
	wire new_net_1112;
	wire new_net_1614;
	wire new_net_1781;
	wire new_net_3312;
	wire new_net_3427;
	wire _0084_;
	wire new_net_1972;
	wire new_net_2476;
	wire new_net_2598;
	wire new_net_1648;
	wire new_net_3399;
	wire _0101_;
	wire new_net_2786;
	wire new_net_3100;
	wire new_net_58;
	wire new_net_1395;
	wire new_net_1550;
	wire new_net_1926;
	wire new_net_3365;
	wire _0125_;
	wire new_net_3385;
	wire _0437_;
	wire _0731_;
	wire _0605_;
	wire _0479_;
	wire _0773_;
	wire new_net_241;
	wire _0647_;
	wire _0521_;
	wire _0689_;
	wire _0143_;
	wire new_net_2678;
	wire new_net_1271;
	wire new_net_3072;
	wire new_net_1625;
	wire new_net_3376;
	wire new_net_2864;
	wire _0166_;
	wire new_net_2399;
	wire new_net_3374;
	wire _0451_;
	wire new_net_1565;
	wire new_net_506;
	wire new_net_3235;
	wire new_net_1826;
	wire new_net_2219;
	wire new_net_1741;
	wire new_net_2915;
	wire new_net_1368;
	wire new_net_419;
	wire new_net_10;
	wire _0468_;
	wire new_net_62;
	wire new_net_524;
	wire new_net_593;
	wire new_net_611;
	wire new_net_767;
	wire new_net_836;
	wire new_net_956;
	wire new_net_1426;
	wire _0492_;
	wire new_net_2157;
	wire new_net_1916;
	wire new_net_2840;
	wire new_net_1380;
	wire new_net_1839;
	wire new_net_3349;
	wire _0509_;
	wire new_net_1901;
	wire new_net_1641;
	wire new_net_2032;
	wire _0533_;
	wire new_net_874;
	wire new_net_2391;
	wire new_net_3135;
	wire _0564_;
	wire _0438_;
	wire _0732_;
	wire _0606_;
	wire _0480_;
	wire _0774_;
	wire _0648_;
	wire _0018_;
	wire _0060_;
	wire _0102_;
	wire new_net_2039;
	wire _0550_;
	wire new_net_2479;
	wire new_net_2677;
	wire new_net_2139;
	wire new_net_2418;
	wire new_net_1585;
	wire new_net_3407;
	wire new_net_3430;
	wire new_net_2175;
	wire new_net_765;
	wire new_net_2278;
	wire new_net_144;
	wire new_net_1959;
	wire new_net_115;
	wire new_net_151;
	wire new_net_172;
	wire new_net_505;
	wire new_net_886;
	wire new_net_904;
	wire new_net_1151;
	wire new_net_1523;
	wire new_net_1810;
	wire new_net_1817;
	wire new_net_1964;
	wire new_net_2618;
	wire new_net_2648;
	wire new_net_2767;
	wire new_net_2948;
	wire new_net_1667;
	wire new_net_2687;
	wire _0329_;
	wire new_net_583;
	wire new_net_2594;
	wire new_net_2263;
	wire _0061_;
	wire new_net_2369;
	wire _0346_;
	wire new_net_590;
	wire _0523_;
	wire _0691_;
	wire _0565_;
	wire _0439_;
	wire _0733_;
	wire _0607_;
	wire _0481_;
	wire _0370_;
	wire _0775_;
	wire new_net_242;
	wire new_net_2199;
	wire new_net_2661;
	wire new_net_2553;
	wire new_net_1455;
	wire new_net_1261;
	wire new_net_2233;
	wire new_net_3317;
	wire _0387_;
	wire new_net_2625;
	wire new_net_3181;
	wire new_net_1789;
	wire _0411_;
	wire new_net_825;
	wire new_net_1588;
	wire _0696_;
	wire new_net_1273;
	wire new_net_1331;
	wire new_net_2674;
	wire new_net_3218;
	wire new_net_63;
	wire new_net_420;
	wire new_net_525;
	wire new_net_594;
	wire new_net_612;
	wire new_net_768;
	wire new_net_837;
	wire _0428_;
	wire new_net_957;
	wire new_net_1745;
	wire new_net_1903;
	wire new_net_2250;
	wire new_net_3292;
	wire _0737_;
	wire new_net_2285;
	wire _0730_;
	wire new_net_2053;
	wire new_net_2355;
	wire new_net_2721;
	wire new_net_3416;
	wire new_net_1998;
	wire _0754_;
	wire new_net_3381;
	wire new_net_2289;
	wire new_net_2401;
	wire new_net_3298;
	wire _0482_;
	wire _0776_;
	wire _0650_;
	wire new_net_316;
	wire _0524_;
	wire _0692_;
	wire _0566_;
	wire new_net_208;
	wire _0440_;
	wire _0734_;
	wire _0778_;
	wire new_net_995;
	wire _0015_;
	wire _0771_;
	wire new_net_240;
	wire new_net_2732;
	wire new_net_3167;
	wire new_net_2920;
	wire new_net_3205;
	wire new_net_2584;
	wire new_net_3233;
	wire _0207_;
	wire _0795_;
	wire new_net_2266;
	wire new_net_1887;
	wire new_net_3087;
	wire new_net_3064;
	wire new_net_3211;
	wire _0224_;
	wire new_net_8;
	wire new_net_116;
	wire new_net_152;
	wire _0248_;
	wire new_net_173;
	wire new_net_887;
	wire new_net_905;
	wire new_net_1018;
	wire new_net_1045;
	wire new_net_1103;
	wire new_net_3142;
	wire new_net_2043;
	wire new_net_3140;
	wire _0265_;
	wire new_net_1025;
	wire new_net_413;
	wire new_net_2484;
	wire _0289_;
	wire new_net_2144;
	wire _0574_;
	wire new_net_1766;
	wire new_net_2570;
	wire _0735_;
	wire _0609_;
	wire _0483_;
	wire _0777_;
	wire new_net_243;
	wire _0651_;
	wire _0306_;
	wire _0525_;
	wire _0693_;
	wire _0567_;
	wire _0591_;
	wire new_net_2017;
	wire new_net_1418;
	wire new_net_1935;
	wire new_net_2456;
	wire _0615_;
	wire new_net_2955;
	wire new_net_2772;
	wire _0608_;
	wire new_net_3340;
	wire new_net_2622;
	wire new_net_3315;
	wire _0632_;
	wire new_net_2300;
	wire new_net_2874;
	wire _0656_;
	wire new_net_64;
	wire new_net_421;
	wire new_net_526;
	wire new_net_595;
	wire new_net_769;
	wire new_net_958;
	wire new_net_1239;
	wire new_net_1508;
	wire _0649_;
	wire new_net_665;
	wire new_net_2900;
	wire new_net_2167;
	wire _0673_;
	wire new_net_2666;
	wire new_net_1391;
	wire new_net_2308;
	wire new_net_3002;
	wire new_net_2235;
	wire new_net_2518;
	wire new_net_1467;
	wire _0690_;
	wire new_net_1507;
	wire new_net_2245;
	wire _0126_;
	wire new_net_1267;
	wire new_net_2239;
	wire new_net_1534;
	wire new_net_3186;
	wire new_net_1658;
	wire new_net_3223;
	wire new_net_1557;
	wire new_net_3107;
	wire _0167_;
	wire new_net_1796;
	wire new_net_2254;
	wire new_net_1422;
	wire new_net_1881;
	wire new_net_3201;
	wire new_net_1292;
	wire new_net_2726;
	wire new_net_515;
	wire new_net_1674;
	wire new_net_2003;
	wire new_net_3060;
	wire new_net_3386;
	wire new_net_317;
	wire new_net_209;
	wire new_net_278;
	wire new_net_368;
	wire new_net_977;
	wire new_net_1086;
	wire new_net_1224;
	wire new_net_1325;
	wire new_net_1367;
	wire new_net_1409;
	wire new_net_2133;
	wire new_net_3303;
	wire new_net_2810;
	wire new_net_1447;
	wire new_net_2630;
	wire new_net_2737;
	wire new_net_3172;
	wire new_net_1813;
	wire new_net_3094;
	wire new_net_2589;
	wire new_net_2697;
	wire new_net_1851;
	wire new_net_2395;
	wire new_net_2448;
	wire new_net_1323;
	wire new_net_1542;
	wire new_net_1816;
	wire new_net_2344;
	wire new_net_11;
	wire new_net_117;
	wire new_net_174;
	wire new_net_261;
	wire new_net_438;
	wire new_net_735;
	wire new_net_906;
	wire new_net_1046;
	wire new_net_1120;
	wire new_net_1143;
	wire new_net_3147;
	wire new_net_2712;
	wire new_net_3290;
	wire new_net_2490;
	wire new_net_2682;
	wire new_net_1768;
	wire new_net_3153;
	wire new_net_3336;
	wire new_net_3258;
	wire new_net_28;
	wire new_net_244;
	wire new_net_352;
	wire new_net_82;
	wire new_net_544;
	wire new_net_613;
	wire new_net_667;
	wire new_net_718;
	wire new_net_1152;
	wire new_net_1168;
	wire new_net_1296;
	wire new_net_1354;
	wire new_net_1694;
	wire _0330_;
	wire new_net_1199;
	wire _0062_;
	wire new_net_2960;
	wire new_net_2328;
	wire _0347_;
	wire new_net_1451;
	wire new_net_1971;
	wire _0371_;
	wire new_net_2881;
	wire new_net_739;
	wire new_net_335;
	wire new_net_386;
	wire new_net_422;
	wire new_net_455;
	wire new_net_560;
	wire new_net_785;
	wire new_net_959;
	wire new_net_1166;
	wire new_net_1784;
	wire new_net_1910;
	wire new_net_1973;
	wire new_net_2376;
	wire _0388_;
	wire new_net_608;
	wire new_net_1385;
	wire new_net_1846;
	wire new_net_2098;
	wire _0412_;
	wire new_net_2523;
	wire new_net_3069;
	wire new_net_3011;
	wire new_net_369;
	wire new_net_279;
	wire new_net_471;
	wire new_net_1180;
	wire new_net_1294;
	wire new_net_1336;
	wire new_net_1170;
	wire new_net_1357;
	wire new_net_1399;
	wire _0738_;
	wire new_net_2758;
	wire new_net_3225;
	wire new_net_850;
	wire new_net_778;
	wire new_net_1562;
	wire new_net_3112;
	wire new_net_1529;
	wire new_net_2839;
	wire new_net_2991;
	wire _0779_;
	wire new_net_1067;
	wire new_net_3419;
	wire new_net_1564;
	wire new_net_930;
	wire _0016_;
	wire new_net_175;
	wire new_net_262;
	wire new_net_631;
	wire new_net_736;
	wire new_net_856;
	wire new_net_907;
	wire new_net_925;
	wire new_net_1047;
	wire new_net_1082;
	wire _0208_;
	wire new_net_2010;
	wire new_net_2160;
	wire new_net_2509;
	wire new_net_2008;
	wire new_net_2731;
	wire new_net_1577;
	wire new_net_2636;
	wire new_net_2927;
	wire new_net_2744;
	wire _0249_;
	wire new_net_1123;
	wire new_net_2742;
	wire new_net_2791;
	wire new_net_1644;
	wire new_net_2670;
	wire new_net_65;
	wire new_net_353;
	wire new_net_245;
	wire new_net_527;
	wire new_net_545;
	wire new_net_614;
	wire new_net_668;
	wire new_net_719;
	wire new_net_770;
	wire _0266_;
	wire new_net_2273;
	wire _0290_;
	wire new_net_1872;
	wire new_net_3332;
	wire new_net_2902;
	wire new_net_2645;
	wire new_net_1414;
	wire new_net_2454;
	wire new_net_2683;
	wire _0307_;
	wire new_net_2495;
	wire new_net_2717;
	wire new_net_2320;
	wire _0592_;
	wire new_net_2493;
	wire new_net_210;
	wire new_net_318;
	wire new_net_336;
	wire new_net_561;
	wire new_net_786;
	wire new_net_650;
	wire new_net_960;
	wire new_net_1068;
	wire new_net_1069;
	wire new_net_1073;
	wire new_net_1636;
	wire new_net_2119;
	wire new_net_3158;
	wire new_net_3414;
	wire new_net_1701;
	wire new_net_2259;
	wire _0633_;
	wire new_net_1774;
	wire new_net_2163;
	wire new_net_2701;
	wire new_net_118;
	wire new_net_280;
	wire new_net_439;
	wire new_net_472;
	wire new_net_1079;
	wire _0674_;
	wire new_net_1092;
	wire new_net_1146;
	wire new_net_1169;
	wire new_net_1326;
	wire new_net_1546;
	wire new_net_2970;
	wire new_net_2886;
	wire new_net_1263;
	wire new_net_2383;
	wire _0103_;
	wire new_net_1589;
	wire new_net_1722;
	wire new_net_2381;
	wire new_net_2451;
	wire new_net_2105;
	wire new_net_3007;
	wire new_net_2211;
	wire new_net_2103;
	wire new_net_2283;
	wire new_net_2530;
	wire new_net_12;
	wire new_net_29;
	wire new_net_83;
	wire new_net_176;
	wire new_net_263;
	wire _0144_;
	wire new_net_632;
	wire new_net_637;
	wire new_net_737;
	wire new_net_857;
	wire new_net_1479;
	wire new_net_2528;
	wire new_net_2657;
	wire new_net_3018;
	wire _0168_;
	wire new_net_1288;
	wire new_net_2763;
	wire new_net_507;
	wire new_net_1670;
	wire new_net_1803;
	wire new_net_1827;
	wire new_net_3230;
	wire _0185_;
	wire new_net_1801;
	wire new_net_3119;
	wire new_net_1807;
	wire new_net_3117;
	wire new_net_387;
	wire new_net_66;
	wire new_net_354;
	wire new_net_423;
	wire new_net_456;
	wire new_net_528;
	wire new_net_546;
	wire new_net_615;
	wire new_net_720;
	wire new_net_771;
	wire new_net_1443;
	wire new_net_2996;
	wire new_net_3424;
	wire new_net_1160;
	wire new_net_2362;
	wire new_net_1319;
	wire new_net_2413;
	wire new_net_1377;
	wire new_net_2136;
	wire new_net_875;
	wire new_net_2514;
	wire new_net_1582;
	wire new_net_1897;
	wire new_net_2603;
	wire new_net_211;
	wire _0552_;
	wire new_net_319;
	wire new_net_337;
	wire new_net_370;
	wire new_net_961;
	wire new_net_979;
	wire new_net_1606;
	wire new_net_1618;
	wire new_net_1661;
	wire new_net_2419;
	wire new_net_2749;
	wire new_net_1931;
	wire new_net_3253;
	wire new_net_766;
	wire new_net_1629;
	wire new_net_145;
	wire new_net_2397;
	wire new_net_1350;
	wire new_net_2982;
	wire new_net_1408;
	wire new_net_1877;
	wire new_net_2183;
	wire new_net_1632;
	wire new_net_1965;
	wire new_net_2907;
	wire new_net_119;
	wire new_net_281;
	wire new_net_440;
	wire new_net_473;
	wire new_net_1130;
	wire new_net_1137;
	wire new_net_1228;
	wire new_net_1295;
	wire new_net_1337;
	wire new_net_1358;
	wire new_net_1605;
	wire new_net_1994;
	wire new_net_2181;
	wire new_net_2435;
	wire new_net_2500;
	wire _0331_;
	wire new_net_584;
	wire new_net_722;
	wire new_net_1603;
	wire new_net_2124;
	wire _0063_;
	wire new_net_3163;
	wire new_net_2845;
	wire _0348_;
	wire new_net_1706;
	wire new_net_2334;
	wire _0372_;
	wire new_net_1381;
	wire new_net_1844;
	wire new_net_30;
	wire new_net_84;
	wire new_net_177;
	wire new_net_246;
	wire new_net_264;
	wire new_net_669;
	wire new_net_738;
	wire new_net_858;
	wire new_net_927;
	wire new_net_1116;
	wire new_net_1750;
	wire new_net_3276;
	wire new_net_2203;
	wire _0389_;
	wire _0413_;
	wire new_net_826;
	wire new_net_1953;
	wire new_net_2893;
	wire _0698_;
	wire new_net_685;
	wire new_net_2820;
	wire new_net_2975;
	wire new_net_2388;
	wire new_net_2069;
	wire new_net_2149;
	wire new_net_833;
	wire new_net_424;
	wire new_net_13;
	wire _0715_;
	wire new_net_388;
	wire new_net_457;
	wire new_net_529;
	wire new_net_562;
	wire new_net_616;
	wire new_net_787;
	wire new_net_842;
	wire new_net_2110;
	wire _0739_;
	wire new_net_2831;
	wire new_net_2535;
	wire new_net_913;
	wire new_net_699;
	wire new_net_1282;
	wire new_net_2829;
	wire new_net_2404;
	wire new_net_3023;
	wire _0000_;
	wire new_net_1172;
	wire new_net_2402;
	wire _0780_;
	wire new_net_996;
	wire new_net_1832;
	wire new_net_212;
	wire new_net_371;
	wire _0017_;
	wire new_net_962;
	wire new_net_980;
	wire new_net_1219;
	wire new_net_1251;
	wire new_net_1437;
	wire new_net_1596;
	wire new_net_1624;
	wire new_net_1890;
	wire new_net_3124;
	wire _0209_;
	wire new_net_1888;
	wire new_net_2408;
	wire new_net_3031;
	wire new_net_1012;
	wire new_net_2036;
	wire new_net_2449;
	wire new_net_2439;
	wire new_net_1313;
	wire new_net_3035;
	wire new_net_2558;
	wire _0250_;
	wire new_net_1019;
	wire new_net_2018;
	wire new_net_1758;
	wire new_net_3322;
	wire new_net_282;
	wire new_net_474;
	wire new_net_633;
	wire new_net_909;
	wire new_net_1327;
	wire new_net_1369;
	wire new_net_1411;
	wire new_net_1453;
	wire new_net_1566;
	wire new_net_1578;
	wire new_net_1854;
	wire new_net_3249;
	wire new_net_1026;
	wire new_net_2488;
	wire new_net_2939;
	wire new_net_1410;
	wire new_net_414;
	wire new_net_2608;
	wire _0291_;
	wire new_net_2754;
	wire _0576_;
	wire new_net_3413;
	wire _0308_;
	wire new_net_2360;
	wire new_net_3166;
	wire _0593_;
	wire new_net_265;
	wire new_net_67;
	wire new_net_85;
	wire new_net_178;
	wire new_net_355;
	wire new_net_247;
	wire new_net_547;
	wire new_net_670;
	wire _0617_;
	wire new_net_721;
	wire new_net_1241;
	wire new_net_2987;
	wire new_net_2188;
	wire new_net_2294;
	wire new_net_2912;
	wire new_net_2540;
	wire new_net_3308;
	wire _0634_;
	wire new_net_2505;
	wire new_net_1941;
	wire new_net_2776;
	wire _0658_;
	wire new_net_666;
	wire new_net_1713;
	wire new_net_320;
	wire new_net_338;
	wire new_net_563;
	wire new_net_617;
	wire new_net_788;
	wire new_net_1060;
	wire new_net_1465;
	wire new_net_1477;
	wire _0675_;
	wire new_net_1490;
	wire new_net_2093;
	wire new_net_2782;
	wire new_net_2850;
	wire new_net_1922;
	wire new_net_3395;
	wire new_net_2854;
	wire new_net_1847;
	wire new_net_2947;
	wire new_net_3041;
	wire new_net_3359;
	wire _0104_;
	wire new_net_1755;
	wire new_net_3281;
	wire new_net_2856;
	wire new_net_2424;
	wire new_net_2898;
	wire new_net_1284;
	wire new_net_120;
	wire new_net_213;
	wire new_net_441;
	wire new_net_963;
	wire new_net_1145;
	wire new_net_1342;
	wire new_net_1520;
	wire new_net_1558;
	wire _0145_;
	wire new_net_1597;
	wire new_net_2074;
	wire new_net_2393;
	wire new_net_2825;
	wire new_net_3232;
	wire new_net_2115;
	wire new_net_3081;
	wire new_net_2836;
	wire _0186_;
	wire new_net_1495;
	wire new_net_2656;
	wire _0471_;
	wire new_net_516;
	wire new_net_5;
	wire new_net_31;
	wire new_net_283;
	wire new_net_475;
	wire new_net_634;
	wire new_net_859;
	wire new_net_910;
	wire new_net_928;
	wire new_net_1074;
	wire new_net_1185;
	wire new_net_1315;
	wire new_net_1373;
	wire new_net_2440;
	wire new_net_3131;
	wire _0512_;
	wire new_net_3129;
	wire _0536_;
	wire new_net_248;
	wire new_net_389;
	wire new_net_14;
	wire new_net_68;
	wire _0553_;
	wire new_net_86;
	wire new_net_179;
	wire new_net_266;
	wire new_net_356;
	wire new_net_425;
	wire new_net_2274;
	wire new_net_1984;
	wire new_net_2563;
	wire new_net_2579;
	wire new_net_1057;
	wire new_net_1346;
	wire new_net_2567;
	wire new_net_1404;
	wire new_net_1963;
	wire new_net_1987;
	wire new_net_2944;
	wire new_net_1663;
	wire new_net_1990;
	wire new_net_2613;
	wire new_net_2691;
	wire new_net_1070;
	wire new_net_321;
	wire new_net_339;
	wire new_net_564;
	wire new_net_618;
	wire new_net_981;
	wire new_net_1187;
	wire new_net_1748;
	wire new_net_2177;
	wire new_net_2026;
	wire new_net_1511;
	wire new_net_2365;
	wire new_net_2917;
	wire _0332_;
	wire new_net_1202;
	wire new_net_3262;
	wire new_net_2659;
	wire new_net_2195;
	wire new_net_2337;
	wire new_net_2164;
	wire new_net_3266;
	wire new_net_2193;
	wire new_net_2549;
	wire _0349_;
	wire new_net_1617;
	wire new_net_2230;
	wire new_net_3313;
	wire new_net_1782;
	wire new_net_121;
	wire _0373_;
	wire new_net_442;
	wire new_net_602;
	wire new_net_740;
	wire new_net_194;
	wire new_net_964;
	wire new_net_1095;
	wire new_net_1129;
	wire new_net_1225;
	wire new_net_1615;
	wire new_net_2950;
	wire new_net_3177;
	wire new_net_2968;
	wire new_net_2338;
	wire new_net_2472;
	wire _0390_;
	wire new_net_1718;
	wire new_net_2599;
	wire new_net_3214;
	wire _0414_;
	wire new_net_1460;
	wire new_net_2787;
	wire new_net_1927;
	wire _0699_;
	wire new_net_3101;
	wire new_net_1226;
	wire new_net_2349;
	wire new_net_3366;
	wire new_net_2212;
	wire new_net_3288;
	wire new_net_3364;
	wire new_net_2208;
	wire new_net_284;
	wire new_net_32;
	wire new_net_476;
	wire new_net_635;
	wire new_net_671;
	wire _0716_;
	wire new_net_860;
	wire new_net_911;
	wire new_net_929;
	wire new_net_1093;
	wire new_net_1278;
	wire new_net_3073;
	wire new_net_772;
	wire new_net_3240;
	wire _0740_;
	wire new_net_3377;
	wire new_net_3375;
	wire new_net_3236;
	wire _0757_;
	wire new_net_2220;
	wire new_net_1433;
	wire new_net_1742;
	wire new_net_2580;
	wire new_net_2916;
	wire _0781_;
	wire new_net_357;
	wire new_net_426;
	wire new_net_15;
	wire new_net_69;
	wire new_net_87;
	wire new_net_180;
	wire new_net_249;
	wire new_net_390;
	wire new_net_459;
	wire new_net_531;
	wire new_net_1912;
	wire new_net_2841;
	wire _0210_;
	wire new_net_1309;
	wire new_net_3350;
	wire new_net_3244;
	wire new_net_1976;
	wire _0227_;
	wire new_net_3136;
	wire _0251_;
	wire new_net_322;
	wire new_net_214;
	wire new_net_373;
	wire new_net_565;
	wire new_net_619;
	wire new_net_982;
	wire new_net_1547;
	wire new_net_1559;
	wire new_net_1866;
	wire new_net_2186;
	wire new_net_2140;
	wire new_net_2480;
	wire new_net_1586;
	wire new_net_3300;
	wire _0268_;
	wire _0292_;
	wire new_net_2279;
	wire _0577_;
	wire _0309_;
	wire new_net_1043;
	wire new_net_2951;
	wire new_net_2768;
	wire new_net_443;
	wire _0594_;
	wire new_net_965;
	wire new_net_1063;
	wire new_net_1072;
	wire new_net_1102;
	wire new_net_1218;
	wire new_net_1512;
	wire new_net_1598;
	wire new_net_1902;
	wire new_net_1908;
	wire _0618_;
	wire new_net_651;
	wire new_net_1668;
	wire new_net_2688;
	wire new_net_2325;
	wire new_net_2870;
	wire new_net_1217;
	wire new_net_2962;
	wire new_net_2329;
	wire new_net_2468;
	wire _0635_;
	wire new_net_658;
	wire new_net_3168;
	wire _0659_;
	wire new_net_2662;
	wire new_net_2200;
	wire new_net_33;
	wire new_net_267;
	wire new_net_285;
	wire new_net_477;
	wire new_net_549;
	wire new_net_636;
	wire new_net_672;
	wire new_net_723;
	wire new_net_861;
	wire new_net_912;
	wire new_net_1462;
	wire _0676_;
	wire new_net_1503;
	wire new_net_2554;
	wire new_net_1975;
	wire new_net_2234;
	wire new_net_548;
	wire new_net_3318;
	wire new_net_3182;
	wire _0105_;
	wire new_net_1790;
	wire new_net_1338;
	wire new_net_60;
	wire new_net_1396;
	wire new_net_2675;
	wire new_net_1654;
	wire new_net_3219;
	wire new_net_16;
	wire new_net_88;
	wire _0153_;
	wire new_net_340;
	wire new_net_532;
	wire new_net_742;
	wire new_net_790;
	wire new_net_1190;
	wire new_net_1749;
	wire new_net_638;
	wire new_net_2478;
	wire _0146_;
	wire new_net_1272;
	wire new_net_2244;
	wire new_net_2319;
	wire new_net_3293;
	wire new_net_2286;
	wire new_net_2079;
	wire _0455_;
	wire new_net_2054;
	wire new_net_1921;
	wire new_net_2154;
	wire new_net_2356;
	wire new_net_508;
	wire new_net_1999;
	wire new_net_2722;
	wire new_net_3417;
	wire new_net_3382;
	wire new_net_3049;
	wire _0187_;
	wire new_net_1525;
	wire new_net_1203;
	wire new_net_3299;
	wire _0472_;
	wire new_net_1427;
	wire new_net_1571;
	wire new_net_215;
	wire new_net_374;
	wire new_net_6;
	wire new_net_323;
	wire new_net_122;
	wire new_net_566;
	wire new_net_983;
	wire _0496_;
	wire new_net_1089;
	wire new_net_1191;
	wire new_net_2229;
	wire new_net_2733;
	wire new_net_2921;
	wire new_net_3090;
	wire new_net_2585;
	wire new_net_2816;
	wire new_net_2267;
	wire new_net_3151;
	wire new_net_3206;
	wire new_net_3088;
	wire _0513_;
	wire new_net_111;
	wire new_net_3212;
	wire _0537_;
	wire new_net_1198;
	wire new_net_1680;
	wire new_net_2272;
	wire new_net_2417;
	wire new_net_444;
	wire new_net_966;
	wire new_net_1939;
	wire new_net_2064;
	wire new_net_1979;
	wire new_net_1400;
	wire new_net_2724;
	wire _0554_;
	wire new_net_2708;
	wire new_net_2044;
	wire new_net_3143;
	wire new_net_3141;
	wire new_net_2486;
	wire new_net_3077;
	wire new_net_2145;
	wire new_net_146;
	wire new_net_1049;
	wire new_net_1690;
	wire new_net_2571;
	wire new_net_3152;
	wire new_net_391;
	wire new_net_70;
	wire new_net_286;
	wire new_net_358;
	wire new_net_427;
	wire new_net_34;
	wire new_net_181;
	wire new_net_250;
	wire new_net_268;
	wire new_net_460;
	wire new_net_578;
	wire new_net_2457;
	wire new_net_2956;
	wire new_net_2773;
	wire _0333_;
	wire new_net_2623;
	wire new_net_1186;
	wire _0350_;
	wire new_net_2372;
	wire new_net_2875;
	wire new_net_1948;
	wire new_net_2061;
	wire new_net_17;
	wire new_net_341;
	wire new_net_620;
	wire _0374_;
	wire new_net_743;
	wire new_net_791;
	wire new_net_1560;
	wire new_net_2042;
	wire new_net_2094;
	wire new_net_2187;
	wire new_net_1456;
	wire new_net_2309;
	wire new_net_2204;
	wire _0391_;
	wire new_net_815;
	wire new_net_2236;
	wire new_net_2209;
	wire new_net_2519;
	wire new_net_3003;
	wire _0415_;
	wire new_net_827;
	wire _0700_;
	wire new_net_686;
	wire new_net_1274;
	wire new_net_2246;
	wire new_net_2240;
	wire new_net_3189;
	wire new_net_123;
	wire new_net_216;
	wire new_net_567;
	wire _0432_;
	wire new_net_834;
	wire new_net_984;
	wire new_net_1107;
	wire new_net_1121;
	wire _0717_;
	wire new_net_1214;
	wire new_net_3104;
	wire new_net_1659;
	wire new_net_843;
	wire new_net_3224;
	wire new_net_2214;
	wire new_net_3108;
	wire _0741_;
	wire new_net_228;
	wire new_net_914;
	wire new_net_700;
	wire _0758_;
	wire new_net_235;
	wire new_net_3202;
	wire new_net_2434;
	wire _0782_;
	wire new_net_862;
	wire new_net_931;
	wire new_net_967;
	wire new_net_1126;
	wire new_net_1144;
	wire new_net_1305;
	wire new_net_1363;
	wire new_net_1675;
	wire _0019_;
	wire new_net_716;
	wire new_net_2004;
	wire new_net_3054;
	wire new_net_3061;
	wire new_net_3304;
	wire new_net_3387;
	wire new_net_2134;
	wire new_net_2409;
	wire new_net_1;
	wire new_net_2631;
	wire new_net_3173;
	wire new_net_3400;
	wire new_net_2738;
	wire new_net_1814;
	wire new_net_673;
	wire new_net_1642;
	wire _0228_;
	wire new_net_2698;
	wire _0252_;
	wire new_net_35;
	wire new_net_182;
	wire new_net_251;
	wire new_net_392;
	wire new_net_71;
	wire new_net_287;
	wire new_net_359;
	wire new_net_428;
	wire new_net_89;
	wire new_net_461;
	wire new_net_1543;
	wire new_net_2345;
	wire new_net_2638;
	wire _0269_;
	wire new_net_1027;
	wire new_net_1127;
	wire new_net_1957;
	wire new_net_415;
	wire new_net_3326;
	wire new_net_3148;
	wire _0293_;
	wire new_net_2713;
	wire _0578_;
	wire new_net_2614;
	wire new_net_1991;
	wire _0310_;
	wire new_net_18;
	wire new_net_324;
	wire new_net_375;
	wire new_net_621;
	wire _0595_;
	wire new_net_744;
	wire new_net_792;
	wire new_net_1231;
	wire new_net_1569;
	wire new_net_1581;
	wire new_net_1697;
	wire new_net_1419;
	wire new_net_3259;
	wire new_net_1695;
	wire _0619_;
	wire new_net_1777;
	wire new_net_2576;
	wire _0636_;
	wire new_net_3050;
	wire _0660_;
	wire new_net_124;
	wire new_net_445;
	wire new_net_568;
	wire new_net_985;
	wire new_net_1062;
	wire new_net_1155;
	wire new_net_1487;
	wire new_net_1977;
	wire new_net_2080;
	wire new_net_2725;
	wire new_net_2882;
	wire _0677_;
	wire new_net_2377;
	wire new_net_52;
	wire new_net_1392;
	wire new_net_1548;
	wire _0113_;
	wire new_net_2099;
	wire new_net_1475;
	wire new_net_1268;
	wire new_net_2524;
	wire new_net_269;
	wire new_net_725;
	wire new_net_863;
	wire new_net_932;
	wire new_net_1066;
	wire new_net_491;
	wire new_net_1149;
	wire new_net_1473;
	wire new_net_1610;
	wire new_net_1665;
	wire new_net_2207;
	wire new_net_2425;
	wire new_net_3012;
	wire new_net_3194;
	wire _0147_;
	wire new_net_2759;
	wire new_net_2216;
	wire new_net_3226;
	wire new_net_3198;
	wire new_net_2953;
	wire _0456_;
	wire new_net_1423;
	wire new_net_1563;
	wire new_net_3113;
	wire _0188_;
	wire new_net_1293;
	wire new_net_2992;
	wire new_net_72;
	wire new_net_288;
	wire new_net_429;
	wire new_net_90;
	wire new_net_36;
	wire new_net_342;
	wire _0473_;
	wire new_net_252;
	wire new_net_462;
	wire new_net_480;
	wire _0497_;
	wire new_net_517;
	wire new_net_1946;
	wire new_net_2441;
	wire new_net_2807;
	wire new_net_2011;
	wire new_net_2510;
	wire new_net_2009;
	wire _0514_;
	wire new_net_1448;
	wire new_net_1893;
	wire new_net_1970;
	wire new_net_2813;
	wire _0538_;
	wire new_net_2637;
	wire new_net_2745;
	wire new_net_2928;
	wire new_net_217;
	wire new_net_325;
	wire new_net_376;
	wire new_net_622;
	wire new_net_745;
	wire new_net_793;
	wire new_net_1324;
	wire new_net_1645;
	wire new_net_2070;
	wire new_net_2511;
	wire _0555_;
	wire new_net_2671;
	wire new_net_2792;
	wire new_net_1873;
	wire new_net_2903;
	wire new_net_2646;
	wire new_net_446;
	wire new_net_569;
	wire new_net_968;
	wire new_net_986;
	wire new_net_1138;
	wire new_net_1240;
	wire new_net_1917;
	wire new_net_2122;
	wire new_net_1599;
	wire new_net_2178;
	wire new_net_2496;
	wire new_net_2867;
	wire new_net_1297;
	wire new_net_2120;
	wire new_net_1355;
	wire new_net_3159;
	wire _0334_;
	wire new_net_1702;
	wire new_net_2260;
	wire new_net_2330;
	wire new_net_803;
	wire new_net_1840;
	wire _0351_;
	wire new_net_1452;
	wire new_net_183;
	wire new_net_270;
	wire new_net_360;
	wire new_net_393;
	wire new_net_552;
	wire new_net_639;
	wire _0375_;
	wire new_net_603;
	wire new_net_726;
	wire new_net_741;
	wire new_net_864;
	wire new_net_2702;
	wire new_net_2897;
	wire new_net_1328;
	wire new_net_2971;
	wire _0392_;
	wire new_net_1386;
	wire new_net_2384;
	wire new_net_2887;
	wire _0416_;
	wire new_net_1723;
	wire new_net_2311;
	wire new_net_2056;
	wire new_net_2106;
	wire new_net_37;
	wire new_net_253;
	wire new_net_343;
	wire new_net_430;
	wire new_net_19;
	wire new_net_463;
	wire new_net_481;
	wire new_net_535;
	wire new_net_676;
	wire new_net_1221;
	wire new_net_2531;
	wire new_net_2676;
	wire new_net_2529;
	wire new_net_3019;
	wire new_net_773;
	wire new_net_3046;
	wire new_net_1359;
	wire new_net_2155;
	wire new_net_1804;
	wire new_net_2764;
	wire new_net_1828;
	wire new_net_3231;
	wire new_net_1524;
	wire new_net_1802;
	wire new_net_2083;
	wire new_net_125;
	wire new_net_218;
	wire new_net_326;
	wire new_net_377;
	wire new_net_623;
	wire new_net_794;
	wire new_net_1113;
	wire new_net_1159;
	wire new_net_1243;
	wire new_net_2443;
	wire _0020_;
	wire new_net_1535;
	wire new_net_2437;
	wire new_net_2667;
	wire new_net_2997;
	wire new_net_1003;
	wire new_net_2414;
	wire _0229_;
	wire new_net_1010;
	wire new_net_2341;
	wire new_net_2040;
	wire new_net_2515;
	wire new_net_570;
	wire new_net_933;
	wire new_net_969;
	wire new_net_987;
	wire new_net_1055;
	wire new_net_1134;
	wire new_net_1222;
	wire new_net_1238;
	wire new_net_1469;
	wire new_net_1481;
	wire new_net_1898;
	wire new_net_2415;
	wire new_net_2604;
	wire new_net_2933;
	wire new_net_2750;
	wire new_net_3098;
	wire new_net_2420;
	wire new_net_478;
	wire _0270_;
	wire new_net_1932;
	wire new_net_3409;
	wire _0294_;
	wire new_net_3254;
	wire new_net_3256;
	wire new_net_1415;
	wire new_net_2983;
	wire new_net_361;
	wire new_net_73;
	wire new_net_91;
	wire new_net_184;
	wire new_net_271;
	wire new_net_289;
	wire new_net_394;
	wire _0311_;
	wire new_net_553;
	wire new_net_640;
	wire new_net_1044;
	wire new_net_1878;
	wire new_net_1966;
	wire new_net_2184;
	wire new_net_2290;
	wire new_net_2908;
	wire new_net_1995;
	wire new_net_2501;
	wire new_net_3187;
	wire new_net_1604;
	wire new_net_2125;
	wire new_net_659;
	wire new_net_1640;
	wire new_net_1709;
	wire new_net_2590;
	wire new_net_2846;
	wire new_net_3164;
	wire new_net_1707;
	wire new_net_1500;
	wire new_net_3391;
	wire new_net_20;
	wire new_net_38;
	wire new_net_254;
	wire new_net_344;
	wire new_net_464;
	wire new_net_482;
	wire new_net_677;
	wire new_net_746;
	wire new_net_1174;
	wire new_net_1237;
	wire new_net_1388;
	wire new_net_2310;
	wire new_net_2303;
	wire new_net_2335;
	wire new_net_3355;
	wire new_net_1751;
	wire new_net_3059;
	wire new_net_3277;
	wire new_net_1264;
	wire new_net_2894;
	wire new_net_2821;
	wire new_net_2976;
	wire new_net_2389;
	wire new_net_126;
	wire new_net_219;
	wire new_net_447;
	wire new_net_795;
	wire new_net_2123;
	wire new_net_2150;
	wire new_net_2429;
	wire new_net_2436;
	wire _0155_;
	wire new_net_2444;
	wire new_net_2111;
	wire new_net_2832;
	wire new_net_1289;
	wire new_net_2536;
	wire new_net_2830;
	wire new_net_2460;
	wire new_net_1485;
	wire new_net_3024;
	wire new_net_509;
	wire new_net_2405;
	wire new_net_3341;
	wire new_net_2669;
	wire _0189_;
	wire new_net_2403;
	wire new_net_571;
	wire new_net_865;
	wire new_net_934;
	wire new_net_970;
	wire new_net_988;
	wire new_net_1128;
	wire new_net_1514;
	wire new_net_1752;
	wire new_net_1904;
	wire new_net_1993;
	wire new_net_2027;
	wire new_net_1444;
	wire new_net_1537;
	wire new_net_2812;
	wire new_net_3125;
	wire new_net_1889;
	wire new_net_112;
	wire new_net_3032;
	wire new_net_2037;
	wire new_net_1320;
	wire new_net_3036;
	wire new_net_2559;
	wire new_net_74;
	wire new_net_92;
	wire new_net_290;
	wire new_net_395;
	wire new_net_431;
	wire new_net_536;
	wire new_net_641;
	wire new_net_917;
	wire new_net_1088;
	wire new_net_1125;
	wire new_net_1759;
	wire new_net_1980;
	wire new_net_3323;
	wire new_net_2639;
	wire new_net_3250;
	wire new_net_761;
	wire new_net_3248;
	wire new_net_1956;
	wire new_net_2641;
	wire new_net_2940;
	wire new_net_2979;
	wire new_net_2609;
	wire new_net_2022;
	wire new_net_900;
	wire new_net_1351;
	wire new_net_39;
	wire new_net_327;
	wire new_net_21;
	wire new_net_378;
	wire _0033_;
	wire new_net_624;
	wire new_net_747;
	wire new_net_1051;
	wire new_net_1300;
	wire new_net_579;
	wire new_net_2321;
	wire new_net_2361;
	wire new_net_3190;
	wire new_net_2988;
	wire new_net_2161;
	wire new_net_2189;
	wire _0335_;
	wire new_net_2295;
	wire new_net_2913;
	wire new_net_3309;
	wire new_net_1153;
	wire new_net_1611;
	wire new_net_1942;
	wire new_net_2777;
	wire _0352_;
	wire new_net_127;
	wire new_net_220;
	wire new_net_448;
	wire new_net_1230;
	wire new_net_1248;
	wire new_net_1488;
	wire new_net_1493;
	wire new_net_1600;
	wire new_net_1612;
	wire _0376_;
	wire new_net_1382;
	wire new_net_1714;
	wire new_net_2595;
	wire new_net_2304;
	wire new_net_3271;
	wire new_net_3396;
	wire new_net_2783;
	wire new_net_2855;
	wire _0393_;
	wire new_net_816;
	wire new_net_1848;
	wire new_net_3067;
	wire new_net_3360;
	wire _0417_;
	wire new_net_828;
	wire new_net_1756;
	wire new_net_3282;
	wire new_net_687;
	wire new_net_2857;
	wire new_net_185;
	wire new_net_272;
	wire new_net_362;
	wire new_net_554;
	wire new_net_572;
	wire new_net_728;
	wire new_net_779;
	wire new_net_866;
	wire new_net_1551;
	wire new_net_835;
	wire new_net_1593;
	wire new_net_2396;
	wire new_net_2077;
	wire new_net_2899;
	wire _0719_;
	wire new_net_694;
	wire new_net_3053;
	wire new_net_3371;
	wire new_net_844;
	wire new_net_1732;
	wire new_net_2075;
	wire new_net_2215;
	wire new_net_1736;
	wire _0760_;
	wire new_net_2837;
	wire new_net_93;
	wire new_net_255;
	wire new_net_291;
	wire new_net_345;
	wire new_net_396;
	wire _0784_;
	wire new_net_432;
	wire new_net_465;
	wire new_net_483;
	wire new_net_537;
	wire new_net_922;
	wire new_net_1496;
	wire new_net_3346;
	wire _0021_;
	wire new_net_717;
	wire new_net_2223;
	wire new_net_1438;
	wire new_net_2410;
	wire new_net_1974;
	wire new_net_2664;
	wire new_net_1676;
	wire new_net_3243;
	wire new_net_3065;
	wire new_net_3132;
	wire new_net_1156;
	wire new_net_1960;
	wire new_net_674;
	wire _0230_;
	wire new_net_1314;
	wire new_net_22;
	wire new_net_379;
	wire new_net_40;
	wire new_net_328;
	wire new_net_625;
	wire new_net_796;
	wire new_net_1162;
	wire new_net_1332;
	wire new_net_1374;
	wire new_net_1416;
	wire new_net_2019;
	wire new_net_3404;
	wire new_net_2275;
	wire new_net_1985;
	wire _0271_;
	wire new_net_1028;
	wire new_net_1594;
	wire new_net_1630;
	wire new_net_2615;
	wire new_net_2945;
	wire new_net_128;
	wire new_net_221;
	wire new_net_449;
	wire new_net_935;
	wire new_net_971;
	wire _0312_;
	wire new_net_989;
	wire new_net_1254;
	wire new_net_1515;
	wire new_net_1649;
	wire new_net_1664;
	wire new_net_1936;
	wire new_net_2684;
	wire new_net_879;
	wire new_net_2366;
	wire new_net_2196;
	wire _0638_;
	wire new_net_2999;
	wire new_net_3267;
	wire new_net_2194;
	wire new_net_2550;
	wire new_net_273;
	wire new_net_75;
	wire new_net_363;
	wire new_net_186;
	wire new_net_555;
	wire new_net_573;
	wire new_net_46;
	wire new_net_729;
	wire new_net_780;
	wire new_net_1078;
	wire new_net_3314;
	wire new_net_3429;
	wire new_net_1616;
	wire new_net_3178;
	wire _0679_;
	wire new_net_1786;
	wire new_net_2339;
	wire new_net_2473;
	wire new_net_2600;
	wire _0115_;
	wire new_net_1650;
	wire new_net_3215;
	wire new_net_2314;
	wire new_net_2788;
	wire new_net_1928;
	wire new_net_2312;
	wire new_net_94;
	wire new_net_256;
	wire new_net_292;
	wire new_net_346;
	wire new_net_397;
	wire new_net_466;
	wire new_net_484;
	wire new_net_538;
	wire new_net_679;
	wire new_net_748;
	wire new_net_2213;
	wire new_net_492;
	wire new_net_1285;
	wire new_net_3289;
	wire new_net_3378;
	wire new_net_1050;
	wire new_net_1567;
	wire new_net_1834;
	wire new_net_3082;
	wire new_net_3237;
	wire new_net_1111;
	wire new_net_2221;
	wire new_net_41;
	wire new_net_23;
	wire new_net_797;
	wire new_net_1104;
	wire new_net_1234;
	wire new_net_1301;
	wire new_net_1343;
	wire new_net_1364;
	wire new_net_1406;
	wire new_net_1471;
	wire new_net_2084;
	wire new_net_518;
	wire new_net_2464;
	wire new_net_2581;
	wire new_net_2842;
	wire new_net_1913;
	wire new_net_1316;
	wire new_net_3208;
	wire new_net_2811;
	wire new_net_3351;
	wire new_net_1087;
	wire new_net_1818;
	wire new_net_3095;
	wire new_net_2342;
	wire new_net_129;
	wire new_net_450;
	wire new_net_867;
	wire new_net_936;
	wire new_net_972;
	wire new_net_990;
	wire new_net_1235;
	wire new_net_1552;
	wire new_net_1622;
	wire new_net_1933;
	wire new_net_3137;
	wire new_net_2416;
	wire new_net_2876;
	wire new_net_2817;
	wire new_net_883;
	wire new_net_2128;
	wire new_net_2481;
	wire new_net_2141;
	wire new_net_1824;
	wire new_net_2796;
	wire new_net_1347;
	wire new_net_1405;
	wire new_net_2280;
	wire new_net_3154;
	wire new_net_364;
	wire new_net_76;
	wire new_net_433;
	wire new_net_643;
	wire new_net_919;
	wire new_net_1061;
	wire new_net_1114;
	wire new_net_1140;
	wire new_net_1829;
	wire new_net_1858;
	wire new_net_2769;
	wire new_net_2952;
	wire new_net_1909;
	wire new_net_1669;
	wire new_net_2689;
	wire _0336_;
	wire new_net_2871;
	wire new_net_2963;
	wire new_net_1378;
	wire new_net_3425;
	wire new_net_380;
	wire new_net_398;
	wire new_net_95;
	wire new_net_257;
	wire new_net_293;
	wire new_net_329;
	wire _0353_;
	wire new_net_485;
	wire new_net_539;
	wire new_net_626;
	wire new_net_1864;
	wire new_net_2170;
	wire _0377_;
	wire new_net_2201;
	wire new_net_2305;
	wire new_net_2663;
	wire new_net_2555;
	wire _0401_;
	wire new_net_820;
	wire new_net_3319;
	wire _0394_;
	wire new_net_749;
	wire new_net_203;
	wire new_net_3183;
	wire _0418_;
	wire new_net_1461;
	wire new_net_2306;
	wire _0703_;
	wire new_net_1164;
	wire new_net_24;
	wire new_net_42;
	wire new_net_222;
	wire new_net_798;
	wire new_net_1245;
	wire new_net_1333;
	wire new_net_1375;
	wire new_net_1417;
	wire new_net_1459;
	wire new_net_1516;
	wire new_net_2862;
	wire new_net_3220;
	wire new_net_2799;
	wire _0720_;
	wire new_net_1279;
	wire new_net_2679;
	wire new_net_774;
	wire new_net_3294;
	wire _0744_;
	wire new_net_2652;
	wire new_net_2801;
	wire new_net_2055;
	wire new_net_2461;
	wire new_net_2723;
	wire new_net_2000;
	wire new_net_1232;
	wire new_net_3057;
	wire _0761_;
	wire new_net_3383;
	wire new_net_187;
	wire new_net_274;
	wire new_net_556;
	wire new_net_574;
	wire new_net_730;
	wire new_net_781;
	wire new_net_868;
	wire new_net_973;
	wire _0785_;
	wire new_net_991;
	wire new_net_1434;
	wire new_net_2130;
	wire new_net_2803;
	wire new_net_3029;
	wire new_net_3169;
	wire new_net_2734;
	wire new_net_2922;
	wire new_net_3091;
	wire new_net_2586;
	wire new_net_1004;
	wire new_net_1310;
	wire new_net_2268;
	wire new_net_3089;
	wire new_net_1819;
	wire new_net_2445;
	wire new_net_2014;
	wire _0231_;
	wire new_net_1011;
	wire new_net_347;
	wire new_net_77;
	wire new_net_434;
	wire new_net_467;
	wire new_net_644;
	wire new_net_680;
	wire new_net_920;
	wire new_net_1184;
	wire new_net_1204;
	wire new_net_1626;
	wire new_net_1821;
	wire new_net_3144;
	wire new_net_2709;
	wire new_net_2045;
	wire new_net_479;
	wire _0272_;
	wire new_net_1247;
	wire new_net_2129;
	wire new_net_2877;
	wire new_net_1157;
	wire new_net_3078;
	wire new_net_2146;
	wire new_net_3333;
	wire new_net_96;
	wire new_net_294;
	wire new_net_330;
	wire new_net_381;
	wire new_net_399;
	wire new_net_486;
	wire new_net_540;
	wire new_net_627;
	wire _0313_;
	wire new_net_1167;
	wire new_net_1691;
	wire new_net_2572;
	wire _0598_;
	wire new_net_1634;
	wire _0622_;
	wire new_net_2957;
	wire new_net_2774;
	wire new_net_724;
	wire new_net_2541;
	wire _0639_;
	wire new_net_660;
	wire new_net_2878;
	wire new_net_130;
	wire new_net_223;
	wire new_net_43;
	wire new_net_451;
	wire _0075_;
	wire _0663_;
	wire new_net_799;
	wire new_net_937;
	wire new_net_1302;
	wire new_net_1344;
	wire new_net_1949;
	wire new_net_2090;
	wire new_net_2373;
	wire new_net_2095;
	wire new_net_1076;
	wire _0680_;
	wire new_net_3193;
	wire new_net_3432;
	wire new_net_2237;
	wire new_net_2520;
	wire new_net_2066;
	wire new_net_3008;
	wire new_net_1339;
	wire new_net_1397;
	wire new_net_188;
	wire new_net_275;
	wire new_net_365;
	wire new_net_557;
	wire _0133_;
	wire new_net_575;
	wire new_net_731;
	wire new_net_782;
	wire new_net_974;
	wire new_net_1080;
	wire new_net_1728;
	wire new_net_2241;
	wire new_net_2755;
	wire new_net_3188;
	wire new_net_1139;
	wire new_net_908;
	wire _0442_;
	wire new_net_3109;
	wire new_net_1255;
	wire new_net_1526;
	wire new_net_915;
	wire new_net_1491;
	wire new_net_510;
	wire new_net_1883;
	wire new_net_258;
	wire new_net_348;
	wire new_net_78;
	wire new_net_468;
	wire new_net_645;
	wire new_net_681;
	wire new_net_1119;
	wire new_net_921;
	wire new_net_1370;
	wire _0476_;
	wire new_net_1428;
	wire new_net_2728;
	wire new_net_2506;
	wire new_net_2005;
	wire new_net_3085;
	wire new_net_3062;
	wire new_net_3055;
	wire new_net_3305;
	wire _0517_;
	wire new_net_113;
	wire new_net_2632;
	wire new_net_2739;
	wire new_net_3174;
	wire new_net_1815;
	wire new_net_3401;
	wire new_net_2699;
	wire new_net_25;
	wire new_net_97;
	wire new_net_331;
	wire new_net_382;
	wire new_net_400;
	wire new_net_541;
	wire new_net_755;
	wire new_net_1215;
	wire new_net_1517;
	wire new_net_1621;
	wire new_net_1544;
	wire new_net_1401;
	wire _0558_;
	wire new_net_2346;
	wire new_net_3040;
	wire new_net_3074;
	wire new_net_762;
	wire new_net_1684;
	wire new_net_2642;
	wire new_net_3327;
	wire new_net_2714;
	wire new_net_2727;
	wire new_net_131;
	wire new_net_224;
	wire new_net_452;
	wire new_net_800;
	wire new_net_869;
	wire new_net_901;
	wire new_net_938;
	wire new_net_992;
	wire new_net_1154;
	wire new_net_1244;
	wire new_net_2116;
	wire new_net_1937;
	wire new_net_3155;
	wire new_net_1698;
	wire new_net_1696;
	wire new_net_2577;
	wire new_net_3264;
	wire new_net_2227;
	wire new_net_189;
	wire new_net_276;
	wire new_net_366;
	wire new_net_435;
	wire new_net_576;
	wire _0354_;
	wire new_net_732;
	wire new_net_1194;
	wire new_net_1200;
	wire new_net_1627;
	wire new_net_2544;
	wire new_net_2966;
	wire _0378_;
	wire new_net_810;
	wire new_net_2883;
	wire new_net_1249;
	wire new_net_1489;
	wire new_net_2378;
	wire _0402_;
	wire new_net_1587;
	wire new_net_1457;
	wire new_net_2065;
	wire new_net_1863;
	wire _0395_;
	wire new_net_817;
	wire new_net_1623;
	wire new_net_2210;
	wire new_net_2100;
	wire _0419_;
	wire new_net_829;
	wire new_net_79;
	wire new_net_295;
	wire new_net_259;
	wire new_net_349;
	wire _0704_;
	wire new_net_487;
	wire new_net_628;
	wire new_net_646;
	wire new_net_688;
	wire new_net_751;
	wire new_net_838;
	wire new_net_2525;
	wire new_net_3015;
	wire new_net_2426;
	wire new_net_3043;
	wire _0436_;
	wire new_net_3013;
	wire _0721_;
	wire new_net_695;
	wire new_net_2050;
	wire new_net_2251;
	wire new_net_3195;
	wire new_net_845;
	wire new_net_2760;
	wire new_net_1628;
	wire _0745_;
	wire new_net_3227;
	wire new_net_2865;
	wire new_net_1430;
	wire new_net_2371;
	wire new_net_3197;
	wire new_net_3114;
	wire new_net_2804;
	wire new_net_26;
	wire _0762_;
	wire new_net_44;
	wire new_net_98;
	wire new_net_332;
	wire new_net_383;
	wire new_net_542;
	wire new_net_1148;
	wire new_net_789;
	wire new_net_1531;
	wire new_net_2465;
	wire _0786_;
	wire new_net_1306;
	wire new_net_2993;
	wire new_net_3421;
	wire new_net_2808;
	wire new_net_2442;
	wire new_net_1811;
	wire new_net_2012;
	wire new_net_1579;
	wire new_net_3422;
	wire new_net_1894;
	wire new_net_675;
	wire new_net_132;
	wire new_net_225;
	wire new_net_453;
	wire new_net_558;
	wire new_net_783;
	wire new_net_801;
	wire new_net_870;
	wire new_net_939;
	wire new_net_1303;
	wire new_net_993;
	wire new_net_1992;
	wire new_net_2746;
	wire new_net_2793;
	wire new_net_1646;
	wire new_net_2672;
	wire new_net_1031;
	wire new_net_1855;
	wire _0273_;
	wire new_net_3408;
	wire new_net_1874;
	wire new_net_2566;
	wire _0582_;
	wire new_net_2904;
	wire new_net_367;
	wire new_net_2;
	wire new_net_190;
	wire new_net_277;
	wire new_net_436;
	wire new_net_469;
	wire new_net_577;
	wire new_net_682;
	wire new_net_733;
	wire new_net_1115;
	wire new_net_2647;
	wire _0314_;
	wire new_net_2719;
	wire _0599_;
	wire new_net_2868;
	wire new_net_2626;
	wire new_net_2121;
	wire _0623_;
	wire new_net_1638;
	wire new_net_2297;
	wire new_net_3160;
	wire new_net_1703;
	wire new_net_2296;
	wire new_net_1256;
	wire new_net_2086;
	wire new_net_2261;
	wire new_net_2331;
	wire new_net_3028;
	wire _0640_;
	wire new_net_1136;
	wire new_net_1841;
	wire new_net_401;
	wire new_net_350;
	wire new_net_80;
	wire new_net_296;
	wire new_net_488;
	wire new_net_629;
	wire new_net_752;
	wire _0664_;
	wire new_net_923;
	wire new_net_1518;
	wire new_net_47;
	wire new_net_3273;
	wire new_net_2703;
	wire _0681_;
	wire new_net_2890;
	wire new_net_1393;
	wire new_net_2972;
	wire new_net_2888;
	wire _0117_;
	wire new_net_2385;
	wire new_net_2705;
	wire new_net_1867;
	wire new_net_45;
	wire new_net_333;
	wire new_net_384;
	wire new_net_543;
	wire new_net_1110;
	wire new_net_1575;
	wire new_net_1679;
	wire _0134_;
	wire new_net_1269;
	wire new_net_1794;
	wire new_net_2107;
	wire new_net_493;
	wire new_net_2532;
	wire new_net_2650;
	wire new_net_2826;
	wire _0443_;
	wire new_net_2458;
	wire new_net_2047;
	wire new_net_3020;
	wire new_net_3047;
	wire _0175_;
	wire new_net_500;
	wire new_net_2400;
	wire _0460_;
	wire new_net_1424;
	wire new_net_2694;
	wire new_net_2049;
	wire new_net_1805;
	wire new_net_2765;
	wire new_net_133;
	wire new_net_559;
	wire new_net_784;
	wire _0484_;
	wire new_net_802;
	wire new_net_926;
	wire new_net_940;
	wire new_net_976;
	wire new_net_994;
	wire new_net_1335;
	wire new_net_3026;
	wire new_net_3121;
	wire _0477_;
	wire new_net_2264;
	wire new_net_2158;
	wire new_net_519;
	wire new_net_3241;
	wire _0501_;
	wire new_net_2438;
	wire _0518_;
	wire new_net_1449;
	wire new_net_1108;
	wire new_net_1509;
	wire new_net_3106;
	wire new_net_2015;
	wire new_net_4;
	wire new_net_191;
	wire new_net_260;
	wire _0542_;
	wire new_net_437;
	wire new_net_470;
	wire new_net_647;
	wire new_net_683;
	wire new_net_734;
	wire new_net_1081;
	wire new_net_1791;
	wire new_net_2516;
	wire new_net_1822;
	wire new_net_1124;
	wire new_net_1513;
	wire new_net_2605;
	wire _0559_;
	wire new_net_884;
	wire new_net_2693;
	wire new_net_2751;
	wire new_net_2934;
	wire new_net_2421;
	wire new_net_140;
	wire new_net_2176;
	wire new_net_1687;
	wire new_net_3410;
	wire new_net_81;
	wire new_net_27;
	wire new_net_99;
	wire new_net_402;
	wire new_net_351;
	wire new_net_630;
	wire new_net_924;
	wire new_net_1555;
	wire new_net_2085;
	wire new_net_2182;
	wire new_net_2257;
	wire new_net_2984;
	wire new_net_1879;
	wire new_net_2185;
	wire new_net_1967;
	wire _0321_;
	wire new_net_2291;
	wire new_net_2619;
	wire new_net_2909;
	wire new_net_1298;
	wire new_net_1356;
	wire new_net_1996;
	wire new_net_1607;
	wire _0053_;
	wire new_net_2502;
	wire new_net_3263;
	wire new_net_2575;
	wire new_net_2126;
	wire _0362_;
	wire new_net_226;
	wire new_net_334;
	wire new_net_385;
	wire new_net_454;
	wire new_net_1085;
	wire new_net_1182;
	wire new_net_1220;
	wire new_net_1710;
	wire _0355_;
	wire new_net_1708;
	wire new_net_2847;
	wire new_net_2779;
	wire new_net_3337;
	wire new_net_1920;
	wire new_net_3392;
	wire new_net_2336;
	wire new_net_3001;
	wire new_net_2172;
	wire new_net_3356;
	wire _0403_;
	wire new_net_821;
	wire new_net_1192;
	wire new_net_3005;
	wire new_net_3278;
	wire new_net_3433;
	wire new_net_550;
	wire new_net_1329;
	wire _0396_;
	wire new_net_1387;
	wire new_net_204;
	wire _0420_;
	input G1;
	input G10;
	input G11;
	input G12;
	input G13;
	input G14;
	input G15;
	input G16;
	input G17;
	input G18;
	input G19;
	input G2;
	input G20;
	input G21;
	input G22;
	input G23;
	input G24;
	input G25;
	input G26;
	input G27;
	input G28;
	input G29;
	input G3;
	input G30;
	input G31;
	input G32;
	input G33;
	input G34;
	input G35;
	input G36;
	input G37;
	input G38;
	input G39;
	input G4;
	input G40;
	input G41;
	input G42;
	input G43;
	input G44;
	input G45;
	input G46;
	input G47;
	input G48;
	input G49;
	input G5;
	input G50;
	input G6;
	input G7;
	input G8;
	input G9;
	output G3519;
	output G3520;
	output G3521;
	output G3522;
	output G3523;
	output G3524;
	output G3525;
	output G3526;
	output G3527;
	output G3528;
	output G3529;
	output G3530;
	output G3531;
	output G3532;
	output G3533;
	output G3534;
	output G3535;
	output G3536;
	output G3537;
	output G3538;
	output G3539;
	output G3540;

	inv _0798_ (
		.din(new_net_52),
		.dout(_0620_)
	);

	and_ii _0799_ (
		.a(new_net_350),
		.b(new_net_595),
		.c(_0631_)
	);

	or_bb _0800_ (
		.a(new_net_772),
		.b(new_net_523),
		.c(new_net_1475)
	);

	and_ii _0801_ (
		.a(new_net_663),
		.b(new_net_36),
		.c(_0652_)
	);

	and_bi _0802_ (
		.a(new_net_217),
		.b(new_net_260),
		.c(_0662_)
	);

	and_bi _0803_ (
		.a(new_net_136),
		.b(new_net_16),
		.c(_0673_)
	);

	and_ii _0804_ (
		.a(new_net_1255),
		.b(_0662_),
		.c(_0684_)
	);

	or_bi _0805_ (
		.a(new_net_597),
		.b(new_net_406),
		.c(_0695_)
	);

	and_bi _0806_ (
		.a(new_net_435),
		.b(new_net_842),
		.c(_0705_)
	);

	or_bi _0807_ (
		.a(new_net_1256),
		.b(_0695_),
		.c(_0716_)
	);

	and_bi _0808_ (
		.a(_0684_),
		.b(_0716_),
		.c(_0727_)
	);

	and_bi _0809_ (
		.a(new_net_292),
		.b(new_net_59),
		.c(_0736_)
	);

	and_bi _0810_ (
		.a(new_net_789),
		.b(new_net_348),
		.c(_0746_)
	);

	or_bb _0811_ (
		.a(_0746_),
		.b(_0736_),
		.c(_0756_)
	);

	and_bi _0812_ (
		.a(new_net_240),
		.b(new_net_890),
		.c(_0764_)
	);

	and_bi _0813_ (
		.a(new_net_86),
		.b(new_net_283),
		.c(_0775_)
	);

	or_bb _0814_ (
		.a(_0775_),
		.b(_0764_),
		.c(_0785_)
	);

	or_bb _0815_ (
		.a(_0785_),
		.b(_0756_),
		.c(_0788_)
	);

	and_bi _0816_ (
		.a(_0727_),
		.b(new_net_1257),
		.c(_0789_)
	);

	or_bb _0817_ (
		.a(_0789_),
		.b(new_net_46),
		.c(_0790_)
	);

	inv _0818_ (
		.din(new_net_31),
		.dout(_0791_)
	);

	or_bi _0819_ (
		.a(new_net_666),
		.b(new_net_494),
		.c(_0792_)
	);

	and_bi _0820_ (
		.a(new_net_685),
		.b(new_net_230),
		.c(_0793_)
	);

	inv _0821_ (
		.din(new_net_285),
		.dout(_0794_)
	);

	and_ii _0822_ (
		.a(new_net_261),
		.b(new_net_14),
		.c(_0795_)
	);

	and_bi _0823_ (
		.a(new_net_717),
		.b(new_net_946),
		.c(_0796_)
	);

	and_bb _0824_ (
		.a(new_net_183),
		.b(new_net_770),
		.c(_0797_)
	);

	and_bi _0825_ (
		.a(new_net_48),
		.b(new_net_495),
		.c(_0000_)
	);

	inv _0826_ (
		.din(new_net_290),
		.dout(_0001_)
	);

	and_ii _0827_ (
		.a(new_net_408),
		.b(new_net_793),
		.c(_0002_)
	);

	or_bb _0828_ (
		.a(new_net_1258),
		.b(new_net_25),
		.c(_0003_)
	);

	and_bi _0829_ (
		.a(new_net_1016),
		.b(new_net_1259),
		.c(_0004_)
	);

	or_bb _0830_ (
		.a(_0004_),
		.b(new_net_1260),
		.c(_0005_)
	);

	and_bi _0831_ (
		.a(new_net_1261),
		.b(_0005_),
		.c(new_net_1481)
	);

	or_bb _0832_ (
		.a(new_net_436),
		.b(new_net_405),
		.c(_0006_)
	);

	and_bb _0833_ (
		.a(new_net_438),
		.b(new_net_407),
		.c(_0007_)
	);

	and_bi _0834_ (
		.a(_0006_),
		.b(_0007_),
		.c(_0008_)
	);

	and_bi _0835_ (
		.a(new_net_293),
		.b(new_net_794),
		.c(_0009_)
	);

	and_bi _0836_ (
		.a(new_net_790),
		.b(new_net_289),
		.c(_0010_)
	);

	and_ii _0837_ (
		.a(_0010_),
		.b(_0009_),
		.c(_0011_)
	);

	or_bi _0838_ (
		.a(new_net_360),
		.b(new_net_489),
		.c(_0012_)
	);

	and_bi _0839_ (
		.a(new_net_361),
		.b(new_net_490),
		.c(_0013_)
	);

	and_bi _0840_ (
		.a(_0012_),
		.b(_0013_),
		.c(_0014_)
	);

	and_bi _0841_ (
		.a(new_net_88),
		.b(new_net_138),
		.c(_0015_)
	);

	and_bi _0842_ (
		.a(new_net_134),
		.b(new_net_83),
		.c(_0016_)
	);

	and_ii _0843_ (
		.a(_0016_),
		.b(_0015_),
		.c(_0017_)
	);

	and_ii _0844_ (
		.a(new_net_241),
		.b(new_net_219),
		.c(_0018_)
	);

	and_bb _0845_ (
		.a(new_net_244),
		.b(new_net_220),
		.c(_0019_)
	);

	and_ii _0846_ (
		.a(_0019_),
		.b(_0018_),
		.c(_0020_)
	);

	and_bi _0847_ (
		.a(new_net_389),
		.b(new_net_103),
		.c(_0021_)
	);

	and_bi _0848_ (
		.a(new_net_104),
		.b(new_net_390),
		.c(_0022_)
	);

	and_ii _0849_ (
		.a(_0022_),
		.b(_0021_),
		.c(_0023_)
	);

	or_bb _0850_ (
		.a(new_net_89),
		.b(new_net_712),
		.c(_0024_)
	);

	and_bb _0851_ (
		.a(new_net_90),
		.b(new_net_713),
		.c(_0025_)
	);

	and_bi _0852_ (
		.a(_0024_),
		.b(_0025_),
		.c(new_net_1477)
	);

	and_bb _0853_ (
		.a(new_net_264),
		.b(new_net_18),
		.c(_0026_)
	);

	and_ii _0854_ (
		.a(new_net_1262),
		.b(new_net_947),
		.c(_0027_)
	);

	or_bb _0855_ (
		.a(new_net_284),
		.b(new_net_896),
		.c(_0028_)
	);

	and_bb _0856_ (
		.a(new_net_278),
		.b(new_net_892),
		.c(_0029_)
	);

	and_bi _0857_ (
		.a(new_net_67),
		.b(new_net_1263),
		.c(_0030_)
	);

	or_bi _0858_ (
		.a(new_net_274),
		.b(new_net_552),
		.c(_0031_)
	);

	and_bi _0859_ (
		.a(new_net_277),
		.b(new_net_553),
		.c(_0032_)
	);

	and_bi _0860_ (
		.a(_0031_),
		.b(_0032_),
		.c(_0033_)
	);

	and_bi _0861_ (
		.a(new_net_596),
		.b(new_net_60),
		.c(_0034_)
	);

	and_bi _0862_ (
		.a(new_net_53),
		.b(new_net_592),
		.c(_0035_)
	);

	and_ii _0863_ (
		.a(_0035_),
		.b(_0034_),
		.c(_0036_)
	);

	and_ii _0864_ (
		.a(new_net_347),
		.b(new_net_843),
		.c(_0037_)
	);

	and_bb _0865_ (
		.a(new_net_351),
		.b(new_net_848),
		.c(_0038_)
	);

	and_ii _0866_ (
		.a(_0038_),
		.b(_0037_),
		.c(_0039_)
	);

	and_ii _0867_ (
		.a(new_net_699),
		.b(new_net_1001),
		.c(_0040_)
	);

	and_bb _0868_ (
		.a(new_net_700),
		.b(new_net_1002),
		.c(_0041_)
	);

	and_ii _0869_ (
		.a(_0041_),
		.b(_0040_),
		.c(_0042_)
	);

	or_bb _0870_ (
		.a(new_net_1020),
		.b(new_net_272),
		.c(_0043_)
	);

	and_bb _0871_ (
		.a(new_net_1021),
		.b(new_net_273),
		.c(_0044_)
	);

	and_bi _0872_ (
		.a(_0043_),
		.b(_0044_),
		.c(new_net_1463)
	);

	and_bi _0873_ (
		.a(new_net_37),
		.b(new_net_231),
		.c(_0045_)
	);

	or_bb _0874_ (
		.a(new_net_91),
		.b(new_net_279),
		.c(_0046_)
	);

	and_bi _0875_ (
		.a(new_net_39),
		.b(new_net_664),
		.c(_0047_)
	);

	or_ii _0876_ (
		.a(new_net_491),
		.b(new_net_658),
		.c(_0048_)
	);

	or_ii _0877_ (
		.a(new_net_665),
		.b(new_net_38),
		.c(_0049_)
	);

	and_bi _0878_ (
		.a(new_net_155),
		.b(_0049_),
		.c(_0050_)
	);

	or_bi _0879_ (
		.a(_0050_),
		.b(new_net_269),
		.c(_0051_)
	);

	and_ii _0880_ (
		.a(new_net_393),
		.b(new_net_578),
		.c(_0052_)
	);

	and_bi _0881_ (
		.a(new_net_286),
		.b(new_net_447),
		.c(_0053_)
	);

	and_bi _0882_ (
		.a(new_net_1264),
		.b(_0053_),
		.c(_0054_)
	);

	and_bi _0883_ (
		.a(new_net_948),
		.b(new_net_287),
		.c(_0055_)
	);

	or_bb _0884_ (
		.a(_0055_),
		.b(new_net_686),
		.c(_0056_)
	);

	or_bb _0885_ (
		.a(new_net_152),
		.b(new_net_40),
		.c(_0057_)
	);

	and_bi _0886_ (
		.a(new_net_613),
		.b(new_net_937),
		.c(_0058_)
	);

	inv _0887_ (
		.din(new_net_17),
		.dout(_0059_)
	);

	or_bi _0888_ (
		.a(new_net_32),
		.b(new_net_149),
		.c(_0060_)
	);

	and_bi _0889_ (
		.a(new_net_800),
		.b(new_net_656),
		.c(_0061_)
	);

	or_bb _0890_ (
		.a(_0061_),
		.b(new_net_1265),
		.c(_0062_)
	);

	and_bi _0891_ (
		.a(new_net_1266),
		.b(_0062_),
		.c(_0063_)
	);

	and_bi _0892_ (
		.a(new_net_394),
		.b(_0063_),
		.c(_0064_)
	);

	or_bb _0893_ (
		.a(_0064_),
		.b(_0054_),
		.c(_0065_)
	);

	or_bb _0894_ (
		.a(new_net_859),
		.b(new_net_804),
		.c(_0066_)
	);

	or_bb _0895_ (
		.a(new_net_127),
		.b(new_net_246),
		.c(_0067_)
	);

	and_bi _0896_ (
		.a(new_net_1267),
		.b(new_net_659),
		.c(_0068_)
	);

	and_bb _0897_ (
		.a(new_net_163),
		.b(new_net_128),
		.c(_0069_)
	);

	or_bb _0898_ (
		.a(new_net_234),
		.b(new_net_270),
		.c(_0070_)
	);

	or_ii _0899_ (
		.a(new_net_332),
		.b(new_net_692),
		.c(_0071_)
	);

	and_bi _0900_ (
		.a(new_net_250),
		.b(new_net_723),
		.c(_0072_)
	);

	or_bi _0901_ (
		.a(new_net_253),
		.b(new_net_87),
		.c(_0073_)
	);

	or_bb _0902_ (
		.a(new_net_1268),
		.b(new_net_156),
		.c(_0074_)
	);

	and_bi _0903_ (
		.a(new_net_1269),
		.b(new_net_414),
		.c(_0075_)
	);

	or_bi _0904_ (
		.a(new_net_176),
		.b(new_net_891),
		.c(_0076_)
	);

	or_ii _0905_ (
		.a(new_net_602),
		.b(new_net_172),
		.c(_0077_)
	);

	or_ii _0906_ (
		.a(new_net_1270),
		.b(new_net_631),
		.c(_0078_)
	);

	or_bb _0907_ (
		.a(_0078_),
		.b(_0075_),
		.c(_0079_)
	);

	and_bi _0908_ (
		.a(new_net_1271),
		.b(_0079_),
		.c(_0080_)
	);

	and_bi _0909_ (
		.a(new_net_334),
		.b(_0080_),
		.c(_0081_)
	);

	or_bb _0910_ (
		.a(new_net_1272),
		.b(new_net_427),
		.c(_0082_)
	);

	and_bi _0911_ (
		.a(new_net_144),
		.b(new_net_316),
		.c(_0083_)
	);

	or_bb _0912_ (
		.a(_0083_),
		.b(new_net_70),
		.c(_0084_)
	);

	and_ii _0913_ (
		.a(new_net_203),
		.b(new_net_419),
		.c(_0085_)
	);

	or_bb _0914_ (
		.a(new_net_1031),
		.b(new_net_317),
		.c(_0086_)
	);

	and_bi _0915_ (
		.a(new_net_72),
		.b(_0086_),
		.c(_0087_)
	);

	and_bi _0916_ (
		.a(new_net_785),
		.b(new_net_465),
		.c(_0088_)
	);

	or_bb _0917_ (
		.a(new_net_448),
		.b(new_net_802),
		.c(_0089_)
	);

	and_bi _0918_ (
		.a(new_net_796),
		.b(new_net_92),
		.c(_0090_)
	);

	or_bi _0919_ (
		.a(new_net_1273),
		.b(_0089_),
		.c(_0091_)
	);

	or_ii _0920_ (
		.a(new_net_275),
		.b(new_net_33),
		.c(_0092_)
	);

	inv _0921_ (
		.din(new_net_265),
		.dout(_0093_)
	);

	and_bi _0922_ (
		.a(new_net_902),
		.b(new_net_652),
		.c(_0094_)
	);

	and_bi _0923_ (
		.a(new_net_673),
		.b(new_net_41),
		.c(_0095_)
	);

	and_bi _0924_ (
		.a(new_net_1043),
		.b(new_net_157),
		.c(_0096_)
	);

	or_bb _0925_ (
		.a(new_net_1274),
		.b(_0094_),
		.c(_0097_)
	);

	and_bi _0926_ (
		.a(new_net_1275),
		.b(_0097_),
		.c(_0098_)
	);

	and_bi _0927_ (
		.a(new_net_398),
		.b(_0098_),
		.c(_0099_)
	);

	or_bi _0928_ (
		.a(_0099_),
		.b(_0091_),
		.c(_0100_)
	);

	or_bi _0929_ (
		.a(new_net_254),
		.b(new_net_137),
		.c(_0101_)
	);

	and_bi _0930_ (
		.a(new_net_603),
		.b(new_net_411),
		.c(_0102_)
	);

	or_bb _0931_ (
		.a(new_net_164),
		.b(new_net_58),
		.c(_0103_)
	);

	and_bi _0932_ (
		.a(new_net_150),
		.b(new_net_84),
		.c(_0104_)
	);

	and_bi _0933_ (
		.a(new_net_883),
		.b(new_net_1276),
		.c(_0105_)
	);

	or_bb _0934_ (
		.a(new_net_1277),
		.b(_0102_),
		.c(_0106_)
	);

	and_bi _0935_ (
		.a(new_net_1278),
		.b(_0106_),
		.c(_0107_)
	);

	and_bi _0936_ (
		.a(new_net_329),
		.b(_0107_),
		.c(_0108_)
	);

	or_bb _0937_ (
		.a(new_net_1279),
		.b(new_net_428),
		.c(_0109_)
	);

	and_bi _0938_ (
		.a(new_net_140),
		.b(new_net_1039),
		.c(_0110_)
	);

	or_bb _0939_ (
		.a(_0110_),
		.b(new_net_533),
		.c(_0111_)
	);

	or_bb _0940_ (
		.a(new_net_1040),
		.b(new_net_1033),
		.c(_0112_)
	);

	and_bi _0941_ (
		.a(new_net_535),
		.b(_0112_),
		.c(_0113_)
	);

	and_bi _0942_ (
		.a(new_net_1280),
		.b(new_net_375),
		.c(_0114_)
	);

	and_bb _0943_ (
		.a(new_net_205),
		.b(new_net_193),
		.c(_0115_)
	);

	inv _0944_ (
		.din(new_net_893),
		.dout(_0116_)
	);

	and_bi _0945_ (
		.a(new_net_395),
		.b(new_net_687),
		.c(_0117_)
	);

	and_ii _0946_ (
		.a(new_net_574),
		.b(new_net_450),
		.c(_0118_)
	);

	or_bb _0947_ (
		.a(_0118_),
		.b(new_net_502),
		.c(_0119_)
	);

	and_bi _0948_ (
		.a(new_net_97),
		.b(new_net_897),
		.c(_0120_)
	);

	or_bb _0949_ (
		.a(new_net_939),
		.b(new_net_15),
		.c(_0121_)
	);

	and_bi _0950_ (
		.a(new_net_525),
		.b(new_net_657),
		.c(_0122_)
	);

	and_bi _0951_ (
		.a(new_net_1281),
		.b(_0122_),
		.c(_0123_)
	);

	and_bi _0952_ (
		.a(new_net_399),
		.b(_0123_),
		.c(_0124_)
	);

	or_bb _0953_ (
		.a(_0124_),
		.b(new_net_1282),
		.c(_0125_)
	);

	or_bi _0954_ (
		.a(_0125_),
		.b(_0119_),
		.c(_0126_)
	);

	or_bi _0955_ (
		.a(new_net_251),
		.b(new_net_242),
		.c(_0127_)
	);

	and_bi _0956_ (
		.a(new_net_139),
		.b(new_net_415),
		.c(_0128_)
	);

	or_bb _0957_ (
		.a(new_net_158),
		.b(new_net_591),
		.c(_0129_)
	);

	and_bi _0958_ (
		.a(new_net_177),
		.b(new_net_221),
		.c(_0130_)
	);

	and_bi _0959_ (
		.a(_0129_),
		.b(_0130_),
		.c(_0131_)
	);

	or_bb _0960_ (
		.a(new_net_1283),
		.b(_0128_),
		.c(_0132_)
	);

	and_bi _0961_ (
		.a(new_net_1284),
		.b(_0132_),
		.c(_0133_)
	);

	and_bi _0962_ (
		.a(new_net_333),
		.b(_0133_),
		.c(_0134_)
	);

	or_bb _0963_ (
		.a(new_net_1285),
		.b(new_net_429),
		.c(_0135_)
	);

	and_bi _0964_ (
		.a(new_net_146),
		.b(new_net_391),
		.c(_0136_)
	);

	or_bb _0965_ (
		.a(_0136_),
		.b(new_net_1045),
		.c(_0137_)
	);

	or_bb _0966_ (
		.a(new_net_392),
		.b(new_net_1034),
		.c(_0138_)
	);

	and_bi _0967_ (
		.a(new_net_1047),
		.b(_0138_),
		.c(_0139_)
	);

	or_bi _0968_ (
		.a(new_net_604),
		.b(new_net_1286),
		.c(_0140_)
	);

	inv _0969_ (
		.din(new_net_93),
		.dout(_0141_)
	);

	and_bi _0970_ (
		.a(new_net_1287),
		.b(new_net_576),
		.c(_0142_)
	);

	or_bb _0971_ (
		.a(new_net_763),
		.b(new_net_262),
		.c(_0143_)
	);

	or_bb _0972_ (
		.a(new_net_940),
		.b(new_net_718),
		.c(_0144_)
	);

	and_bi _0973_ (
		.a(new_net_894),
		.b(new_net_653),
		.c(_0145_)
	);

	and_bi _0974_ (
		.a(new_net_1288),
		.b(_0145_),
		.c(_0146_)
	);

	and_bi _0975_ (
		.a(new_net_396),
		.b(_0146_),
		.c(_0147_)
	);

	and_bi _0976_ (
		.a(new_net_449),
		.b(new_net_907),
		.c(_0148_)
	);

	or_bb _0977_ (
		.a(_0148_),
		.b(_0147_),
		.c(_0149_)
	);

	and_bi _0978_ (
		.a(_0143_),
		.b(new_net_1289),
		.c(_0150_)
	);

	inv _0979_ (
		.din(new_net_218),
		.dout(_0151_)
	);

	or_bb _0980_ (
		.a(new_net_252),
		.b(new_net_258),
		.c(_0152_)
	);

	and_bi _0981_ (
		.a(new_net_85),
		.b(new_net_410),
		.c(_0153_)
	);

	or_bb _0982_ (
		.a(new_net_165),
		.b(new_net_352),
		.c(_0154_)
	);

	and_bi _0983_ (
		.a(new_net_151),
		.b(new_net_135),
		.c(_0155_)
	);

	and_bi _0984_ (
		.a(new_net_340),
		.b(new_net_1290),
		.c(_0156_)
	);

	or_bb _0985_ (
		.a(_0156_),
		.b(_0153_),
		.c(_0157_)
	);

	and_bi _0986_ (
		.a(new_net_1291),
		.b(_0157_),
		.c(_0158_)
	);

	and_bi _0987_ (
		.a(new_net_330),
		.b(_0158_),
		.c(_0159_)
	);

	or_bb _0988_ (
		.a(new_net_1292),
		.b(new_net_430),
		.c(_0160_)
	);

	and_bi _0989_ (
		.a(new_net_141),
		.b(new_net_387),
		.c(_0161_)
	);

	and_bi _0990_ (
		.a(new_net_11),
		.b(_0161_),
		.c(_0162_)
	);

	and_ii _0991_ (
		.a(new_net_388),
		.b(new_net_1032),
		.c(_0163_)
	);

	and_bi _0992_ (
		.a(_0163_),
		.b(new_net_13),
		.c(_0164_)
	);

	or_bb _0993_ (
		.a(new_net_812),
		.b(new_net_869),
		.c(_0165_)
	);

	or_bb _0994_ (
		.a(new_net_862),
		.b(new_net_320),
		.c(_0166_)
	);

	and_bi _0995_ (
		.a(new_net_423),
		.b(new_net_1293),
		.c(_0167_)
	);

	inv _0996_ (
		.din(new_net_968),
		.dout(_0168_)
	);

	and_bi _0997_ (
		.a(new_net_773),
		.b(new_net_54),
		.c(_0169_)
	);

	or_bb _0998_ (
		.a(_0169_),
		.b(new_net_689),
		.c(_0170_)
	);

	and_bi _0999_ (
		.a(new_net_903),
		.b(new_net_938),
		.c(_0171_)
	);

	inv _1000_ (
		.din(new_net_353),
		.dout(_0172_)
	);

	and_bi _1001_ (
		.a(new_net_187),
		.b(new_net_654),
		.c(_0173_)
	);

	or_bb _1002_ (
		.a(_0173_),
		.b(new_net_1294),
		.c(_0174_)
	);

	and_bi _1003_ (
		.a(new_net_1295),
		.b(_0174_),
		.c(_0175_)
	);

	or_bi _1004_ (
		.a(_0175_),
		.b(new_net_400),
		.c(_0176_)
	);

	and_bi _1005_ (
		.a(new_net_159),
		.b(new_net_660),
		.c(_0177_)
	);

	or_bb _1006_ (
		.a(new_net_1296),
		.b(new_net_98),
		.c(_0178_)
	);

	or_bb _1007_ (
		.a(_0178_),
		.b(new_net_397),
		.c(_0179_)
	);

	and_bi _1008_ (
		.a(new_net_61),
		.b(new_net_483),
		.c(_0180_)
	);

	and_bi _1009_ (
		.a(new_net_94),
		.b(new_net_55),
		.c(_0181_)
	);

	or_bb _1010_ (
		.a(new_net_1297),
		.b(_0180_),
		.c(_0182_)
	);

	or_bi _1011_ (
		.a(_0182_),
		.b(new_net_1298),
		.c(_0183_)
	);

	or_bb _1012_ (
		.a(new_net_416),
		.b(new_net_259),
		.c(_0184_)
	);

	or_bb _1013_ (
		.a(new_net_160),
		.b(new_net_844),
		.c(_0185_)
	);

	and_bi _1014_ (
		.a(new_net_178),
		.b(new_net_243),
		.c(_0186_)
	);

	and_bi _1015_ (
		.a(_0185_),
		.b(_0186_),
		.c(_0187_)
	);

	and_bi _1016_ (
		.a(_0184_),
		.b(new_net_1299),
		.c(_0188_)
	);

	or_bb _1017_ (
		.a(new_net_661),
		.b(new_net_247),
		.c(_0189_)
	);

	or_bb _1018_ (
		.a(new_net_226),
		.b(new_net_693),
		.c(_0190_)
	);

	and_ii _1019_ (
		.a(new_net_662),
		.b(new_net_249),
		.c(_0191_)
	);

	and_bi _1020_ (
		.a(new_net_26),
		.b(new_net_73),
		.c(_0192_)
	);

	and_bi _1021_ (
		.a(_0190_),
		.b(_0192_),
		.c(_0193_)
	);

	and_bi _1022_ (
		.a(_0188_),
		.b(new_net_1300),
		.c(_0194_)
	);

	and_bi _1023_ (
		.a(new_net_331),
		.b(_0194_),
		.c(_0195_)
	);

	or_bb _1024_ (
		.a(new_net_99),
		.b(new_net_1035),
		.c(_0196_)
	);

	and_bi _1025_ (
		.a(new_net_833),
		.b(new_net_1301),
		.c(_0197_)
	);

	or_bi _1026_ (
		.a(new_net_100),
		.b(new_net_145),
		.c(_0198_)
	);

	and_bi _1027_ (
		.a(new_net_1302),
		.b(new_net_834),
		.c(_0199_)
	);

	and_ii _1028_ (
		.a(new_net_467),
		.b(new_net_583),
		.c(_0200_)
	);

	and_bi _1029_ (
		.a(new_net_188),
		.b(new_net_95),
		.c(_0201_)
	);

	and_bi _1030_ (
		.a(new_net_486),
		.b(new_net_190),
		.c(_0202_)
	);

	or_bb _1031_ (
		.a(_0202_),
		.b(new_net_1303),
		.c(_0203_)
	);

	and_bb _1032_ (
		.a(new_net_354),
		.b(new_net_598),
		.c(_0204_)
	);

	or_bb _1033_ (
		.a(new_net_1304),
		.b(new_net_774),
		.c(_0205_)
	);

	and_bi _1034_ (
		.a(new_net_575),
		.b(new_net_458),
		.c(_0206_)
	);

	and_bi _1035_ (
		.a(new_net_688),
		.b(new_net_271),
		.c(_0207_)
	);

	and_bb _1036_ (
		.a(new_net_173),
		.b(new_net_599),
		.c(_0208_)
	);

	and_bi _1037_ (
		.a(new_net_632),
		.b(new_net_1305),
		.c(_0209_)
	);

	and_bi _1038_ (
		.a(new_net_950),
		.b(_0209_),
		.c(_0210_)
	);

	or_bb _1039_ (
		.a(new_net_1306),
		.b(_0206_),
		.c(_0211_)
	);

	and_bi _1040_ (
		.a(_0203_),
		.b(new_net_1307),
		.c(_0212_)
	);

	or_bb _1041_ (
		.a(new_net_227),
		.b(new_net_126),
		.c(_0213_)
	);

	and_ii _1042_ (
		.a(new_net_114),
		.b(new_net_724),
		.c(_0214_)
	);

	or_ii _1043_ (
		.a(new_net_115),
		.b(new_net_791),
		.c(_0215_)
	);

	and_bi _1044_ (
		.a(new_net_245),
		.b(new_net_417),
		.c(_0216_)
	);

	or_bb _1045_ (
		.a(new_net_536),
		.b(new_net_168),
		.c(_0217_)
	);

	and_bi _1046_ (
		.a(new_net_166),
		.b(new_net_294),
		.c(_0218_)
	);

	and_bi _1047_ (
		.a(_0217_),
		.b(new_net_1308),
		.c(_0219_)
	);

	or_bb _1048_ (
		.a(new_net_1309),
		.b(_0216_),
		.c(_0220_)
	);

	and_bi _1049_ (
		.a(new_net_1310),
		.b(_0220_),
		.c(_0221_)
	);

	and_bi _1050_ (
		.a(new_net_335),
		.b(_0221_),
		.c(_0222_)
	);

	or_bb _1051_ (
		.a(new_net_1311),
		.b(new_net_588),
		.c(_0223_)
	);

	or_bb _1052_ (
		.a(new_net_609),
		.b(new_net_1036),
		.c(_0224_)
	);

	and_ii _1053_ (
		.a(_0224_),
		.b(new_net_49),
		.c(_0225_)
	);

	and_bi _1054_ (
		.a(new_net_147),
		.b(new_net_610),
		.c(_0226_)
	);

	and_bi _1055_ (
		.a(new_net_50),
		.b(_0226_),
		.c(_0227_)
	);

	or_bb _1056_ (
		.a(new_net_1312),
		.b(new_net_705),
		.c(_0228_)
	);

	and_bi _1057_ (
		.a(new_net_527),
		.b(new_net_856),
		.c(_0229_)
	);

	or_bb _1058_ (
		.a(new_net_764),
		.b(new_net_600),
		.c(_0230_)
	);

	and_bi _1059_ (
		.a(new_net_593),
		.b(new_net_484),
		.c(_0231_)
	);

	and_bb _1060_ (
		.a(new_net_174),
		.b(new_net_847),
		.c(_0232_)
	);

	and_bi _1061_ (
		.a(new_net_884),
		.b(new_net_1313),
		.c(_0233_)
	);

	and_bi _1062_ (
		.a(new_net_952),
		.b(_0233_),
		.c(_0234_)
	);

	or_bb _1063_ (
		.a(new_net_1314),
		.b(_0231_),
		.c(_0235_)
	);

	and_bi _1064_ (
		.a(_0230_),
		.b(_0235_),
		.c(_0236_)
	);

	or_ii _1065_ (
		.a(new_net_117),
		.b(new_net_404),
		.c(_0237_)
	);

	and_bb _1066_ (
		.a(new_net_179),
		.b(new_net_795),
		.c(_0238_)
	);

	and_bi _1067_ (
		.a(new_net_380),
		.b(new_net_161),
		.c(_0239_)
	);

	or_bb _1068_ (
		.a(_0239_),
		.b(_0238_),
		.c(_0240_)
	);

	and_bi _1069_ (
		.a(new_net_291),
		.b(new_net_412),
		.c(_0241_)
	);

	or_bb _1070_ (
		.a(_0241_),
		.b(new_net_1315),
		.c(_0242_)
	);

	and_bi _1071_ (
		.a(new_net_1316),
		.b(_0242_),
		.c(_0243_)
	);

	and_bi _1072_ (
		.a(new_net_336),
		.b(_0243_),
		.c(_0244_)
	);

	or_bb _1073_ (
		.a(new_net_624),
		.b(new_net_590),
		.c(_0245_)
	);

	or_bb _1074_ (
		.a(new_net_682),
		.b(new_net_1037),
		.c(_0246_)
	);

	or_bb _1075_ (
		.a(_0246_),
		.b(new_net_108),
		.c(_0247_)
	);

	and_bi _1076_ (
		.a(new_net_148),
		.b(new_net_683),
		.c(_0248_)
	);

	and_bi _1077_ (
		.a(new_net_110),
		.b(_0248_),
		.c(_0249_)
	);

	and_bi _1078_ (
		.a(new_net_767),
		.b(new_net_1317),
		.c(_0250_)
	);

	or_ii _1079_ (
		.a(new_net_915),
		.b(new_net_879),
		.c(_0251_)
	);

	inv _1080_ (
		.din(new_net_849),
		.dout(_0252_)
	);

	and_bi _1081_ (
		.a(new_net_485),
		.b(new_net_577),
		.c(_0253_)
	);

	or_bb _1082_ (
		.a(_0253_),
		.b(new_net_911),
		.c(_0254_)
	);

	and_bi _1083_ (
		.a(new_net_96),
		.b(new_net_845),
		.c(_0255_)
	);

	and_bb _1084_ (
		.a(new_net_542),
		.b(new_net_175),
		.c(_0256_)
	);

	and_bi _1085_ (
		.a(new_net_341),
		.b(new_net_1318),
		.c(_0257_)
	);

	and_bi _1086_ (
		.a(new_net_951),
		.b(_0257_),
		.c(_0258_)
	);

	or_bb _1087_ (
		.a(_0258_),
		.b(_0255_),
		.c(_0259_)
	);

	and_bi _1088_ (
		.a(_0254_),
		.b(new_net_1319),
		.c(_0260_)
	);

	or_ii _1089_ (
		.a(new_net_116),
		.b(new_net_437),
		.c(_0261_)
	);

	and_bb _1090_ (
		.a(new_net_153),
		.b(new_net_409),
		.c(_0262_)
	);

	and_bi _1091_ (
		.a(new_net_633),
		.b(new_net_169),
		.c(_0263_)
	);

	or_bb _1092_ (
		.a(_0263_),
		.b(_0262_),
		.c(_0264_)
	);

	and_bi _1093_ (
		.a(new_net_792),
		.b(new_net_413),
		.c(_0265_)
	);

	or_bb _1094_ (
		.a(_0265_),
		.b(new_net_1320),
		.c(_0266_)
	);

	and_bi _1095_ (
		.a(new_net_1321),
		.b(_0266_),
		.c(_0267_)
	);

	and_bi _1096_ (
		.a(new_net_337),
		.b(_0267_),
		.c(_0268_)
	);

	or_bb _1097_ (
		.a(new_net_759),
		.b(new_net_589),
		.c(_0269_)
	);

	or_bb _1098_ (
		.a(new_net_925),
		.b(new_net_1038),
		.c(_0270_)
	);

	or_bb _1099_ (
		.a(_0270_),
		.b(new_net_365),
		.c(_0271_)
	);

	or_bb _1100_ (
		.a(new_net_885),
		.b(new_net_680),
		.c(_0272_)
	);

	and_bi _1101_ (
		.a(new_net_880),
		.b(new_net_769),
		.c(_0273_)
	);

	and_bi _1102_ (
		.a(new_net_707),
		.b(new_net_468),
		.c(_0274_)
	);

	or_bb _1103_ (
		.a(_0274_),
		.b(new_net_584),
		.c(_0275_)
	);

	or_bb _1104_ (
		.a(new_net_1322),
		.b(_0273_),
		.c(_0276_)
	);

	and_bi _1105_ (
		.a(_0272_),
		.b(new_net_1323),
		.c(_0277_)
	);

	and_ii _1106_ (
		.a(new_net_120),
		.b(new_net_1013),
		.c(_0278_)
	);

	and_bi _1107_ (
		.a(new_net_606),
		.b(new_net_870),
		.c(_0279_)
	);

	and_ii _1108_ (
		.a(_0279_),
		.b(new_net_814),
		.c(_0280_)
	);

	and_bi _1109_ (
		.a(new_net_424),
		.b(new_net_1324),
		.c(_0281_)
	);

	and_bb _1110_ (
		.a(new_net_376),
		.b(new_net_786),
		.c(_0282_)
	);

	or_bb _1111_ (
		.a(_0282_),
		.b(new_net_466),
		.c(_0283_)
	);

	or_bb _1112_ (
		.a(new_net_1325),
		.b(_0281_),
		.c(_0284_)
	);

	or_bb _1113_ (
		.a(new_net_806),
		.b(_0278_),
		.c(new_net_1465)
	);

	or_ii _1114_ (
		.a(new_net_111),
		.b(new_net_44),
		.c(_0285_)
	);

	and_bi _1115_ (
		.a(new_net_1018),
		.b(new_net_9),
		.c(_0286_)
	);

	inv _1116_ (
		.din(new_net_628),
		.dout(_0287_)
	);

	or_bb _1117_ (
		.a(new_net_760),
		.b(new_net_625),
		.c(_0288_)
	);

	or_bb _1118_ (
		.a(new_net_102),
		.b(new_net_422),
		.c(_0289_)
	);

	or_bb _1119_ (
		.a(_0289_),
		.b(_0288_),
		.c(_0290_)
	);

	or_bb _1120_ (
		.a(_0290_),
		.b(new_net_611),
		.c(_0291_)
	);

	and_bb _1121_ (
		.a(new_net_926),
		.b(new_net_684),
		.c(_0292_)
	);

	or_ii _1122_ (
		.a(new_net_101),
		.b(new_net_420),
		.c(_0293_)
	);

	or_bi _1123_ (
		.a(new_net_1326),
		.b(new_net_612),
		.c(_0294_)
	);

	and_bi _1124_ (
		.a(_0292_),
		.b(_0294_),
		.c(_0295_)
	);

	and_bi _1125_ (
		.a(new_net_1327),
		.b(_0295_),
		.c(_0296_)
	);

	and_bi _1126_ (
		.a(new_net_480),
		.b(_0296_),
		.c(_0297_)
	);

	and_bi _1127_ (
		.a(new_net_142),
		.b(new_net_927),
		.c(_0298_)
	);

	and_bi _1128_ (
		.a(new_net_367),
		.b(_0298_),
		.c(_0299_)
	);

	and_bi _1129_ (
		.a(new_net_886),
		.b(new_net_1328),
		.c(_0300_)
	);

	inv _1130_ (
		.din(new_net_549),
		.dout(_0301_)
	);

	or_bb _1131_ (
		.a(new_net_1329),
		.b(new_net_681),
		.c(_0302_)
	);

	and_bi _1132_ (
		.a(new_net_630),
		.b(new_net_358),
		.c(_0303_)
	);

	or_bb _1133_ (
		.a(_0303_),
		.b(new_net_1330),
		.c(_0304_)
	);

	and_bi _1134_ (
		.a(new_net_996),
		.b(new_net_439),
		.c(_0305_)
	);

	or_bb _1135_ (
		.a(new_net_473),
		.b(new_net_12),
		.c(_0306_)
	);

	and_bi _1136_ (
		.a(new_net_999),
		.b(new_net_863),
		.c(_0307_)
	);

	and_bi _1137_ (
		.a(new_net_864),
		.b(new_net_1000),
		.c(_0308_)
	);

	and_ii _1138_ (
		.a(_0308_),
		.b(_0307_),
		.c(_0309_)
	);

	and_bi _1139_ (
		.a(new_net_1046),
		.b(new_net_472),
		.c(_0310_)
	);

	and_bi _1140_ (
		.a(new_net_322),
		.b(new_net_761),
		.c(_0311_)
	);

	and_bi _1141_ (
		.a(new_net_762),
		.b(new_net_321),
		.c(_0312_)
	);

	or_bb _1142_ (
		.a(_0312_),
		.b(_0311_),
		.c(_0313_)
	);

	or_bb _1143_ (
		.a(new_net_643),
		.b(new_net_708),
		.c(_0314_)
	);

	or_ii _1144_ (
		.a(new_net_1019),
		.b(new_net_112),
		.c(_0315_)
	);

	and_bi _1145_ (
		.a(new_net_534),
		.b(new_net_989),
		.c(_0316_)
	);

	or_bb _1146_ (
		.a(new_net_29),
		.b(new_net_207),
		.c(_0317_)
	);

	and_bb _1147_ (
		.a(new_net_30),
		.b(new_net_206),
		.c(_0318_)
	);

	and_bi _1148_ (
		.a(_0317_),
		.b(_0318_),
		.c(_0319_)
	);

	inv _1149_ (
		.din(new_net_210),
		.dout(_0320_)
	);

	and_ii _1150_ (
		.a(new_net_1331),
		.b(new_net_874),
		.c(_0321_)
	);

	or_ii _1151_ (
		.a(new_net_1007),
		.b(new_net_941),
		.c(_0322_)
	);

	or_bi _1152_ (
		.a(new_net_875),
		.b(new_net_945),
		.c(_0323_)
	);

	and_bb _1153_ (
		.a(new_net_471),
		.b(new_net_813),
		.c(_0324_)
	);

	and_bb _1154_ (
		.a(new_net_481),
		.b(new_net_605),
		.c(_0325_)
	);

	and_ii _1155_ (
		.a(new_net_931),
		.b(new_net_710),
		.c(_0326_)
	);

	and_ii _1156_ (
		.a(_0326_),
		.b(new_net_1332),
		.c(_0327_)
	);

	and_bi _1157_ (
		.a(new_net_213),
		.b(new_net_560),
		.c(_0328_)
	);

	and_bi _1158_ (
		.a(new_net_561),
		.b(new_net_212),
		.c(_0329_)
	);

	or_bb _1159_ (
		.a(new_net_1333),
		.b(new_net_647),
		.c(_0330_)
	);

	and_bi _1160_ (
		.a(new_net_378),
		.b(new_net_1334),
		.c(_0331_)
	);

	and_bi _1161_ (
		.a(new_net_324),
		.b(_0331_),
		.c(_0332_)
	);

	or_bb _1162_ (
		.a(new_net_74),
		.b(new_net_579),
		.c(_0333_)
	);

	and_bi _1163_ (
		.a(new_net_233),
		.b(_0333_),
		.c(_0334_)
	);

	inv _1164_ (
		.din(new_net_129),
		.dout(_0335_)
	);

	and_bi _1165_ (
		.a(new_net_1017),
		.b(new_net_1335),
		.c(_0336_)
	);

	inv _1166_ (
		.din(new_net_1010),
		.dout(_0337_)
	);

	and_bi _1167_ (
		.a(new_net_474),
		.b(new_net_121),
		.c(_0338_)
	);

	and_ii _1168_ (
		.a(new_net_1025),
		.b(new_net_645),
		.c(_0339_)
	);

	or_bb _1169_ (
		.a(new_net_118),
		.b(new_net_932),
		.c(_0340_)
	);

	and_bi _1170_ (
		.a(new_net_943),
		.b(new_net_646),
		.c(_0341_)
	);

	and_bi _1171_ (
		.a(new_net_711),
		.b(_0341_),
		.c(_0342_)
	);

	or_bi _1172_ (
		.a(_0342_),
		.b(new_net_379),
		.c(_0343_)
	);

	or_bi _1173_ (
		.a(new_net_454),
		.b(new_net_181),
		.c(_0344_)
	);

	and_bi _1174_ (
		.a(new_net_455),
		.b(new_net_182),
		.c(_0345_)
	);

	and_bi _1175_ (
		.a(_0344_),
		.b(_0345_),
		.c(_0346_)
	);

	and_bi _1176_ (
		.a(new_net_1015),
		.b(new_net_1027),
		.c(_0347_)
	);

	and_ii _1177_ (
		.a(_0347_),
		.b(new_net_807),
		.c(_0348_)
	);

	or_bi _1178_ (
		.a(new_net_544),
		.b(new_net_944),
		.c(_0349_)
	);

	and_bi _1179_ (
		.a(new_net_585),
		.b(new_net_451),
		.c(_0350_)
	);

	and_bb _1180_ (
		.a(new_net_669),
		.b(new_net_21),
		.c(_0351_)
	);

	and_ii _1181_ (
		.a(_0351_),
		.b(new_net_919),
		.c(_0352_)
	);

	and_ii _1182_ (
		.a(_0352_),
		.b(new_net_580),
		.c(_0353_)
	);

	and_bi _1183_ (
		.a(new_net_20),
		.b(new_net_670),
		.c(_0354_)
	);

	and_bb _1184_ (
		.a(new_net_777),
		.b(new_net_581),
		.c(_0355_)
	);

	or_bi _1185_ (
		.a(new_net_492),
		.b(new_net_170),
		.c(_0356_)
	);

	or_bi _1186_ (
		.a(new_net_236),
		.b(new_net_211),
		.c(_0357_)
	);

	and_bi _1187_ (
		.a(new_net_34),
		.b(new_net_204),
		.c(_0358_)
	);

	or_bb _1188_ (
		.a(new_net_1336),
		.b(new_net_232),
		.c(_0359_)
	);

	or_ii _1189_ (
		.a(new_net_35),
		.b(new_net_805),
		.c(_0360_)
	);

	and_bb _1190_ (
		.a(new_net_421),
		.b(new_net_42),
		.c(_0361_)
	);

	or_bb _1191_ (
		.a(new_net_775),
		.b(new_net_860),
		.c(_0362_)
	);

	and_ii _1192_ (
		.a(new_net_1029),
		.b(new_net_130),
		.c(_0363_)
	);

	and_bi _1193_ (
		.a(new_net_349),
		.b(new_net_381),
		.c(_0364_)
	);

	inv _1194_ (
		.din(_0364_),
		.dout(_0365_)
	);

	and_bi _1195_ (
		.a(new_net_721),
		.b(new_net_297),
		.c(_0366_)
	);

	or_bi _1196_ (
		.a(new_net_776),
		.b(new_net_861),
		.c(_0367_)
	);

	and_bi _1197_ (
		.a(new_net_131),
		.b(new_net_185),
		.c(_0368_)
	);

	and_bi _1198_ (
		.a(new_net_509),
		.b(new_net_690),
		.c(_0369_)
	);

	and_bi _1199_ (
		.a(new_net_524),
		.b(new_net_562),
		.c(_0370_)
	);

	or_bb _1200_ (
		.a(new_net_626),
		.b(new_net_1337),
		.c(_0371_)
	);

	and_bi _1201_ (
		.a(new_net_132),
		.b(new_net_1030),
		.c(_0372_)
	);

	and_bi _1202_ (
		.a(new_net_913),
		.b(new_net_740),
		.c(_0373_)
	);

	and_ii _1203_ (
		.a(new_net_186),
		.b(new_net_133),
		.c(_0374_)
	);

	and_bi _1204_ (
		.a(new_net_906),
		.b(new_net_817),
		.c(_0375_)
	);

	and_ii _1205_ (
		.a(new_net_143),
		.b(new_net_418),
		.c(_0376_)
	);

	or_bb _1206_ (
		.a(_0376_),
		.b(new_net_691),
		.c(_0377_)
	);

	and_bi _1207_ (
		.a(new_net_503),
		.b(new_net_956),
		.c(_0378_)
	);

	or_bb _1208_ (
		.a(new_net_781),
		.b(new_net_865),
		.c(_0379_)
	);

	or_bb _1209_ (
		.a(_0379_),
		.b(new_net_1338),
		.c(_0380_)
	);

	and_bi _1210_ (
		.a(new_net_541),
		.b(new_net_522),
		.c(_0381_)
	);

	inv _1211_ (
		.din(new_net_162),
		.dout(_0382_)
	);

	inv _1212_ (
		.din(new_net_601),
		.dout(_0383_)
	);

	and_bi _1213_ (
		.a(new_net_971),
		.b(new_net_824),
		.c(_0384_)
	);

	or_bb _1214_ (
		.a(new_net_267),
		.b(new_net_200),
		.c(_0385_)
	);

	or_bb _1215_ (
		.a(_0385_),
		.b(new_net_1339),
		.c(_0386_)
	);

	or_bb _1216_ (
		.a(_0386_),
		.b(_0380_),
		.c(_0387_)
	);

	or_bb _1217_ (
		.a(new_net_1340),
		.b(_0371_),
		.c(_0388_)
	);

	or_bi _1218_ (
		.a(new_net_306),
		.b(new_net_318),
		.c(_0389_)
	);

	and_bi _1219_ (
		.a(new_net_355),
		.b(new_net_506),
		.c(_0390_)
	);

	and_bi _1220_ (
		.a(new_net_675),
		.b(new_net_962),
		.c(_0391_)
	);

	or_bb _1221_ (
		.a(new_net_1341),
		.b(_0390_),
		.c(_0392_)
	);

	and_bi _1222_ (
		.a(new_net_1342),
		.b(_0392_),
		.c(_0393_)
	);

	and_bi _1223_ (
		.a(new_net_460),
		.b(new_net_301),
		.c(_0394_)
	);

	or_bb _1224_ (
		.a(_0394_),
		.b(new_net_154),
		.c(_0395_)
	);

	and_bi _1225_ (
		.a(new_net_615),
		.b(new_net_564),
		.c(_0396_)
	);

	and_bi _1226_ (
		.a(new_net_401),
		.b(new_net_741),
		.c(_0397_)
	);

	and_bi _1227_ (
		.a(new_net_280),
		.b(new_net_441),
		.c(_0398_)
	);

	and_ii _1228_ (
		.a(new_net_469),
		.b(new_net_819),
		.c(_0399_)
	);

	or_bb _1229_ (
		.a(_0399_),
		.b(_0397_),
		.c(_0400_)
	);

	or_bb _1230_ (
		.a(new_net_1343),
		.b(_0396_),
		.c(_0401_)
	);

	or_bb _1231_ (
		.a(_0401_),
		.b(new_net_787),
		.c(_0402_)
	);

	and_bi _1232_ (
		.a(new_net_1344),
		.b(_0402_),
		.c(_0403_)
	);

	and_bi _1233_ (
		.a(_0388_),
		.b(_0403_),
		.c(_0404_)
	);

	and_bi _1234_ (
		.a(new_net_79),
		.b(_0404_),
		.c(_0405_)
	);

	and_bi _1235_ (
		.a(new_net_1012),
		.b(new_net_248),
		.c(_0406_)
	);

	inv _1236_ (
		.din(new_net_342),
		.dout(_0407_)
	);

	or_bb _1237_ (
		.a(new_net_981),
		.b(_0405_),
		.c(_0408_)
	);

	and_bi _1238_ (
		.a(_0357_),
		.b(new_net_1345),
		.c(_0409_)
	);

	or_bb _1239_ (
		.a(new_net_1346),
		.b(_0355_),
		.c(_0410_)
	);

	or_bb _1240_ (
		.a(_0410_),
		.b(new_net_1347),
		.c(new_net_1)
	);

	and_bi _1241_ (
		.a(new_net_71),
		.b(new_net_991),
		.c(_0411_)
	);

	or_bb _1242_ (
		.a(new_net_558),
		.b(new_net_194),
		.c(_0412_)
	);

	or_ii _1243_ (
		.a(new_net_559),
		.b(new_net_195),
		.c(_0413_)
	);

	or_ii _1244_ (
		.a(_0413_),
		.b(_0412_),
		.c(_0414_)
	);

	or_bb _1245_ (
		.a(new_net_725),
		.b(new_net_237),
		.c(_0415_)
	);

	and_ii _1246_ (
		.a(new_net_674),
		.b(new_net_403),
		.c(_0416_)
	);

	and_ii _1247_ (
		.a(new_net_810),
		.b(new_net_823),
		.c(_0417_)
	);

	and_bi _1248_ (
		.a(new_net_319),
		.b(new_net_521),
		.c(_0418_)
	);

	and_bi _1249_ (
		.a(new_net_461),
		.b(new_net_563),
		.c(_0419_)
	);

	or_bb _1250_ (
		.a(_0419_),
		.b(new_net_1348),
		.c(_0420_)
	);

	and_bi _1251_ (
		.a(new_net_357),
		.b(new_net_738),
		.c(_0421_)
	);

	or_bb _1252_ (
		.a(new_net_1349),
		.b(new_net_443),
		.c(_0422_)
	);

	and_bi _1253_ (
		.a(new_net_1350),
		.b(new_net_302),
		.c(_0423_)
	);

	or_bb _1254_ (
		.a(_0423_),
		.b(new_net_1351),
		.c(_0424_)
	);

	or_bi _1255_ (
		.a(new_net_957),
		.b(new_net_614),
		.c(_0425_)
	);

	or_ii _1256_ (
		.a(_0425_),
		.b(new_net_235),
		.c(_0426_)
	);

	or_bb _1257_ (
		.a(new_net_1352),
		.b(_0424_),
		.c(_0427_)
	);

	or_bb _1258_ (
		.a(new_net_1353),
		.b(_0420_),
		.c(_0428_)
	);

	or_bb _1259_ (
		.a(_0428_),
		.b(new_net_1354),
		.c(_0429_)
	);

	and_bi _1260_ (
		.a(new_net_505),
		.b(new_net_571),
		.c(_0430_)
	);

	and_bi _1261_ (
		.a(new_net_125),
		.b(new_net_370),
		.c(_0431_)
	);

	and_bi _1262_ (
		.a(new_net_908),
		.b(new_net_964),
		.c(_0432_)
	);

	and_bi _1263_ (
		.a(new_net_909),
		.b(new_net_511),
		.c(_0433_)
	);

	or_bb _1264_ (
		.a(_0433_),
		.b(new_net_547),
		.c(_0434_)
	);

	and_bi _1265_ (
		.a(new_net_973),
		.b(new_net_731),
		.c(_0435_)
	);

	and_bi _1266_ (
		.a(new_net_189),
		.b(new_net_818),
		.c(_0436_)
	);

	or_bb _1267_ (
		.a(new_net_808),
		.b(new_net_1355),
		.c(_0437_)
	);

	or_bb _1268_ (
		.a(_0437_),
		.b(_0434_),
		.c(_0438_)
	);

	and_bi _1269_ (
		.a(new_net_56),
		.b(new_net_537),
		.c(_0439_)
	);

	and_ii _1270_ (
		.a(new_net_888),
		.b(new_net_307),
		.c(_0440_)
	);

	and_bi _1271_ (
		.a(new_net_797),
		.b(new_net_825),
		.c(_0441_)
	);

	or_bb _1272_ (
		.a(_0441_),
		.b(new_net_167),
		.c(_0442_)
	);

	or_bb _1273_ (
		.a(new_net_694),
		.b(new_net_1356),
		.c(_0443_)
	);

	or_bb _1274_ (
		.a(_0443_),
		.b(_0438_),
		.c(_0444_)
	);

	and_bi _1275_ (
		.a(_0431_),
		.b(new_net_1357),
		.c(_0445_)
	);

	and_bi _1276_ (
		.a(_0429_),
		.b(_0445_),
		.c(_0446_)
	);

	and_bi _1277_ (
		.a(new_net_75),
		.b(_0446_),
		.c(_0447_)
	);

	or_bb _1278_ (
		.a(_0447_),
		.b(new_net_985),
		.c(_0448_)
	);

	and_bi _1279_ (
		.a(_0415_),
		.b(new_net_1358),
		.c(_0449_)
	);

	and_bi _1280_ (
		.a(new_net_452),
		.b(new_net_587),
		.c(_0450_)
	);

	and_bi _1281_ (
		.a(new_net_582),
		.b(new_net_586),
		.c(_0451_)
	);

	and_bi _1282_ (
		.a(new_net_23),
		.b(_0451_),
		.c(_0452_)
	);

	and_bi _1283_ (
		.a(new_net_1359),
		.b(new_net_554),
		.c(_0453_)
	);

	or_bb _1284_ (
		.a(_0453_),
		.b(new_net_923),
		.c(_0454_)
	);

	and_bb _1285_ (
		.a(new_net_990),
		.b(new_net_377),
		.c(_0455_)
	);

	and_ii _1286_ (
		.a(new_net_1360),
		.b(new_net_648),
		.c(_0456_)
	);

	or_bi _1287_ (
		.a(new_net_1003),
		.b(new_net_726),
		.c(_0457_)
	);

	and_bi _1288_ (
		.a(new_net_1004),
		.b(new_net_727),
		.c(_0458_)
	);

	and_bi _1289_ (
		.a(_0457_),
		.b(_0458_),
		.c(_0459_)
	);

	or_bi _1290_ (
		.a(new_net_326),
		.b(new_net_697),
		.c(_0460_)
	);

	and_bi _1291_ (
		.a(new_net_325),
		.b(new_net_698),
		.c(_0461_)
	);

	and_bi _1292_ (
		.a(_0460_),
		.b(_0461_),
		.c(_0462_)
	);

	and_bi _1293_ (
		.a(_0454_),
		.b(new_net_1361),
		.c(_0463_)
	);

	or_bb _1294_ (
		.a(_0463_),
		.b(new_net_1362),
		.c(new_net_0)
	);

	or_bb _1295_ (
		.a(new_net_374),
		.b(new_net_900),
		.c(_0464_)
	);

	or_bb _1296_ (
		.a(new_net_239),
		.b(new_net_644),
		.c(_0465_)
	);

	and_bi _1297_ (
		.a(new_net_462),
		.b(new_net_730),
		.c(_0466_)
	);

	and_bi _1298_ (
		.a(new_net_801),
		.b(new_net_963),
		.c(_0467_)
	);

	and_bi _1299_ (
		.a(new_net_444),
		.b(new_net_512),
		.c(_0468_)
	);

	or_bb _1300_ (
		.a(_0468_),
		.b(new_net_1363),
		.c(_0469_)
	);

	or_bb _1301_ (
		.a(_0469_),
		.b(new_net_1364),
		.c(_0470_)
	);

	and_bi _1302_ (
		.a(new_net_720),
		.b(new_net_570),
		.c(_0471_)
	);

	and_bi _1303_ (
		.a(new_net_671),
		.b(new_net_310),
		.c(_0472_)
	);

	or_bb _1304_ (
		.a(_0472_),
		.b(new_net_180),
		.c(_0473_)
	);

	and_bi _1305_ (
		.a(new_net_402),
		.b(new_net_303),
		.c(_0474_)
	);

	or_bi _1306_ (
		.a(new_net_617),
		.b(new_net_266),
		.c(_0475_)
	);

	and_bi _1307_ (
		.a(new_net_1365),
		.b(new_net_826),
		.c(_0476_)
	);

	or_bb _1308_ (
		.a(new_net_1366),
		.b(_0474_),
		.c(_0477_)
	);

	or_bb _1309_ (
		.a(new_net_1367),
		.b(new_net_487),
		.c(_0478_)
	);

	or_bb _1310_ (
		.a(_0478_),
		.b(_0471_),
		.c(_0479_)
	);

	or_bb _1311_ (
		.a(_0479_),
		.b(new_net_1368),
		.c(_0480_)
	);

	and_bi _1312_ (
		.a(new_net_191),
		.b(new_net_965),
		.c(_0481_)
	);

	or_bi _1313_ (
		.a(new_net_739),
		.b(new_net_383),
		.c(_0482_)
	);

	and_bi _1314_ (
		.a(_0482_),
		.b(new_net_881),
		.c(_0483_)
	);

	and_bi _1315_ (
		.a(new_net_634),
		.b(new_net_513),
		.c(_0484_)
	);

	and_ii _1316_ (
		.a(new_net_889),
		.b(new_net_828),
		.c(_0485_)
	);

	or_bb _1317_ (
		.a(new_net_1369),
		.b(_0484_),
		.c(_0486_)
	);

	and_bi _1318_ (
		.a(new_net_1370),
		.b(_0486_),
		.c(_0487_)
	);

	and_bi _1319_ (
		.a(new_net_974),
		.b(new_net_565),
		.c(_0488_)
	);

	and_bi _1320_ (
		.a(new_net_850),
		.b(new_net_755),
		.c(_0489_)
	);

	and_ii _1321_ (
		.a(new_net_295),
		.b(new_net_298),
		.c(_0490_)
	);

	or_bb _1322_ (
		.a(_0490_),
		.b(new_net_202),
		.c(_0491_)
	);

	or_bb _1323_ (
		.a(new_net_1371),
		.b(_0488_),
		.c(_0492_)
	);

	and_bi _1324_ (
		.a(new_net_1372),
		.b(_0492_),
		.c(_0493_)
	);

	and_bi _1325_ (
		.a(_0480_),
		.b(_0493_),
		.c(_0494_)
	);

	and_bi _1326_ (
		.a(new_net_81),
		.b(_0494_),
		.c(_0495_)
	);

	or_bb _1327_ (
		.a(_0495_),
		.b(new_net_983),
		.c(_0496_)
	);

	and_bi _1328_ (
		.a(_0465_),
		.b(new_net_1373),
		.c(_0497_)
	);

	inv _1329_ (
		.din(new_net_994),
		.dout(_0498_)
	);

	and_bi _1330_ (
		.a(new_net_440),
		.b(new_net_1374),
		.c(_0499_)
	);

	and_bb _1331_ (
		.a(new_net_1022),
		.b(new_net_323),
		.c(_0500_)
	);

	and_ii _1332_ (
		.a(new_net_1375),
		.b(new_net_119),
		.c(_0501_)
	);

	or_bi _1333_ (
		.a(new_net_456),
		.b(new_net_867),
		.c(_0502_)
	);

	and_bi _1334_ (
		.a(new_net_457),
		.b(new_net_868),
		.c(_0503_)
	);

	or_bb _1335_ (
		.a(_0503_),
		.b(new_net_344),
		.c(_0504_)
	);

	and_bi _1336_ (
		.a(new_net_1376),
		.b(_0504_),
		.c(_0505_)
	);

	or_bb _1337_ (
		.a(_0505_),
		.b(new_net_1377),
		.c(new_net_3)
	);

	and_bi _1338_ (
		.a(new_net_778),
		.b(new_net_555),
		.c(_0506_)
	);

	or_bb _1339_ (
		.a(new_net_238),
		.b(new_net_709),
		.c(_0507_)
	);

	and_bi _1340_ (
		.a(new_net_540),
		.b(new_net_735),
		.c(_0508_)
	);

	and_bi _1341_ (
		.a(new_net_382),
		.b(new_net_514),
		.c(_0509_)
	);

	or_bb _1342_ (
		.a(_0509_),
		.b(new_net_1378),
		.c(_0510_)
	);

	or_ii _1343_ (
		.a(new_net_846),
		.b(new_net_895),
		.c(_0511_)
	);

	and_bi _1344_ (
		.a(new_net_1379),
		.b(new_net_820),
		.c(_0512_)
	);

	and_bi _1345_ (
		.a(new_net_526),
		.b(new_net_958),
		.c(_0513_)
	);

	or_bb _1346_ (
		.a(new_net_779),
		.b(_0512_),
		.c(_0514_)
	);

	or_bb _1347_ (
		.a(new_net_1380),
		.b(_0510_),
		.c(_0515_)
	);

	and_bi _1348_ (
		.a(new_net_192),
		.b(new_net_572),
		.c(_0516_)
	);

	and_bi _1349_ (
		.a(new_net_594),
		.b(new_net_635),
		.c(_0517_)
	);

	and_ii _1350_ (
		.a(new_net_746),
		.b(new_net_312),
		.c(_0518_)
	);

	or_bb _1351_ (
		.a(_0518_),
		.b(new_net_196),
		.c(_0519_)
	);

	or_bb _1352_ (
		.a(new_net_1381),
		.b(_0516_),
		.c(_0520_)
	);

	or_bb _1353_ (
		.a(_0520_),
		.b(new_net_1382),
		.c(_0521_)
	);

	or_bi _1354_ (
		.a(new_net_308),
		.b(new_net_356),
		.c(_0522_)
	);

	and_bi _1355_ (
		.a(new_net_442),
		.b(new_net_732),
		.c(_0523_)
	);

	and_bi _1356_ (
		.a(new_net_618),
		.b(new_net_309),
		.c(_0524_)
	);

	or_bb _1357_ (
		.a(new_net_933),
		.b(new_net_1383),
		.c(_0525_)
	);

	and_bi _1358_ (
		.a(new_net_1384),
		.b(_0525_),
		.c(_0526_)
	);

	and_ii _1359_ (
		.a(new_net_811),
		.b(new_net_507),
		.c(_0527_)
	);

	or_bb _1360_ (
		.a(_0527_),
		.b(new_net_1044),
		.c(_0528_)
	);

	and_bi _1361_ (
		.a(new_net_716),
		.b(new_net_959),
		.c(_0529_)
	);

	and_bi _1362_ (
		.a(new_net_464),
		.b(new_net_829),
		.c(_0530_)
	);

	or_bb _1363_ (
		.a(_0530_),
		.b(new_net_1385),
		.c(_0531_)
	);

	or_bb _1364_ (
		.a(new_net_1386),
		.b(_0528_),
		.c(_0532_)
	);

	or_bb _1365_ (
		.a(_0532_),
		.b(new_net_695),
		.c(_0533_)
	);

	and_bi _1366_ (
		.a(_0526_),
		.b(_0533_),
		.c(_0534_)
	);

	and_bi _1367_ (
		.a(_0521_),
		.b(new_net_1387),
		.c(_0535_)
	);

	and_bi _1368_ (
		.a(new_net_80),
		.b(_0535_),
		.c(_0536_)
	);

	or_bb _1369_ (
		.a(_0536_),
		.b(new_net_982),
		.c(_0537_)
	);

	and_bi _1370_ (
		.a(_0507_),
		.b(new_net_1388),
		.c(_0538_)
	);

	and_bi _1371_ (
		.a(new_net_922),
		.b(new_net_453),
		.c(_0539_)
	);

	or_bb _1372_ (
		.a(_0539_),
		.b(new_net_1389),
		.c(_0540_)
	);

	or_bb _1373_ (
		.a(new_net_1390),
		.b(_0506_),
		.c(new_net_2)
	);

	or_bb _1374_ (
		.a(new_net_873),
		.b(new_net_106),
		.c(_0541_)
	);

	or_bb _1375_ (
		.a(new_net_475),
		.b(new_net_109),
		.c(_0542_)
	);

	and_bi _1376_ (
		.a(new_net_831),
		.b(new_net_918),
		.c(_0543_)
	);

	and_bi _1377_ (
		.a(new_net_917),
		.b(new_net_832),
		.c(_0544_)
	);

	or_bb _1378_ (
		.a(_0544_),
		.b(_0543_),
		.c(_0545_)
	);

	and_ii _1379_ (
		.a(new_net_476),
		.b(new_net_366),
		.c(_0546_)
	);

	or_bb _1380_ (
		.a(new_net_497),
		.b(new_net_551),
		.c(_0547_)
	);

	and_bb _1381_ (
		.a(new_net_498),
		.b(new_net_550),
		.c(_0548_)
	);

	and_bi _1382_ (
		.a(_0547_),
		.b(_0548_),
		.c(_0549_)
	);

	or_ii _1383_ (
		.a(new_net_620),
		.b(new_net_995),
		.c(_0550_)
	);

	and_bi _1384_ (
		.a(new_net_953),
		.b(_0550_),
		.c(new_net_4)
	);

	and_ii _1385_ (
		.a(new_net_477),
		.b(new_net_51),
		.c(_0551_)
	);

	or_bi _1386_ (
		.a(new_net_228),
		.b(new_net_858),
		.c(_0552_)
	);

	and_bi _1387_ (
		.a(new_net_229),
		.b(new_net_857),
		.c(_0553_)
	);

	or_bi _1388_ (
		.a(_0553_),
		.b(_0552_),
		.c(_0554_)
	);

	and_bi _1389_ (
		.a(new_net_478),
		.b(new_net_887),
		.c(_0555_)
	);

	or_bi _1390_ (
		.a(new_net_1041),
		.b(new_net_955),
		.c(_0556_)
	);

	and_bi _1391_ (
		.a(new_net_479),
		.b(new_net_768),
		.c(_0557_)
	);

	and_bi _1392_ (
		.a(new_net_445),
		.b(new_net_1391),
		.c(_0558_)
	);

	and_bi _1393_ (
		.a(new_net_362),
		.b(new_net_753),
		.c(_0559_)
	);

	and_bi _1394_ (
		.a(new_net_754),
		.b(new_net_364),
		.c(_0560_)
	);

	and_ii _1395_ (
		.a(new_net_1392),
		.b(new_net_607),
		.c(_0561_)
	);

	and_bi _1396_ (
		.a(new_net_433),
		.b(new_net_979),
		.c(_0562_)
	);

	and_bi _1397_ (
		.a(new_net_980),
		.b(new_net_434),
		.c(_0563_)
	);

	or_bb _1398_ (
		.a(new_net_928),
		.b(new_net_1393),
		.c(_0564_)
	);

	and_bi _1399_ (
		.a(new_net_993),
		.b(new_net_623),
		.c(_0565_)
	);

	inv _1400_ (
		.din(new_net_368),
		.dout(_0566_)
	);

	and_bb _1401_ (
		.a(new_net_1042),
		.b(new_net_916),
		.c(_0567_)
	);

	or_bi _1402_ (
		.a(new_net_1394),
		.b(new_net_446),
		.c(_0568_)
	);

	or_ii _1403_ (
		.a(new_net_838),
		.b(new_net_935),
		.c(_0569_)
	);

	and_bi _1404_ (
		.a(new_net_369),
		.b(new_net_839),
		.c(_0570_)
	);

	and_bi _1405_ (
		.a(_0569_),
		.b(_0570_),
		.c(_0571_)
	);

	or_bb _1406_ (
		.a(new_net_214),
		.b(new_net_1026),
		.c(_0572_)
	);

	or_ii _1407_ (
		.a(new_net_255),
		.b(new_net_19),
		.c(_0573_)
	);

	and_ii _1408_ (
		.a(new_net_1395),
		.b(new_net_122),
		.c(_0574_)
	);

	or_bb _1409_ (
		.a(new_net_655),
		.b(new_net_493),
		.c(_0575_)
	);

	or_bb _1410_ (
		.a(new_net_222),
		.b(new_net_363),
		.c(_0576_)
	);

	and_bi _1411_ (
		.a(new_net_616),
		.b(new_net_515),
		.c(_0577_)
	);

	and_bi _1412_ (
		.a(new_net_803),
		.b(new_net_313),
		.c(_0578_)
	);

	or_ii _1413_ (
		.a(new_net_281),
		.b(new_net_57),
		.c(_0579_)
	);

	and_bi _1414_ (
		.a(new_net_1396),
		.b(new_net_821),
		.c(_0580_)
	);

	or_bb _1415_ (
		.a(new_net_1397),
		.b(_0578_),
		.c(_0581_)
	);

	or_bb _1416_ (
		.a(_0581_),
		.b(new_net_1398),
		.c(_0582_)
	);

	and_bi _1417_ (
		.a(new_net_904),
		.b(new_net_566),
		.c(_0583_)
	);

	and_bi _1418_ (
		.a(new_net_676),
		.b(new_net_736),
		.c(_0584_)
	);

	or_bb _1419_ (
		.a(_0584_),
		.b(new_net_782),
		.c(_0585_)
	);

	or_bb _1420_ (
		.a(new_net_1399),
		.b(new_net_788),
		.c(_0586_)
	);

	or_bb _1421_ (
		.a(_0586_),
		.b(_0583_),
		.c(_0587_)
	);

	or_bb _1422_ (
		.a(_0587_),
		.b(new_net_1400),
		.c(_0588_)
	);

	or_bi _1423_ (
		.a(new_net_733),
		.b(new_net_757),
		.c(_0589_)
	);

	or_bb _1424_ (
		.a(new_net_851),
		.b(new_net_386),
		.c(_0590_)
	);

	and_bi _1425_ (
		.a(new_net_1401),
		.b(new_net_299),
		.c(_0591_)
	);

	and_bi _1426_ (
		.a(new_net_1402),
		.b(_0591_),
		.c(_0592_)
	);

	and_bi _1427_ (
		.a(new_net_62),
		.b(new_net_516),
		.c(_0593_)
	);

	and_bi _1428_ (
		.a(new_net_912),
		.b(new_net_966),
		.c(_0594_)
	);

	or_bb _1429_ (
		.a(new_net_1403),
		.b(_0593_),
		.c(_0595_)
	);

	and_bi _1430_ (
		.a(_0592_),
		.b(_0595_),
		.c(_0596_)
	);

	and_bi _1431_ (
		.a(new_net_538),
		.b(new_net_567),
		.c(_0597_)
	);

	and_ii _1432_ (
		.a(new_net_747),
		.b(new_net_830),
		.c(_0598_)
	);

	or_bb _1433_ (
		.a(_0598_),
		.b(new_net_197),
		.c(_0599_)
	);

	or_bb _1434_ (
		.a(new_net_1404),
		.b(_0597_),
		.c(_0600_)
	);

	and_bi _1435_ (
		.a(new_net_1405),
		.b(_0600_),
		.c(_0601_)
	);

	and_bi _1436_ (
		.a(_0588_),
		.b(_0601_),
		.c(_0602_)
	);

	and_bi _1437_ (
		.a(new_net_76),
		.b(_0602_),
		.c(_0603_)
	);

	or_bb _1438_ (
		.a(_0603_),
		.b(new_net_986),
		.c(_0604_)
	);

	and_bi _1439_ (
		.a(_0576_),
		.b(new_net_1406),
		.c(_0605_)
	);

	and_bi _1440_ (
		.a(new_net_22),
		.b(new_net_257),
		.c(_0606_)
	);

	and_ii _1441_ (
		.a(_0606_),
		.b(new_net_921),
		.c(_0607_)
	);

	and_bi _1442_ (
		.a(new_net_123),
		.b(new_net_1407),
		.c(_0608_)
	);

	or_bb _1443_ (
		.a(_0608_),
		.b(new_net_1408),
		.c(_0609_)
	);

	or_bb _1444_ (
		.a(_0609_),
		.b(new_net_1409),
		.c(new_net_6)
	);

	and_bb _1445_ (
		.a(new_net_215),
		.b(new_net_1023),
		.c(_0610_)
	);

	or_bi _1446_ (
		.a(_0610_),
		.b(new_net_24),
		.c(_0611_)
	);

	and_bi _1447_ (
		.a(new_net_1024),
		.b(new_net_124),
		.c(_0612_)
	);

	and_ii _1448_ (
		.a(_0612_),
		.b(new_net_27),
		.c(_0613_)
	);

	or_bb _1449_ (
		.a(_0613_),
		.b(new_net_920),
		.c(_0614_)
	);

	and_bi _1450_ (
		.a(new_net_706),
		.b(new_net_629),
		.c(_0615_)
	);

	or_bb _1451_ (
		.a(new_net_1410),
		.b(new_net_608),
		.c(_0616_)
	);

	and_bi _1452_ (
		.a(new_net_835),
		.b(new_net_482),
		.c(_0617_)
	);

	inv _1453_ (
		.din(_0617_),
		.dout(_0618_)
	);

	and_bi _1454_ (
		.a(new_net_431),
		.b(new_net_528),
		.c(_0619_)
	);

	and_bi _1455_ (
		.a(new_net_529),
		.b(new_net_432),
		.c(_0621_)
	);

	and_ii _1456_ (
		.a(_0621_),
		.b(_0619_),
		.c(_0622_)
	);

	or_bb _1457_ (
		.a(new_net_649),
		.b(new_net_338),
		.c(_0623_)
	);

	and_bb _1458_ (
		.a(new_net_650),
		.b(new_net_339),
		.c(_0624_)
	);

	and_bi _1459_ (
		.a(_0623_),
		.b(_0624_),
		.c(_0625_)
	);

	or_ii _1460_ (
		.a(new_net_345),
		.b(new_net_929),
		.c(_0626_)
	);

	or_bb _1461_ (
		.a(new_net_346),
		.b(new_net_930),
		.c(_0627_)
	);

	and_bb _1462_ (
		.a(_0627_),
		.b(_0626_),
		.c(_0628_)
	);

	and_bi _1463_ (
		.a(_0614_),
		.b(new_net_1411),
		.c(_0629_)
	);

	or_bi _1464_ (
		.a(new_net_223),
		.b(new_net_651),
		.c(_0630_)
	);

	and_ii _1465_ (
		.a(new_net_470),
		.b(new_net_311),
		.c(_0632_)
	);

	and_bi _1466_ (
		.a(new_net_619),
		.b(new_net_742),
		.c(_0633_)
	);

	and_bi _1467_ (
		.a(new_net_463),
		.b(new_net_508),
		.c(_0634_)
	);

	or_bb _1468_ (
		.a(_0634_),
		.b(new_net_1412),
		.c(_0635_)
	);

	or_bb _1469_ (
		.a(_0635_),
		.b(new_net_1413),
		.c(_0636_)
	);

	or_bi _1470_ (
		.a(new_net_677),
		.b(new_net_898),
		.c(_0637_)
	);

	and_bi _1471_ (
		.a(new_net_1414),
		.b(new_net_815),
		.c(_0638_)
	);

	or_bb _1472_ (
		.a(new_net_1415),
		.b(_0636_),
		.c(_0639_)
	);

	and_bi _1473_ (
		.a(new_net_798),
		.b(new_net_568),
		.c(_0640_)
	);

	or_bb _1474_ (
		.a(_0640_),
		.b(new_net_548),
		.c(_0641_)
	);

	or_bb _1475_ (
		.a(_0641_),
		.b(new_net_171),
		.c(_0642_)
	);

	or_bb _1476_ (
		.a(_0642_),
		.b(new_net_1416),
		.c(_0643_)
	);

	and_ii _1477_ (
		.a(new_net_539),
		.b(new_net_64),
		.c(_0644_)
	);

	or_bb _1478_ (
		.a(new_net_840),
		.b(new_net_314),
		.c(_0645_)
	);

	and_bi _1479_ (
		.a(new_net_722),
		.b(new_net_816),
		.c(_0646_)
	);

	and_bi _1480_ (
		.a(_0645_),
		.b(new_net_1417),
		.c(_0647_)
	);

	and_bi _1481_ (
		.a(new_net_756),
		.b(new_net_517),
		.c(_0648_)
	);

	and_bi _1482_ (
		.a(new_net_636),
		.b(new_net_743),
		.c(_0649_)
	);

	or_bb _1483_ (
		.a(new_net_1418),
		.b(_0648_),
		.c(_0650_)
	);

	and_bi _1484_ (
		.a(new_net_914),
		.b(new_net_573),
		.c(_0651_)
	);

	and_bi _1485_ (
		.a(new_net_972),
		.b(new_net_960),
		.c(_0653_)
	);

	or_bb _1486_ (
		.a(_0653_),
		.b(new_net_201),
		.c(_0654_)
	);

	or_bb _1487_ (
		.a(new_net_1419),
		.b(_0651_),
		.c(_0655_)
	);

	or_bb _1488_ (
		.a(_0655_),
		.b(new_net_1420),
		.c(_0656_)
	);

	and_bi _1489_ (
		.a(new_net_1421),
		.b(_0656_),
		.c(_0657_)
	);

	and_bi _1490_ (
		.a(_0643_),
		.b(_0657_),
		.c(_0658_)
	);

	and_bi _1491_ (
		.a(new_net_77),
		.b(_0658_),
		.c(_0659_)
	);

	or_bb _1492_ (
		.a(_0659_),
		.b(new_net_987),
		.c(_0660_)
	);

	and_bi _1493_ (
		.a(_0630_),
		.b(new_net_1422),
		.c(_0661_)
	);

	or_bb _1494_ (
		.a(new_net_1423),
		.b(_0629_),
		.c(new_net_5)
	);

	or_bb _1495_ (
		.a(new_net_500),
		.b(new_net_532),
		.c(_0663_)
	);

	or_bi _1496_ (
		.a(new_net_225),
		.b(new_net_621),
		.c(_0664_)
	);

	and_ii _1497_ (
		.a(new_net_841),
		.b(new_net_827),
		.c(_0665_)
	);

	and_bi _1498_ (
		.a(new_net_637),
		.b(new_net_43),
		.c(_0666_)
	);

	or_bb _1499_ (
		.a(new_net_1424),
		.b(new_net_198),
		.c(_0667_)
	);

	or_bb _1500_ (
		.a(new_net_1425),
		.b(_0665_),
		.c(_0668_)
	);

	and_bi _1501_ (
		.a(new_net_384),
		.b(new_net_961),
		.c(_0669_)
	);

	and_bi _1502_ (
		.a(new_net_853),
		.b(new_net_744),
		.c(_0670_)
	);

	or_bb _1503_ (
		.a(_0670_),
		.b(new_net_1426),
		.c(_0671_)
	);

	and_ii _1504_ (
		.a(new_net_638),
		.b(new_net_1427),
		.c(_0672_)
	);

	and_ii _1505_ (
		.a(new_net_783),
		.b(new_net_518),
		.c(_0674_)
	);

	or_bb _1506_ (
		.a(new_net_1428),
		.b(new_net_758),
		.c(_0675_)
	);

	and_bi _1507_ (
		.a(new_net_1429),
		.b(new_net_300),
		.c(_0676_)
	);

	or_bb _1508_ (
		.a(_0676_),
		.b(_0674_),
		.c(_0677_)
	);

	or_bb _1509_ (
		.a(_0677_),
		.b(new_net_1430),
		.c(_0678_)
	);

	or_bb _1510_ (
		.a(_0678_),
		.b(new_net_1431),
		.c(_0679_)
	);

	and_ii _1511_ (
		.a(new_net_268),
		.b(new_net_627),
		.c(_0680_)
	);

	and_bi _1512_ (
		.a(new_net_719),
		.b(new_net_510),
		.c(_0681_)
	);

	or_bb _1513_ (
		.a(_0681_),
		.b(new_net_866),
		.c(_0682_)
	);

	and_bi _1514_ (
		.a(new_net_504),
		.b(new_net_315),
		.c(_0683_)
	);

	and_bi _1515_ (
		.a(new_net_799),
		.b(new_net_734),
		.c(_0685_)
	);

	or_bb _1516_ (
		.a(new_net_1432),
		.b(_0683_),
		.c(_0686_)
	);

	or_bb _1517_ (
		.a(_0686_),
		.b(_0682_),
		.c(_0687_)
	);

	or_bb _1518_ (
		.a(new_net_882),
		.b(new_net_488),
		.c(_0688_)
	);

	or_bb _1519_ (
		.a(_0688_),
		.b(new_net_1433),
		.c(_0689_)
	);

	and_bi _1520_ (
		.a(_0680_),
		.b(new_net_1434),
		.c(_0690_)
	);

	and_bi _1521_ (
		.a(new_net_1435),
		.b(_0690_),
		.c(_0691_)
	);

	and_bi _1522_ (
		.a(new_net_82),
		.b(_0691_),
		.c(_0692_)
	);

	or_bb _1523_ (
		.a(_0692_),
		.b(new_net_984),
		.c(_0693_)
	);

	and_bi _1524_ (
		.a(_0664_),
		.b(new_net_1436),
		.c(_0694_)
	);

	and_bi _1525_ (
		.a(new_net_622),
		.b(new_net_992),
		.c(_0696_)
	);

	or_bb _1526_ (
		.a(_0696_),
		.b(new_net_343),
		.c(_0697_)
	);

	and_bi _1527_ (
		.a(new_net_936),
		.b(new_net_1437),
		.c(_0698_)
	);

	or_bb _1528_ (
		.a(_0698_),
		.b(new_net_1438),
		.c(new_net_8)
	);

	and_bi _1529_ (
		.a(new_net_256),
		.b(new_net_28),
		.c(_0699_)
	);

	and_bi _1530_ (
		.a(new_net_924),
		.b(new_net_216),
		.c(_0700_)
	);

	or_bb _1531_ (
		.a(new_net_224),
		.b(new_net_954),
		.c(_0701_)
	);

	and_bi _1532_ (
		.a(new_net_543),
		.b(new_net_967),
		.c(_0702_)
	);

	and_bi _1533_ (
		.a(new_net_852),
		.b(new_net_519),
		.c(_0703_)
	);

	or_bb _1534_ (
		.a(_0703_),
		.b(new_net_1439),
		.c(_0704_)
	);

	and_ii _1535_ (
		.a(new_net_784),
		.b(new_net_304),
		.c(_0706_)
	);

	and_bi _1536_ (
		.a(new_net_63),
		.b(new_net_737),
		.c(_0707_)
	);

	or_bb _1537_ (
		.a(new_net_1440),
		.b(_0706_),
		.c(_0708_)
	);

	or_bb _1538_ (
		.a(_0708_),
		.b(_0704_),
		.c(_0709_)
	);

	and_bi _1539_ (
		.a(new_net_385),
		.b(new_net_569),
		.c(_0710_)
	);

	and_ii _1540_ (
		.a(new_net_296),
		.b(new_net_822),
		.c(_0711_)
	);

	or_bb _1541_ (
		.a(_0711_),
		.b(new_net_199),
		.c(_0712_)
	);

	or_bb _1542_ (
		.a(new_net_1441),
		.b(_0710_),
		.c(_0713_)
	);

	or_bb _1543_ (
		.a(_0713_),
		.b(new_net_1442),
		.c(_0714_)
	);

	or_bb _1544_ (
		.a(new_net_745),
		.b(new_net_288),
		.c(_0715_)
	);

	and_bi _1545_ (
		.a(new_net_672),
		.b(new_net_520),
		.c(_0717_)
	);

	and_bi _1546_ (
		.a(new_net_1443),
		.b(_0717_),
		.c(_0718_)
	);

	and_bi _1547_ (
		.a(new_net_905),
		.b(new_net_305),
		.c(_0719_)
	);

	or_bb _1548_ (
		.a(_0719_),
		.b(new_net_809),
		.c(_0720_)
	);

	and_bi _1549_ (
		.a(_0718_),
		.b(_0720_),
		.c(_0721_)
	);

	or_bb _1550_ (
		.a(new_net_934),
		.b(new_net_780),
		.c(_0722_)
	);

	or_bb _1551_ (
		.a(_0722_),
		.b(new_net_696),
		.c(_0723_)
	);

	or_bb _1552_ (
		.a(new_net_1444),
		.b(new_net_371),
		.c(_0724_)
	);

	and_bi _1553_ (
		.a(new_net_1445),
		.b(_0724_),
		.c(_0725_)
	);

	and_bi _1554_ (
		.a(new_net_1446),
		.b(_0725_),
		.c(_0726_)
	);

	and_bi _1555_ (
		.a(new_net_78),
		.b(_0726_),
		.c(_0728_)
	);

	or_bb _1556_ (
		.a(_0728_),
		.b(new_net_988),
		.c(_0729_)
	);

	and_bi _1557_ (
		.a(_0701_),
		.b(new_net_1447),
		.c(_0730_)
	);

	or_bb _1558_ (
		.a(new_net_1448),
		.b(_0700_),
		.c(_0731_)
	);

	or_bb _1559_ (
		.a(new_net_1449),
		.b(_0699_),
		.c(new_net_7)
	);

	or_bb _1560_ (
		.a(new_net_751),
		.b(new_net_976),
		.c(_0732_)
	);

	or_bb _1561_ (
		.a(new_net_854),
		.b(new_net_678),
		.c(_0733_)
	);

	or_bb _1562_ (
		.a(new_net_1450),
		.b(new_net_748),
		.c(_0734_)
	);

	and_ii _1563_ (
		.a(_0734_),
		.b(new_net_876),
		.c(_0735_)
	);

	inv _1564_ (
		.din(new_net_997),
		.dout(new_net_1479)
	);

	and_bi _1565_ (
		.a(new_net_45),
		.b(new_net_877),
		.c(_0737_)
	);

	or_bi _1566_ (
		.a(new_net_998),
		.b(new_net_113),
		.c(_0738_)
	);

	or_bb _1567_ (
		.a(_0738_),
		.b(new_net_1451),
		.c(new_net_1473)
	);

	and_bb _1568_ (
		.a(new_net_373),
		.b(new_net_901),
		.c(_0739_)
	);

	and_bi _1569_ (
		.a(new_net_878),
		.b(new_net_1452),
		.c(_0740_)
	);

	and_bb _1570_ (
		.a(new_net_872),
		.b(new_net_107),
		.c(_0741_)
	);

	or_bi _1571_ (
		.a(new_net_1453),
		.b(new_net_749),
		.c(_0742_)
	);

	and_bb _1572_ (
		.a(new_net_752),
		.b(new_net_977),
		.c(_0743_)
	);

	or_bi _1573_ (
		.a(new_net_1454),
		.b(new_net_855),
		.c(_0744_)
	);

	and_bb _1574_ (
		.a(new_net_501),
		.b(new_net_531),
		.c(_0745_)
	);

	and_bi _1575_ (
		.a(new_net_679),
		.b(new_net_1455),
		.c(_0747_)
	);

	and_ii _1576_ (
		.a(new_net_556),
		.b(new_net_425),
		.c(_0748_)
	);

	and_bb _1577_ (
		.a(new_net_557),
		.b(new_net_426),
		.c(_0749_)
	);

	or_bb _1578_ (
		.a(_0749_),
		.b(_0748_),
		.c(_0750_)
	);

	or_bb _1579_ (
		.a(new_net_728),
		.b(new_net_65),
		.c(_0751_)
	);

	and_bb _1580_ (
		.a(new_net_729),
		.b(new_net_66),
		.c(_0752_)
	);

	and_bi _1581_ (
		.a(_0751_),
		.b(_0752_),
		.c(_0753_)
	);

	or_bb _1582_ (
		.a(new_net_701),
		.b(new_net_639),
		.c(_0754_)
	);

	and_bb _1583_ (
		.a(new_net_703),
		.b(new_net_642),
		.c(_0755_)
	);

	and_bi _1584_ (
		.a(_0754_),
		.b(_0755_),
		.c(new_net_1469)
	);

	and_bi _1585_ (
		.a(new_net_949),
		.b(new_net_69),
		.c(new_net_1467)
	);

	and_bi _1586_ (
		.a(new_net_970),
		.b(new_net_359),
		.c(new_net_1471)
	);

	and_bi _1587_ (
		.a(new_net_184),
		.b(new_net_1011),
		.c(_0757_)
	);

	and_bi _1588_ (
		.a(new_net_1028),
		.b(new_net_667),
		.c(_0758_)
	);

	or_bb _1589_ (
		.a(_0758_),
		.b(new_net_1456),
		.c(new_net_1483)
	);

	or_ii _1590_ (
		.a(new_net_1008),
		.b(new_net_969),
		.c(_0759_)
	);

	and_bi _1591_ (
		.a(new_net_1014),
		.b(new_net_1009),
		.c(_0760_)
	);

	and_bi _1592_ (
		.a(_0759_),
		.b(_0760_),
		.c(_0761_)
	);

	and_bi _1593_ (
		.a(new_net_942),
		.b(new_net_1457),
		.c(_0762_)
	);

	and_bi _1594_ (
		.a(new_net_545),
		.b(new_net_1006),
		.c(_0763_)
	);

	and_bi _1595_ (
		.a(new_net_1005),
		.b(new_net_546),
		.c(_0765_)
	);

	and_ii _1596_ (
		.a(_0765_),
		.b(_0763_),
		.c(_0766_)
	);

	or_ii _1597_ (
		.a(new_net_765),
		.b(new_net_836),
		.c(_0767_)
	);

	or_bb _1598_ (
		.a(new_net_766),
		.b(new_net_837),
		.c(_0768_)
	);

	or_ii _1599_ (
		.a(_0768_),
		.b(_0767_),
		.c(_0769_)
	);

	and_ii _1600_ (
		.a(new_net_496),
		.b(new_net_668),
		.c(_0770_)
	);

	or_bb _1601_ (
		.a(new_net_714),
		.b(new_net_47),
		.c(_0771_)
	);

	and_bi _1602_ (
		.a(_0769_),
		.b(new_net_1458),
		.c(_0772_)
	);

	or_bi _1603_ (
		.a(new_net_263),
		.b(new_net_282),
		.c(_0773_)
	);

	and_ii _1604_ (
		.a(new_net_68),
		.b(new_net_276),
		.c(_0774_)
	);

	and_bi _1605_ (
		.a(new_net_1459),
		.b(_0774_),
		.c(_0776_)
	);

	and_bi _1606_ (
		.a(new_net_715),
		.b(_0776_),
		.c(_0777_)
	);

	or_ii _1607_ (
		.a(new_net_771),
		.b(new_net_910),
		.c(_0778_)
	);

	and_bi _1608_ (
		.a(new_net_459),
		.b(_0778_),
		.c(_0779_)
	);

	or_bb _1609_ (
		.a(new_net_1460),
		.b(_0777_),
		.c(_0780_)
	);

	or_bb _1610_ (
		.a(new_net_1461),
		.b(_0772_),
		.c(new_net_1485)
	);

	or_ii _1611_ (
		.a(new_net_640),
		.b(new_net_208),
		.c(_0781_)
	);

	and_ii _1612_ (
		.a(new_net_641),
		.b(new_net_209),
		.c(_0782_)
	);

	or_bi _1613_ (
		.a(_0782_),
		.b(new_net_10),
		.c(_0783_)
	);

	and_bi _1614_ (
		.a(new_net_1462),
		.b(_0783_),
		.c(_0784_)
	);

	or_ii _1615_ (
		.a(new_net_327),
		.b(new_net_704),
		.c(_0786_)
	);

	or_bb _1616_ (
		.a(new_net_328),
		.b(new_net_702),
		.c(_0787_)
	);

	or_ii _1617_ (
		.a(_0787_),
		.b(_0786_),
		.c(G3539)
	);

	spl2 _0784__v_fanout (
		.a(_0784_),
		.b(new_net_328),
		.c(new_net_327)
	);

	spl2 new_net_1254_v_fanout (
		.a(new_net_1254),
		.b(new_net_704),
		.c(new_net_702)
	);

	bfr new_net_1487_bfr_before (
		.din(new_net_1487),
		.dout(new_net_1254)
	);

	spl3L _0753__v_fanout (
		.a(_0753_),
		.b(new_net_703),
		.c(new_net_1487),
		.d(new_net_701)
	);

	spl2 new_net_1253_v_fanout (
		.a(new_net_1253),
		.b(new_net_642),
		.c(new_net_639)
	);

	spl2 _0735__v_fanout (
		.a(_0735_),
		.b(new_net_998),
		.c(new_net_997)
	);

	bfr new_net_1488_bfr_before (
		.din(new_net_1488),
		.dout(new_net_1253)
	);

	spl3L _0740__v_fanout (
		.a(_0740_),
		.b(new_net_1488),
		.c(new_net_640),
		.d(new_net_641)
	);

	spl2 _0742__v_fanout (
		.a(_0742_),
		.b(new_net_66),
		.c(new_net_65)
	);

	spl3L _0464__v_fanout (
		.a(_0464_),
		.b(new_net_878),
		.c(new_net_877),
		.d(new_net_876)
	);

	bfr new_net_1489_bfr_after (
		.din(_0750_),
		.dout(new_net_1489)
	);

	bfr new_net_1490_bfr_after (
		.din(new_net_1489),
		.dout(new_net_1490)
	);

	spl2 _0750__v_fanout (
		.a(new_net_1490),
		.b(new_net_729),
		.c(new_net_728)
	);

	spl2 _0541__v_fanout (
		.a(_0541_),
		.b(new_net_749),
		.c(new_net_748)
	);

	bfr new_net_1491_bfr_before (
		.din(new_net_1491),
		.dout(G3534)
	);

	bfr new_net_1492_bfr_before (
		.din(new_net_1492),
		.dout(new_net_1491)
	);

	bfr new_net_1493_bfr_before (
		.din(new_net_1493),
		.dout(new_net_1492)
	);

	bfr new_net_1494_bfr_before (
		.din(new_net_1494),
		.dout(new_net_1493)
	);

	bfr new_net_1495_bfr_before (
		.din(new_net_1495),
		.dout(new_net_1494)
	);

	bfr new_net_1496_bfr_before (
		.din(new_net_1496),
		.dout(new_net_1495)
	);

	bfr new_net_1497_bfr_before (
		.din(new_net_1497),
		.dout(new_net_1496)
	);

	bfr new_net_1498_bfr_before (
		.din(new_net_1498),
		.dout(new_net_1497)
	);

	bfr new_net_1499_bfr_before (
		.din(new_net_1499),
		.dout(new_net_1498)
	);

	bfr new_net_1500_bfr_before (
		.din(new_net_1500),
		.dout(new_net_1499)
	);

	spl3L new_net_1_v_fanout (
		.a(new_net_1),
		.b(new_net_900),
		.c(new_net_901),
		.d(new_net_1500)
	);

	bfr new_net_1501_bfr_before (
		.din(new_net_1501),
		.dout(G3536)
	);

	bfr new_net_1502_bfr_before (
		.din(new_net_1502),
		.dout(new_net_1501)
	);

	bfr new_net_1503_bfr_before (
		.din(new_net_1503),
		.dout(new_net_1502)
	);

	bfr new_net_1504_bfr_before (
		.din(new_net_1504),
		.dout(new_net_1503)
	);

	bfr new_net_1505_bfr_before (
		.din(new_net_1505),
		.dout(new_net_1504)
	);

	bfr new_net_1506_bfr_before (
		.din(new_net_1506),
		.dout(new_net_1505)
	);

	bfr new_net_1507_bfr_before (
		.din(new_net_1507),
		.dout(new_net_1506)
	);

	bfr new_net_1508_bfr_before (
		.din(new_net_1508),
		.dout(new_net_1507)
	);

	bfr new_net_1509_bfr_before (
		.din(new_net_1509),
		.dout(new_net_1508)
	);

	bfr new_net_1510_bfr_before (
		.din(new_net_1510),
		.dout(new_net_1509)
	);

	bfr new_net_1511_bfr_before (
		.din(new_net_1511),
		.dout(new_net_1510)
	);

	spl3L new_net_2_v_fanout (
		.a(new_net_2),
		.b(new_net_872),
		.c(new_net_873),
		.d(new_net_1511)
	);

	bfr new_net_1512_bfr_after (
		.din(new_net_0),
		.dout(new_net_1512)
	);

	bfr new_net_1513_bfr_before (
		.din(new_net_1513),
		.dout(G3535)
	);

	bfr new_net_1514_bfr_before (
		.din(new_net_1514),
		.dout(new_net_1513)
	);

	bfr new_net_1515_bfr_before (
		.din(new_net_1515),
		.dout(new_net_1514)
	);

	bfr new_net_1516_bfr_before (
		.din(new_net_1516),
		.dout(new_net_1515)
	);

	bfr new_net_1517_bfr_before (
		.din(new_net_1517),
		.dout(new_net_1516)
	);

	bfr new_net_1518_bfr_before (
		.din(new_net_1518),
		.dout(new_net_1517)
	);

	bfr new_net_1519_bfr_before (
		.din(new_net_1519),
		.dout(new_net_1518)
	);

	bfr new_net_1520_bfr_before (
		.din(new_net_1520),
		.dout(new_net_1519)
	);

	bfr new_net_1521_bfr_before (
		.din(new_net_1521),
		.dout(new_net_1520)
	);

	bfr new_net_1522_bfr_before (
		.din(new_net_1522),
		.dout(new_net_1521)
	);

	spl3L new_net_0_v_fanout (
		.a(new_net_1512),
		.b(new_net_373),
		.c(new_net_374),
		.d(new_net_1522)
	);

	spl2 _0747__v_fanout (
		.a(_0747_),
		.b(new_net_557),
		.c(new_net_556)
	);

	spl2 _0663__v_fanout (
		.a(_0663_),
		.b(new_net_679),
		.c(new_net_678)
	);

	spl2 _0354__v_fanout (
		.a(_0354_),
		.b(new_net_778),
		.c(new_net_777)
	);

	spl2 new_net_1252_v_fanout (
		.a(new_net_1252),
		.b(new_net_581),
		.c(new_net_580)
	);

	spl2 _0350__v_fanout (
		.a(_0350_),
		.b(new_net_670),
		.c(new_net_669)
	);

	bfr new_net_1523_bfr_before (
		.din(new_net_1523),
		.dout(new_net_555)
	);

	bfr new_net_1524_bfr_before (
		.din(new_net_1524),
		.dout(new_net_1523)
	);

	spl2 _0450__v_fanout (
		.a(_0450_),
		.b(new_net_1524),
		.c(new_net_554)
	);

	bfr new_net_1525_bfr_before (
		.din(new_net_1525),
		.dout(G3531)
	);

	bfr new_net_1526_bfr_before (
		.din(new_net_1526),
		.dout(new_net_1525)
	);

	bfr new_net_1527_bfr_before (
		.din(new_net_1527),
		.dout(new_net_1526)
	);

	bfr new_net_1528_bfr_before (
		.din(new_net_1528),
		.dout(new_net_1527)
	);

	bfr new_net_1529_bfr_before (
		.din(new_net_1529),
		.dout(new_net_1528)
	);

	bfr new_net_1530_bfr_before (
		.din(new_net_1530),
		.dout(new_net_1529)
	);

	bfr new_net_1531_bfr_before (
		.din(new_net_1531),
		.dout(new_net_1530)
	);

	bfr new_net_1532_bfr_before (
		.din(new_net_1532),
		.dout(new_net_1531)
	);

	bfr new_net_1533_bfr_before (
		.din(new_net_1533),
		.dout(new_net_1532)
	);

	bfr new_net_1534_bfr_before (
		.din(new_net_1534),
		.dout(new_net_1533)
	);

	bfr new_net_1535_bfr_before (
		.din(new_net_1535),
		.dout(new_net_1534)
	);

	bfr new_net_1536_bfr_before (
		.din(new_net_1536),
		.dout(new_net_1535)
	);

	bfr new_net_1537_bfr_before (
		.din(new_net_1537),
		.dout(new_net_1536)
	);

	bfr new_net_1538_bfr_before (
		.din(new_net_1538),
		.dout(new_net_1537)
	);

	bfr new_net_1539_bfr_before (
		.din(new_net_1539),
		.dout(new_net_1538)
	);

	bfr new_net_1540_bfr_before (
		.din(new_net_1540),
		.dout(new_net_1539)
	);

	spl3L new_net_5_v_fanout (
		.a(new_net_5),
		.b(new_net_500),
		.c(new_net_501),
		.d(new_net_1540)
	);

	spl2 new_net_1197_v_fanout (
		.a(new_net_1197),
		.b(new_net_923),
		.c(new_net_919)
	);

	spl2 new_net_1228_v_fanout (
		.a(new_net_1228),
		.b(new_net_21),
		.c(new_net_20)
	);

	bfr new_net_1541_bfr_after (
		.din(_0744_),
		.dout(new_net_1541)
	);

	bfr new_net_1542_bfr_after (
		.din(new_net_1541),
		.dout(new_net_1542)
	);

	bfr new_net_1543_bfr_after (
		.din(new_net_1542),
		.dout(new_net_1543)
	);

	bfr new_net_1544_bfr_after (
		.din(new_net_1543),
		.dout(new_net_1544)
	);

	bfr new_net_1545_bfr_after (
		.din(new_net_1544),
		.dout(new_net_1545)
	);

	spl2 _0744__v_fanout (
		.a(new_net_1545),
		.b(new_net_426),
		.c(new_net_425)
	);

	bfr new_net_1546_bfr_after (
		.din(new_net_6),
		.dout(new_net_1546)
	);

	bfr new_net_1547_bfr_after (
		.din(new_net_1546),
		.dout(new_net_1547)
	);

	bfr new_net_1548_bfr_before (
		.din(new_net_1548),
		.dout(G3533)
	);

	bfr new_net_1549_bfr_before (
		.din(new_net_1549),
		.dout(new_net_1548)
	);

	bfr new_net_1550_bfr_before (
		.din(new_net_1550),
		.dout(new_net_1549)
	);

	bfr new_net_1551_bfr_before (
		.din(new_net_1551),
		.dout(new_net_1550)
	);

	bfr new_net_1552_bfr_before (
		.din(new_net_1552),
		.dout(new_net_1551)
	);

	bfr new_net_1553_bfr_before (
		.din(new_net_1553),
		.dout(new_net_1552)
	);

	bfr new_net_1554_bfr_before (
		.din(new_net_1554),
		.dout(new_net_1553)
	);

	bfr new_net_1555_bfr_before (
		.din(new_net_1555),
		.dout(new_net_1554)
	);

	bfr new_net_1556_bfr_before (
		.din(new_net_1556),
		.dout(new_net_1555)
	);

	bfr new_net_1557_bfr_before (
		.din(new_net_1557),
		.dout(new_net_1556)
	);

	bfr new_net_1558_bfr_before (
		.din(new_net_1558),
		.dout(new_net_1557)
	);

	bfr new_net_1559_bfr_before (
		.din(new_net_1559),
		.dout(new_net_1558)
	);

	bfr new_net_1560_bfr_before (
		.din(new_net_1560),
		.dout(new_net_1559)
	);

	bfr new_net_1561_bfr_before (
		.din(new_net_1561),
		.dout(new_net_1560)
	);

	bfr new_net_1562_bfr_before (
		.din(new_net_1562),
		.dout(new_net_1561)
	);

	bfr new_net_1563_bfr_before (
		.din(new_net_1563),
		.dout(new_net_1562)
	);

	spl3L new_net_6_v_fanout (
		.a(new_net_1547),
		.b(new_net_531),
		.c(new_net_532),
		.d(new_net_1563)
	);

	spl2 new_net_1251_v_fanout (
		.a(new_net_1251),
		.b(new_net_587),
		.c(new_net_585)
	);

	spl3L _0346__v_fanout (
		.a(_0346_),
		.b(new_net_452),
		.c(new_net_453),
		.d(new_net_451)
	);

	bfr new_net_1564_bfr_after (
		.din(new_net_3),
		.dout(new_net_1564)
	);

	bfr new_net_1565_bfr_after (
		.din(new_net_1564),
		.dout(new_net_1565)
	);

	bfr new_net_1566_bfr_after (
		.din(new_net_1565),
		.dout(new_net_1566)
	);

	bfr new_net_1567_bfr_after (
		.din(new_net_1566),
		.dout(new_net_1567)
	);

	bfr new_net_1568_bfr_after (
		.din(new_net_1567),
		.dout(new_net_1568)
	);

	bfr new_net_1569_bfr_after (
		.din(new_net_1568),
		.dout(new_net_1569)
	);

	bfr new_net_1570_bfr_after (
		.din(new_net_1569),
		.dout(new_net_1570)
	);

	bfr new_net_1571_bfr_after (
		.din(new_net_1570),
		.dout(new_net_1571)
	);

	bfr new_net_1572_bfr_before (
		.din(new_net_1572),
		.dout(G3529)
	);

	bfr new_net_1573_bfr_before (
		.din(new_net_1573),
		.dout(new_net_1572)
	);

	bfr new_net_1574_bfr_before (
		.din(new_net_1574),
		.dout(new_net_1573)
	);

	bfr new_net_1575_bfr_before (
		.din(new_net_1575),
		.dout(new_net_1574)
	);

	bfr new_net_1576_bfr_before (
		.din(new_net_1576),
		.dout(new_net_1575)
	);

	bfr new_net_1577_bfr_before (
		.din(new_net_1577),
		.dout(new_net_1576)
	);

	bfr new_net_1578_bfr_before (
		.din(new_net_1578),
		.dout(new_net_1577)
	);

	bfr new_net_1579_bfr_before (
		.din(new_net_1579),
		.dout(new_net_1578)
	);

	bfr new_net_1580_bfr_before (
		.din(new_net_1580),
		.dout(new_net_1579)
	);

	bfr new_net_1581_bfr_before (
		.din(new_net_1581),
		.dout(new_net_1580)
	);

	bfr new_net_1582_bfr_before (
		.din(new_net_1582),
		.dout(new_net_1581)
	);

	spl3L new_net_3_v_fanout (
		.a(new_net_1571),
		.b(new_net_106),
		.c(new_net_107),
		.d(new_net_1582)
	);

	bfr new_net_1583_bfr_before (
		.din(new_net_1583),
		.dout(new_net_854)
	);

	bfr new_net_1584_bfr_before (
		.din(new_net_1584),
		.dout(new_net_1583)
	);

	bfr new_net_1585_bfr_before (
		.din(new_net_1585),
		.dout(new_net_1584)
	);

	bfr new_net_1586_bfr_before (
		.din(new_net_1586),
		.dout(new_net_1585)
	);

	bfr new_net_1587_bfr_before (
		.din(new_net_1587),
		.dout(new_net_1586)
	);

	spl2 _0732__v_fanout (
		.a(_0732_),
		.b(new_net_855),
		.c(new_net_1587)
	);

	bfr new_net_1588_bfr_before (
		.din(new_net_1588),
		.dout(new_net_1197)
	);

	bfr new_net_1589_bfr_before (
		.din(new_net_1589),
		.dout(new_net_1588)
	);

	spl2 new_net_1196_v_fanout (
		.a(new_net_1196),
		.b(new_net_922),
		.c(new_net_1589)
	);

	bfr new_net_1590_bfr_before (
		.din(new_net_1590),
		.dout(new_net_1196)
	);

	spl2 new_net_1195_v_fanout (
		.a(new_net_1195),
		.b(new_net_920),
		.c(new_net_1590)
	);

	bfr new_net_1591_bfr_before (
		.din(new_net_1591),
		.dout(new_net_1252)
	);

	bfr new_net_1592_bfr_before (
		.din(new_net_1592),
		.dout(new_net_1591)
	);

	bfr new_net_1593_bfr_before (
		.din(new_net_1593),
		.dout(new_net_1592)
	);

	bfr new_net_1594_bfr_before (
		.din(new_net_1594),
		.dout(new_net_1593)
	);

	bfr new_net_1595_bfr_before (
		.din(new_net_1595),
		.dout(new_net_1594)
	);

	spl2 _0332__v_fanout (
		.a(_0332_),
		.b(new_net_1595),
		.c(new_net_582)
	);

	bfr new_net_1596_bfr_before (
		.din(new_net_1596),
		.dout(new_net_1228)
	);

	bfr new_net_1597_bfr_before (
		.din(new_net_1597),
		.dout(new_net_1596)
	);

	spl2 new_net_1227_v_fanout (
		.a(new_net_1227),
		.b(new_net_1597),
		.c(new_net_23)
	);

	spl2 _0343__v_fanout (
		.a(_0343_),
		.b(new_net_182),
		.c(new_net_181)
	);

	bfr new_net_1598_bfr_before (
		.din(new_net_1598),
		.dout(G3532)
	);

	bfr new_net_1599_bfr_before (
		.din(new_net_1599),
		.dout(new_net_1598)
	);

	bfr new_net_1600_bfr_before (
		.din(new_net_1600),
		.dout(new_net_1599)
	);

	bfr new_net_1601_bfr_before (
		.din(new_net_1601),
		.dout(new_net_1600)
	);

	bfr new_net_1602_bfr_before (
		.din(new_net_1602),
		.dout(new_net_1601)
	);

	bfr new_net_1603_bfr_before (
		.din(new_net_1603),
		.dout(new_net_1602)
	);

	bfr new_net_1604_bfr_before (
		.din(new_net_1604),
		.dout(new_net_1603)
	);

	bfr new_net_1605_bfr_before (
		.din(new_net_1605),
		.dout(new_net_1604)
	);

	bfr new_net_1606_bfr_before (
		.din(new_net_1606),
		.dout(new_net_1605)
	);

	bfr new_net_1607_bfr_before (
		.din(new_net_1607),
		.dout(new_net_1606)
	);

	bfr new_net_1608_bfr_before (
		.din(new_net_1608),
		.dout(new_net_1607)
	);

	bfr new_net_1609_bfr_before (
		.din(new_net_1609),
		.dout(new_net_1608)
	);

	bfr new_net_1610_bfr_before (
		.din(new_net_1610),
		.dout(new_net_1609)
	);

	bfr new_net_1611_bfr_before (
		.din(new_net_1611),
		.dout(new_net_1610)
	);

	bfr new_net_1612_bfr_before (
		.din(new_net_1612),
		.dout(new_net_1611)
	);

	bfr new_net_1613_bfr_before (
		.din(new_net_1613),
		.dout(new_net_1612)
	);

	bfr new_net_1614_bfr_before (
		.din(new_net_1614),
		.dout(new_net_1613)
	);

	bfr new_net_1615_bfr_before (
		.din(new_net_1615),
		.dout(new_net_1614)
	);

	bfr new_net_1616_bfr_before (
		.din(new_net_1616),
		.dout(new_net_1615)
	);

	bfr new_net_1617_bfr_before (
		.din(new_net_1617),
		.dout(new_net_1616)
	);

	bfr new_net_1618_bfr_before (
		.din(new_net_1618),
		.dout(new_net_1617)
	);

	spl3L new_net_7_v_fanout (
		.a(new_net_7),
		.b(new_net_751),
		.c(new_net_752),
		.d(new_net_1618)
	);

	spl2 _0766__v_fanout (
		.a(_0766_),
		.b(new_net_766),
		.c(new_net_765)
	);

	spl3L _0564__v_fanout (
		.a(_0564_),
		.b(new_net_124),
		.c(new_net_123),
		.d(new_net_122)
	);

	spl2 new_net_1250_v_fanout (
		.a(new_net_1250),
		.b(new_net_930),
		.c(new_net_929)
	);

	spl2 _0625__v_fanout (
		.a(_0625_),
		.b(new_net_346),
		.c(new_net_345)
	);

	bfr new_net_1619_bfr_after (
		.din(_0349_),
		.dout(new_net_1619)
	);

	bfr new_net_1620_bfr_after (
		.din(new_net_1619),
		.dout(new_net_1620)
	);

	bfr new_net_1621_bfr_after (
		.din(new_net_1620),
		.dout(new_net_1621)
	);

	bfr new_net_1622_bfr_before (
		.din(new_net_1622),
		.dout(new_net_1251)
	);

	spl2 _0349__v_fanout (
		.a(new_net_1621),
		.b(new_net_586),
		.c(new_net_1622)
	);

	bfr new_net_1623_bfr_before (
		.din(new_net_1623),
		.dout(new_net_324)
	);

	spl3L _0322__v_fanout (
		.a(_0322_),
		.b(new_net_325),
		.c(new_net_326),
		.d(new_net_1623)
	);

	bfr new_net_1624_bfr_after (
		.din(_0762_),
		.dout(new_net_1624)
	);

	spl2 _0762__v_fanout (
		.a(new_net_1624),
		.b(new_net_837),
		.c(new_net_836)
	);

	spl2 _0323__v_fanout (
		.a(_0323_),
		.b(new_net_379),
		.c(new_net_378)
	);

	spl2 _0563__v_fanout (
		.a(_0563_),
		.b(new_net_1250),
		.c(new_net_928)
	);

	spl2 _0501__v_fanout (
		.a(_0501_),
		.b(new_net_868),
		.c(new_net_867)
	);

	bfr new_net_1625_bfr_before (
		.din(new_net_1625),
		.dout(new_net_27)
	);

	bfr new_net_1626_bfr_before (
		.din(new_net_1626),
		.dout(new_net_1625)
	);

	bfr new_net_1627_bfr_before (
		.din(new_net_1627),
		.dout(new_net_1626)
	);

	spl2 _0611__v_fanout (
		.a(_0611_),
		.b(new_net_28),
		.c(new_net_1627)
	);

	bfr new_net_1628_bfr_after (
		.din(_0459_),
		.dout(new_net_1628)
	);

	spl2 _0459__v_fanout (
		.a(new_net_1628),
		.b(new_net_698),
		.c(new_net_697)
	);

	bfr new_net_1629_bfr_after (
		.din(_0340_),
		.dout(new_net_1629)
	);

	bfr new_net_1630_bfr_after (
		.din(new_net_1629),
		.dout(new_net_1630)
	);

	bfr new_net_1631_bfr_after (
		.din(new_net_1630),
		.dout(new_net_1631)
	);

	spl2 _0340__v_fanout (
		.a(new_net_1631),
		.b(new_net_455),
		.c(new_net_454)
	);

	bfr new_net_1632_bfr_before (
		.din(new_net_1632),
		.dout(new_net_1195)
	);

	bfr new_net_1633_bfr_before (
		.din(new_net_1633),
		.dout(new_net_1632)
	);

	bfr new_net_1634_bfr_before (
		.din(new_net_1634),
		.dout(new_net_1633)
	);

	spl2 new_net_1194_v_fanout (
		.a(new_net_1194),
		.b(new_net_1634),
		.c(new_net_921)
	);

	spl2 new_net_1247_v_fanout (
		.a(new_net_1247),
		.b(new_net_1005),
		.c(new_net_1006)
	);

	spl3L new_net_1249_v_fanout (
		.a(new_net_1249),
		.b(new_net_942),
		.c(new_net_945),
		.d(new_net_941)
	);

	bfr new_net_1635_bfr_before (
		.din(new_net_1635),
		.dout(new_net_1227)
	);

	bfr new_net_1636_bfr_before (
		.din(new_net_1636),
		.dout(new_net_1635)
	);

	bfr new_net_1637_bfr_before (
		.din(new_net_1637),
		.dout(new_net_1636)
	);

	bfr new_net_1638_bfr_before (
		.din(new_net_1638),
		.dout(new_net_1637)
	);

	bfr new_net_1639_bfr_before (
		.din(new_net_1639),
		.dout(new_net_1638)
	);

	spl3L new_net_1226_v_fanout (
		.a(new_net_1226),
		.b(new_net_22),
		.c(new_net_19),
		.d(new_net_1639)
	);

	bfr new_net_1640_bfr_before (
		.din(new_net_1640),
		.dout(new_net_256)
	);

	spl3L _0572__v_fanout (
		.a(_0572_),
		.b(new_net_1640),
		.c(new_net_257),
		.d(new_net_255)
	);

	spl3L _0348__v_fanout (
		.a(_0348_),
		.b(new_net_545),
		.c(new_net_546),
		.d(new_net_544)
	);

	spl2 new_net_1248_v_fanout (
		.a(new_net_1248),
		.b(new_net_943),
		.c(new_net_944)
	);

	spl2 new_net_1240_v_fanout (
		.a(new_net_1240),
		.b(new_net_650),
		.c(new_net_649)
	);

	spl2 _0339__v_fanout (
		.a(_0339_),
		.b(new_net_119),
		.c(new_net_118)
	);

	spl2 _0561__v_fanout (
		.a(_0561_),
		.b(new_net_434),
		.c(new_net_433)
	);

	spl2 _0616__v_fanout (
		.a(_0616_),
		.b(new_net_339),
		.c(new_net_338)
	);

	bfr new_net_1641_bfr_after (
		.din(_0499_),
		.dout(new_net_1641)
	);

	bfr new_net_1642_bfr_after (
		.din(new_net_1641),
		.dout(new_net_1642)
	);

	spl2 _0499__v_fanout (
		.a(new_net_1642),
		.b(new_net_457),
		.c(new_net_456)
	);

	spl2 _0305__v_fanout (
		.a(_0305_),
		.b(new_net_1249),
		.c(new_net_1248)
	);

	bfr new_net_1643_bfr_after (
		.din(new_net_8),
		.dout(new_net_1643)
	);

	bfr new_net_1644_bfr_after (
		.din(new_net_1643),
		.dout(new_net_1644)
	);

	bfr new_net_1645_bfr_after (
		.din(new_net_1644),
		.dout(new_net_1645)
	);

	bfr new_net_1646_bfr_after (
		.din(new_net_1645),
		.dout(new_net_1646)
	);

	bfr new_net_1647_bfr_after (
		.din(new_net_1646),
		.dout(new_net_1647)
	);

	bfr new_net_1648_bfr_after (
		.din(new_net_1647),
		.dout(new_net_1648)
	);

	bfr new_net_1649_bfr_before (
		.din(new_net_1649),
		.dout(G3528)
	);

	bfr new_net_1650_bfr_before (
		.din(new_net_1650),
		.dout(new_net_1649)
	);

	bfr new_net_1651_bfr_before (
		.din(new_net_1651),
		.dout(new_net_1650)
	);

	bfr new_net_1652_bfr_before (
		.din(new_net_1652),
		.dout(new_net_1651)
	);

	bfr new_net_1653_bfr_before (
		.din(new_net_1653),
		.dout(new_net_1652)
	);

	bfr new_net_1654_bfr_before (
		.din(new_net_1654),
		.dout(new_net_1653)
	);

	bfr new_net_1655_bfr_before (
		.din(new_net_1655),
		.dout(new_net_1654)
	);

	bfr new_net_1656_bfr_before (
		.din(new_net_1656),
		.dout(new_net_1655)
	);

	bfr new_net_1657_bfr_before (
		.din(new_net_1657),
		.dout(new_net_1656)
	);

	bfr new_net_1658_bfr_before (
		.din(new_net_1658),
		.dout(new_net_1657)
	);

	bfr new_net_1659_bfr_before (
		.din(new_net_1659),
		.dout(new_net_1658)
	);

	bfr new_net_1660_bfr_before (
		.din(new_net_1660),
		.dout(new_net_1659)
	);

	bfr new_net_1661_bfr_before (
		.din(new_net_1661),
		.dout(new_net_1660)
	);

	bfr new_net_1662_bfr_before (
		.din(new_net_1662),
		.dout(new_net_1661)
	);

	bfr new_net_1663_bfr_before (
		.din(new_net_1663),
		.dout(new_net_1662)
	);

	bfr new_net_1664_bfr_before (
		.din(new_net_1664),
		.dout(new_net_1663)
	);

	bfr new_net_1665_bfr_before (
		.din(new_net_1665),
		.dout(new_net_1664)
	);

	bfr new_net_1666_bfr_before (
		.din(new_net_1666),
		.dout(new_net_1665)
	);

	bfr new_net_1667_bfr_before (
		.din(new_net_1667),
		.dout(new_net_1666)
	);

	bfr new_net_1668_bfr_before (
		.din(new_net_1668),
		.dout(new_net_1667)
	);

	bfr new_net_1669_bfr_before (
		.din(new_net_1669),
		.dout(new_net_1668)
	);

	spl3L new_net_8_v_fanout (
		.a(new_net_1648),
		.b(new_net_976),
		.c(new_net_977),
		.d(new_net_1669)
	);

	bfr new_net_1670_bfr_before (
		.din(new_net_1670),
		.dout(new_net_1247)
	);

	spl3L _0456__v_fanout (
		.a(_0456_),
		.b(new_net_1670),
		.c(new_net_1004),
		.d(new_net_1003)
	);

	bfr new_net_1671_bfr_before (
		.din(new_net_1671),
		.dout(new_net_1024)
	);

	bfr new_net_1672_bfr_before (
		.din(new_net_1672),
		.dout(new_net_1671)
	);

	bfr new_net_1673_bfr_before (
		.din(new_net_1673),
		.dout(new_net_1672)
	);

	bfr new_net_1674_bfr_before (
		.din(new_net_1674),
		.dout(new_net_1673)
	);

	bfr new_net_1675_bfr_before (
		.din(new_net_1675),
		.dout(new_net_1674)
	);

	spl4L new_net_1246_v_fanout (
		.a(new_net_1246),
		.b(new_net_1028),
		.c(new_net_1026),
		.d(new_net_1675),
		.e(new_net_1023)
	);

	spl3L _0571__v_fanout (
		.a(_0571_),
		.b(new_net_215),
		.c(new_net_216),
		.d(new_net_214)
	);

	spl2 new_net_1242_v_fanout (
		.a(new_net_1242),
		.b(new_net_726),
		.c(new_net_727)
	);

	bfr new_net_1676_bfr_before (
		.din(new_net_1676),
		.dout(new_net_646)
	);

	bfr new_net_1677_bfr_before (
		.din(new_net_1677),
		.dout(new_net_1676)
	);

	bfr new_net_1678_bfr_before (
		.din(new_net_1678),
		.dout(new_net_1677)
	);

	spl2 new_net_1243_v_fanout (
		.a(new_net_1243),
		.b(new_net_645),
		.c(new_net_1678)
	);

	spl2 _0304__v_fanout (
		.a(_0304_),
		.b(new_net_440),
		.c(new_net_439)
	);

	spl2 _0559__v_fanout (
		.a(_0559_),
		.b(new_net_608),
		.c(new_net_607)
	);

	spl4L _0338__v_fanout (
		.a(_0338_),
		.b(new_net_1246),
		.c(new_net_1027),
		.d(new_net_1022),
		.e(new_net_1025)
	);

	spl2 _0328__v_fanout (
		.a(_0328_),
		.b(new_net_648),
		.c(new_net_647)
	);

	spl2 _0558__v_fanout (
		.a(_0558_),
		.b(new_net_754),
		.c(new_net_753)
	);

	spl2 _0568__v_fanout (
		.a(_0568_),
		.b(new_net_839),
		.c(new_net_838)
	);

	spl2 new_net_1244_v_fanout (
		.a(new_net_1244),
		.b(new_net_364),
		.c(new_net_362)
	);

	spl2 _0566__v_fanout (
		.a(_0566_),
		.b(new_net_936),
		.c(new_net_935)
	);

	bfr new_net_1679_bfr_before (
		.din(new_net_1679),
		.dout(new_net_1007)
	);

	bfr new_net_1680_bfr_before (
		.din(new_net_1680),
		.dout(new_net_1679)
	);

	bfr new_net_1681_bfr_before (
		.din(new_net_1681),
		.dout(new_net_1680)
	);

	bfr new_net_1682_bfr_before (
		.din(new_net_1682),
		.dout(new_net_1681)
	);

	bfr new_net_1683_bfr_before (
		.din(new_net_1683),
		.dout(new_net_1682)
	);

	spl3L _0321__v_fanout (
		.a(_0321_),
		.b(new_net_1009),
		.c(new_net_1008),
		.d(new_net_1683)
	);

	spl2 _0277__v_fanout (
		.a(_0277_),
		.b(new_net_121),
		.c(new_net_120)
	);

	bfr new_net_1684_bfr_after (
		.din(_0168_),
		.dout(new_net_1684)
	);

	bfr new_net_1685_bfr_before (
		.din(new_net_1685),
		.dout(new_net_1015)
	);

	bfr new_net_1686_bfr_before (
		.din(new_net_1686),
		.dout(new_net_1685)
	);

	spl3L _0168__v_fanout (
		.a(new_net_1684),
		.b(new_net_1686),
		.c(new_net_1014),
		.d(new_net_1013)
	);

	spl2 new_net_1241_v_fanout (
		.a(new_net_1241),
		.b(new_net_212),
		.c(new_net_213)
	);

	spl2 _0327__v_fanout (
		.a(_0327_),
		.b(new_net_561),
		.c(new_net_560)
	);

	bfr new_net_1687_bfr_before (
		.din(new_net_1687),
		.dout(new_net_969)
	);

	spl2 new_net_1245_v_fanout (
		.a(new_net_1245),
		.b(new_net_1687),
		.c(new_net_970)
	);

	bfr new_net_1688_bfr_after (
		.din(new_net_4),
		.dout(new_net_1688)
	);

	bfr new_net_1689_bfr_after (
		.din(new_net_1688),
		.dout(new_net_1689)
	);

	bfr new_net_1690_bfr_after (
		.din(new_net_1689),
		.dout(new_net_1690)
	);

	bfr new_net_1691_bfr_after (
		.din(new_net_1690),
		.dout(new_net_1691)
	);

	bfr new_net_1692_bfr_after (
		.din(new_net_1691),
		.dout(new_net_1692)
	);

	bfr new_net_1693_bfr_before (
		.din(new_net_1693),
		.dout(G3526)
	);

	bfr new_net_1694_bfr_before (
		.din(new_net_1694),
		.dout(new_net_1693)
	);

	bfr new_net_1695_bfr_before (
		.din(new_net_1695),
		.dout(new_net_1694)
	);

	bfr new_net_1696_bfr_before (
		.din(new_net_1696),
		.dout(new_net_1695)
	);

	bfr new_net_1697_bfr_before (
		.din(new_net_1697),
		.dout(new_net_1696)
	);

	bfr new_net_1698_bfr_before (
		.din(new_net_1698),
		.dout(new_net_1697)
	);

	bfr new_net_1699_bfr_before (
		.din(new_net_1699),
		.dout(new_net_1698)
	);

	bfr new_net_1700_bfr_before (
		.din(new_net_1700),
		.dout(new_net_1699)
	);

	bfr new_net_1701_bfr_before (
		.din(new_net_1701),
		.dout(new_net_1700)
	);

	bfr new_net_1702_bfr_before (
		.din(new_net_1702),
		.dout(new_net_1701)
	);

	bfr new_net_1703_bfr_before (
		.din(new_net_1703),
		.dout(new_net_1702)
	);

	bfr new_net_1704_bfr_before (
		.din(new_net_1704),
		.dout(new_net_1703)
	);

	bfr new_net_1705_bfr_before (
		.din(new_net_1705),
		.dout(new_net_1704)
	);

	bfr new_net_1706_bfr_before (
		.din(new_net_1706),
		.dout(new_net_1705)
	);

	bfr new_net_1707_bfr_before (
		.din(new_net_1707),
		.dout(new_net_1706)
	);

	bfr new_net_1708_bfr_before (
		.din(new_net_1708),
		.dout(new_net_1707)
	);

	bfr new_net_1709_bfr_before (
		.din(new_net_1709),
		.dout(new_net_1708)
	);

	bfr new_net_1710_bfr_before (
		.din(new_net_1710),
		.dout(new_net_1709)
	);

	bfr new_net_1711_bfr_before (
		.din(new_net_1711),
		.dout(new_net_1710)
	);

	bfr new_net_1712_bfr_before (
		.din(new_net_1712),
		.dout(new_net_1711)
	);

	bfr new_net_1713_bfr_before (
		.din(new_net_1713),
		.dout(new_net_1712)
	);

	bfr new_net_1714_bfr_before (
		.din(new_net_1714),
		.dout(new_net_1713)
	);

	bfr new_net_1715_bfr_before (
		.din(new_net_1715),
		.dout(new_net_1714)
	);

	bfr new_net_1716_bfr_before (
		.din(new_net_1716),
		.dout(new_net_1715)
	);

	bfr new_net_1717_bfr_before (
		.din(new_net_1717),
		.dout(new_net_1716)
	);

	bfr new_net_1718_bfr_before (
		.din(new_net_1718),
		.dout(new_net_1717)
	);

	spl3L new_net_4_v_fanout (
		.a(new_net_1692),
		.b(new_net_979),
		.c(new_net_980),
		.d(new_net_1718)
	);

	spl2 _0302__v_fanout (
		.a(_0302_),
		.b(new_net_359),
		.c(new_net_358)
	);

	bfr new_net_1719_bfr_before (
		.din(new_net_1719),
		.dout(new_net_875)
	);

	bfr new_net_1720_bfr_before (
		.din(new_net_1720),
		.dout(new_net_1719)
	);

	bfr new_net_1721_bfr_before (
		.din(new_net_1721),
		.dout(new_net_1720)
	);

	bfr new_net_1722_bfr_before (
		.din(new_net_1722),
		.dout(new_net_1721)
	);

	bfr new_net_1723_bfr_before (
		.din(new_net_1723),
		.dout(new_net_1722)
	);

	bfr new_net_1724_bfr_before (
		.din(new_net_1724),
		.dout(new_net_1723)
	);

	bfr new_net_1725_bfr_before (
		.din(new_net_1725),
		.dout(new_net_1724)
	);

	spl2 _0314__v_fanout (
		.a(_0314_),
		.b(new_net_1725),
		.c(new_net_874)
	);

	bfr new_net_1726_bfr_before (
		.din(new_net_1726),
		.dout(new_net_369)
	);

	bfr new_net_1727_bfr_before (
		.din(new_net_1727),
		.dout(new_net_1726)
	);

	spl2 _0565__v_fanout (
		.a(_0565_),
		.b(new_net_1727),
		.c(new_net_368)
	);

	spl2 _0556__v_fanout (
		.a(_0556_),
		.b(new_net_446),
		.c(new_net_445)
	);

	bfr new_net_1728_bfr_after (
		.din(_0284_),
		.dout(new_net_1728)
	);

	bfr new_net_1729_bfr_after (
		.din(new_net_1728),
		.dout(new_net_1729)
	);

	bfr new_net_1730_bfr_after (
		.din(new_net_1729),
		.dout(new_net_1730)
	);

	bfr new_net_1731_bfr_before (
		.din(new_net_1731),
		.dout(new_net_807)
	);

	bfr new_net_1732_bfr_before (
		.din(new_net_1732),
		.dout(new_net_1731)
	);

	spl2 _0284__v_fanout (
		.a(new_net_1730),
		.b(new_net_1732),
		.c(new_net_806)
	);

	bfr new_net_1733_bfr_before (
		.din(new_net_1733),
		.dout(new_net_344)
	);

	bfr new_net_1734_bfr_before (
		.din(new_net_1734),
		.dout(new_net_1733)
	);

	bfr new_net_1735_bfr_before (
		.din(new_net_1735),
		.dout(new_net_1734)
	);

	bfr new_net_1736_bfr_before (
		.din(new_net_1736),
		.dout(new_net_1735)
	);

	bfr new_net_1737_bfr_before (
		.din(new_net_1737),
		.dout(new_net_1736)
	);

	bfr new_net_1738_bfr_before (
		.din(new_net_1738),
		.dout(new_net_1737)
	);

	bfr new_net_1739_bfr_before (
		.din(new_net_1739),
		.dout(new_net_1738)
	);

	bfr new_net_1740_bfr_before (
		.din(new_net_1740),
		.dout(new_net_1739)
	);

	bfr new_net_1741_bfr_before (
		.din(new_net_1741),
		.dout(new_net_1740)
	);

	bfr new_net_1742_bfr_before (
		.din(new_net_1742),
		.dout(new_net_1741)
	);

	spl2 new_net_1221_v_fanout (
		.a(new_net_1221),
		.b(new_net_343),
		.c(new_net_1742)
	);

	spl2 _0251__v_fanout (
		.a(_0251_),
		.b(new_net_681),
		.c(new_net_680)
	);

	bfr new_net_1743_bfr_before (
		.din(new_net_1743),
		.dout(new_net_1245)
	);

	spl2 _0167__v_fanout (
		.a(_0167_),
		.b(new_net_1743),
		.c(new_net_968)
	);

	bfr new_net_1744_bfr_before (
		.din(new_net_1744),
		.dout(new_net_953)
	);

	spl3L _0545__v_fanout (
		.a(_0545_),
		.b(new_net_954),
		.c(new_net_955),
		.d(new_net_1744)
	);

	bfr new_net_1745_bfr_before (
		.din(new_net_1745),
		.dout(new_net_1241)
	);

	bfr new_net_1746_bfr_before (
		.din(new_net_1746),
		.dout(new_net_1745)
	);

	spl3L _0319__v_fanout (
		.a(_0319_),
		.b(new_net_211),
		.c(new_net_210),
		.d(new_net_1746)
	);

	bfr new_net_1747_bfr_before (
		.din(new_net_1747),
		.dout(new_net_711)
	);

	bfr new_net_1748_bfr_before (
		.din(new_net_1748),
		.dout(new_net_1747)
	);

	bfr new_net_1749_bfr_before (
		.din(new_net_1749),
		.dout(new_net_1748)
	);

	bfr new_net_1750_bfr_before (
		.din(new_net_1750),
		.dout(new_net_1749)
	);

	bfr new_net_1751_bfr_before (
		.din(new_net_1751),
		.dout(new_net_1750)
	);

	bfr new_net_1752_bfr_before (
		.din(new_net_1752),
		.dout(new_net_1751)
	);

	bfr new_net_1753_bfr_before (
		.din(new_net_1753),
		.dout(new_net_1752)
	);

	bfr new_net_1754_bfr_before (
		.din(new_net_1754),
		.dout(new_net_1753)
	);

	bfr new_net_1755_bfr_before (
		.din(new_net_1755),
		.dout(new_net_1754)
	);

	bfr new_net_1756_bfr_before (
		.din(new_net_1756),
		.dout(new_net_1755)
	);

	spl4L _0309__v_fanout (
		.a(_0309_),
		.b(new_net_1756),
		.c(new_net_709),
		.d(new_net_708),
		.e(new_net_710)
	);

	bfr new_net_1757_bfr_before (
		.din(new_net_1757),
		.dout(new_net_1240)
	);

	bfr new_net_1758_bfr_before (
		.din(new_net_1758),
		.dout(new_net_1757)
	);

	bfr new_net_1759_bfr_before (
		.din(new_net_1759),
		.dout(new_net_1758)
	);

	bfr new_net_1760_bfr_before (
		.din(new_net_1760),
		.dout(new_net_1759)
	);

	bfr new_net_1761_bfr_before (
		.din(new_net_1761),
		.dout(new_net_1760)
	);

	bfr new_net_1762_bfr_before (
		.din(new_net_1762),
		.dout(new_net_1761)
	);

	bfr new_net_1763_bfr_before (
		.din(new_net_1763),
		.dout(new_net_1762)
	);

	spl2 _0622__v_fanout (
		.a(_0622_),
		.b(new_net_651),
		.c(new_net_1763)
	);

	bfr new_net_1764_bfr_before (
		.din(new_net_1764),
		.dout(new_net_1243)
	);

	bfr new_net_1765_bfr_before (
		.din(new_net_1765),
		.dout(new_net_1764)
	);

	bfr new_net_1766_bfr_before (
		.din(new_net_1766),
		.dout(new_net_1765)
	);

	bfr new_net_1767_bfr_before (
		.din(new_net_1767),
		.dout(new_net_1766)
	);

	bfr new_net_1768_bfr_before (
		.din(new_net_1768),
		.dout(new_net_1767)
	);

	spl3L _0313__v_fanout (
		.a(_0313_),
		.b(new_net_1768),
		.c(new_net_644),
		.d(new_net_643)
	);

	bfr new_net_1769_bfr_before (
		.din(new_net_1769),
		.dout(new_net_1244)
	);

	bfr new_net_1770_bfr_before (
		.din(new_net_1770),
		.dout(new_net_1769)
	);

	bfr new_net_1771_bfr_before (
		.din(new_net_1771),
		.dout(new_net_1770)
	);

	spl2 _0554__v_fanout (
		.a(_0554_),
		.b(new_net_363),
		.c(new_net_1771)
	);

	spl4L _0549__v_fanout (
		.a(_0549_),
		.b(new_net_621),
		.c(new_net_622),
		.d(new_net_620),
		.e(new_net_623)
	);

	bfr new_net_1772_bfr_before (
		.din(new_net_1772),
		.dout(new_net_1242)
	);

	bfr new_net_1773_bfr_before (
		.din(new_net_1773),
		.dout(new_net_1772)
	);

	bfr new_net_1774_bfr_before (
		.din(new_net_1774),
		.dout(new_net_1773)
	);

	bfr new_net_1775_bfr_before (
		.din(new_net_1775),
		.dout(new_net_1774)
	);

	bfr new_net_1776_bfr_before (
		.din(new_net_1776),
		.dout(new_net_1775)
	);

	bfr new_net_1777_bfr_before (
		.din(new_net_1777),
		.dout(new_net_1776)
	);

	spl2 _0414__v_fanout (
		.a(_0414_),
		.b(new_net_1777),
		.c(new_net_725)
	);

	spl2 _0229__v_fanout (
		.a(_0229_),
		.b(new_net_880),
		.c(new_net_879)
	);

	spl2 _0115__v_fanout (
		.a(_0115_),
		.b(new_net_424),
		.c(new_net_423)
	);

	spl3L new_net_1234_v_fanout (
		.a(new_net_1234),
		.b(new_net_984),
		.c(new_net_988),
		.d(new_net_987)
	);

	bfr new_net_1778_bfr_before (
		.din(new_net_1778),
		.dout(new_net_996)
	);

	bfr new_net_1779_bfr_before (
		.din(new_net_1779),
		.dout(new_net_1778)
	);

	bfr new_net_1780_bfr_before (
		.din(new_net_1780),
		.dout(new_net_1779)
	);

	bfr new_net_1781_bfr_before (
		.din(new_net_1781),
		.dout(new_net_1780)
	);

	bfr new_net_1782_bfr_before (
		.din(new_net_1782),
		.dout(new_net_1781)
	);

	bfr new_net_1783_bfr_before (
		.din(new_net_1783),
		.dout(new_net_1782)
	);

	spl4L new_net_1066_v_fanout (
		.a(new_net_1066),
		.b(new_net_995),
		.c(new_net_1783),
		.d(new_net_992),
		.e(new_net_993)
	);

	spl2 new_net_1233_v_fanout (
		.a(new_net_1233),
		.b(new_net_981),
		.c(new_net_985)
	);

	spl3L _0228__v_fanout (
		.a(_0228_),
		.b(new_net_857),
		.c(new_net_858),
		.d(new_net_856)
	);

	bfr new_net_1784_bfr_before (
		.din(new_net_1784),
		.dout(new_net_323)
	);

	bfr new_net_1785_bfr_before (
		.din(new_net_1785),
		.dout(new_net_1784)
	);

	bfr new_net_1786_bfr_before (
		.din(new_net_1786),
		.dout(new_net_1785)
	);

	bfr new_net_1787_bfr_before (
		.din(new_net_1787),
		.dout(new_net_1786)
	);

	bfr new_net_1788_bfr_before (
		.din(new_net_1788),
		.dout(new_net_1787)
	);

	bfr new_net_1789_bfr_before (
		.din(new_net_1789),
		.dout(new_net_1788)
	);

	bfr new_net_1790_bfr_before (
		.din(new_net_1790),
		.dout(new_net_1789)
	);

	bfr new_net_1791_bfr_before (
		.din(new_net_1791),
		.dout(new_net_1790)
	);

	bfr new_net_1792_bfr_before (
		.din(new_net_1792),
		.dout(new_net_1791)
	);

	spl4L _0140__v_fanout (
		.a(_0140_),
		.b(new_net_321),
		.c(new_net_322),
		.d(new_net_320),
		.e(new_net_1792)
	);

	spl3L _0300__v_fanout (
		.a(_0300_),
		.b(new_net_550),
		.c(new_net_551),
		.d(new_net_549)
	);

	spl2 new_net_1235_v_fanout (
		.a(new_net_1235),
		.b(new_net_982),
		.c(new_net_986)
	);

	spl3L _0114__v_fanout (
		.a(_0114_),
		.b(new_net_206),
		.c(new_net_207),
		.d(new_net_205)
	);

	spl3L _0088__v_fanout (
		.a(_0088_),
		.b(new_net_195),
		.c(new_net_194),
		.d(new_net_193)
	);

	spl3L _0165__v_fanout (
		.a(_0165_),
		.b(new_net_863),
		.c(new_net_864),
		.d(new_net_862)
	);

	bfr new_net_1793_bfr_before (
		.din(new_net_1793),
		.dout(new_net_915)
	);

	bfr new_net_1794_bfr_before (
		.din(new_net_1794),
		.dout(new_net_1793)
	);

	spl4L _0250__v_fanout (
		.a(_0250_),
		.b(new_net_918),
		.c(new_net_916),
		.d(new_net_1794),
		.e(new_net_917)
	);

	spl3L _0200__v_fanout (
		.a(_0200_),
		.b(new_net_528),
		.c(new_net_529),
		.d(new_net_527)
	);

	spl3L new_net_1236_v_fanout (
		.a(new_net_1236),
		.b(new_net_983),
		.c(new_net_1234),
		.d(new_net_1233)
	);

	bfr new_net_1795_bfr_after (
		.din(_0325_),
		.dout(new_net_1795)
	);

	bfr new_net_1796_bfr_after (
		.din(new_net_1795),
		.dout(new_net_1796)
	);

	bfr new_net_1797_bfr_after (
		.din(new_net_1796),
		.dout(new_net_1797)
	);

	bfr new_net_1798_bfr_before (
		.din(new_net_1798),
		.dout(new_net_932)
	);

	bfr new_net_1799_bfr_before (
		.din(new_net_1799),
		.dout(new_net_1798)
	);

	bfr new_net_1800_bfr_before (
		.din(new_net_1800),
		.dout(new_net_1799)
	);

	bfr new_net_1801_bfr_before (
		.din(new_net_1801),
		.dout(new_net_1800)
	);

	bfr new_net_1802_bfr_before (
		.din(new_net_1802),
		.dout(new_net_1801)
	);

	bfr new_net_1803_bfr_before (
		.din(new_net_1803),
		.dout(new_net_1802)
	);

	bfr new_net_1804_bfr_before (
		.din(new_net_1804),
		.dout(new_net_1803)
	);

	bfr new_net_1805_bfr_before (
		.din(new_net_1805),
		.dout(new_net_1804)
	);

	spl2 _0325__v_fanout (
		.a(new_net_1797),
		.b(new_net_1805),
		.c(new_net_931)
	);

	bfr new_net_1806_bfr_before (
		.din(new_net_1806),
		.dout(new_net_1041)
	);

	bfr new_net_1807_bfr_before (
		.din(new_net_1807),
		.dout(new_net_1806)
	);

	bfr new_net_1808_bfr_before (
		.din(new_net_1808),
		.dout(new_net_1807)
	);

	spl2 _0555__v_fanout (
		.a(_0555_),
		.b(new_net_1042),
		.c(new_net_1808)
	);

	bfr new_net_1809_bfr_after (
		.din(_0618_),
		.dout(new_net_1809)
	);

	spl2 _0618__v_fanout (
		.a(new_net_1809),
		.b(new_net_432),
		.c(new_net_431)
	);

	bfr new_net_1810_bfr_before (
		.din(new_net_1810),
		.dout(new_net_82)
	);

	spl2 new_net_1178_v_fanout (
		.a(new_net_1178),
		.b(new_net_1810),
		.c(new_net_81)
	);

	spl2 _0084__v_fanout (
		.a(_0084_),
		.b(new_net_786),
		.c(new_net_785)
	);

	bfr new_net_1811_bfr_before (
		.din(new_net_1811),
		.dout(new_net_814)
	);

	spl3L _0164__v_fanout (
		.a(_0164_),
		.b(new_net_1811),
		.c(new_net_813),
		.d(new_net_812)
	);

	bfr new_net_1812_bfr_before (
		.din(new_net_1812),
		.dout(new_net_769)
	);

	bfr new_net_1813_bfr_before (
		.din(new_net_1813),
		.dout(new_net_1812)
	);

	bfr new_net_1814_bfr_before (
		.din(new_net_1814),
		.dout(new_net_1813)
	);

	bfr new_net_1815_bfr_before (
		.din(new_net_1815),
		.dout(new_net_1814)
	);

	spl3L _0247__v_fanout (
		.a(_0247_),
		.b(new_net_768),
		.c(new_net_1815),
		.d(new_net_767)
	);

	spl2 _0199__v_fanout (
		.a(_0199_),
		.b(new_net_468),
		.c(new_net_467)
	);

	bfr new_net_1816_bfr_after (
		.din(_0542_),
		.dout(new_net_1816)
	);

	bfr new_net_1817_bfr_after (
		.din(new_net_1816),
		.dout(new_net_1817)
	);

	spl2 _0542__v_fanout (
		.a(new_net_1817),
		.b(new_net_832),
		.c(new_net_831)
	);

	bfr new_net_1818_bfr_before (
		.din(new_net_1818),
		.dout(new_net_466)
	);

	spl2 _0087__v_fanout (
		.a(_0087_),
		.b(new_net_1818),
		.c(new_net_465)
	);

	bfr new_net_1819_bfr_after (
		.din(_0546_),
		.dout(new_net_1819)
	);

	bfr new_net_1820_bfr_after (
		.din(new_net_1819),
		.dout(new_net_1820)
	);

	spl2 _0546__v_fanout (
		.a(new_net_1820),
		.b(new_net_498),
		.c(new_net_497)
	);

	bfr new_net_1821_bfr_before (
		.din(new_net_1821),
		.dout(new_net_75)
	);

	bfr new_net_1822_bfr_before (
		.din(new_net_1822),
		.dout(new_net_78)
	);

	bfr new_net_1823_bfr_before (
		.din(new_net_1823),
		.dout(new_net_77)
	);

	spl4L new_net_1179_v_fanout (
		.a(new_net_1179),
		.b(new_net_76),
		.c(new_net_1823),
		.d(new_net_1821),
		.e(new_net_1822)
	);

	spl4L new_net_1224_v_fanout (
		.a(new_net_1224),
		.b(new_net_478),
		.c(new_net_479),
		.d(new_net_471),
		.e(new_net_480)
	);

	bfr new_net_1824_bfr_after (
		.din(_0551_),
		.dout(new_net_1824)
	);

	bfr new_net_1825_bfr_after (
		.din(new_net_1824),
		.dout(new_net_1825)
	);

	spl2 _0551__v_fanout (
		.a(new_net_1825),
		.b(new_net_229),
		.c(new_net_228)
	);

	spl3L _0139__v_fanout (
		.a(_0139_),
		.b(new_net_606),
		.c(new_net_605),
		.d(new_net_604)
	);

	spl3L _0225__v_fanout (
		.a(_0225_),
		.b(new_net_706),
		.c(new_net_707),
		.d(new_net_705)
	);

	bfr new_net_1826_bfr_before (
		.din(new_net_1826),
		.dout(new_net_630)
	);

	bfr new_net_1827_bfr_before (
		.din(new_net_1827),
		.dout(new_net_1826)
	);

	bfr new_net_1828_bfr_before (
		.din(new_net_1828),
		.dout(new_net_1827)
	);

	bfr new_net_1829_bfr_before (
		.din(new_net_1829),
		.dout(new_net_1828)
	);

	bfr new_net_1830_bfr_before (
		.din(new_net_1830),
		.dout(new_net_1829)
	);

	bfr new_net_1831_bfr_before (
		.din(new_net_1831),
		.dout(new_net_1830)
	);

	bfr new_net_1832_bfr_before (
		.din(new_net_1832),
		.dout(new_net_1831)
	);

	bfr new_net_1833_bfr_before (
		.din(new_net_1833),
		.dout(new_net_1832)
	);

	spl2 new_net_1220_v_fanout (
		.a(new_net_1220),
		.b(new_net_1833),
		.c(new_net_629)
	);

	spl3L _0113__v_fanout (
		.a(_0113_),
		.b(new_net_376),
		.c(new_net_377),
		.d(new_net_375)
	);

	bfr new_net_1834_bfr_after (
		.din(_0306_),
		.dout(new_net_1834)
	);

	bfr new_net_1835_bfr_after (
		.din(new_net_1834),
		.dout(new_net_1835)
	);

	spl2 _0306__v_fanout (
		.a(new_net_1835),
		.b(new_net_1000),
		.c(new_net_999)
	);

	bfr new_net_1836_bfr_before (
		.din(new_net_1836),
		.dout(new_net_584)
	);

	spl2 _0197__v_fanout (
		.a(_0197_),
		.b(new_net_1836),
		.c(new_net_583)
	);

	bfr new_net_1837_bfr_before (
		.din(new_net_1837),
		.dout(new_net_474)
	);

	bfr new_net_1838_bfr_before (
		.din(new_net_1838),
		.dout(new_net_1837)
	);

	bfr new_net_1839_bfr_before (
		.din(new_net_1839),
		.dout(new_net_1838)
	);

	bfr new_net_1840_bfr_before (
		.din(new_net_1840),
		.dout(new_net_1839)
	);

	bfr new_net_1841_bfr_before (
		.din(new_net_1841),
		.dout(new_net_1840)
	);

	bfr new_net_1842_bfr_before (
		.din(new_net_1842),
		.dout(new_net_1841)
	);

	bfr new_net_1843_bfr_before (
		.din(new_net_1843),
		.dout(new_net_1842)
	);

	bfr new_net_1844_bfr_before (
		.din(new_net_1844),
		.dout(new_net_1843)
	);

	bfr new_net_1845_bfr_before (
		.din(new_net_1845),
		.dout(new_net_1844)
	);

	spl2 new_net_1223_v_fanout (
		.a(new_net_1223),
		.b(new_net_481),
		.c(new_net_1845)
	);

	spl2 _0162__v_fanout (
		.a(_0162_),
		.b(new_net_870),
		.c(new_net_869)
	);

	bfr new_net_1846_bfr_before (
		.din(new_net_1846),
		.dout(new_net_885)
	);

	bfr new_net_1847_bfr_before (
		.din(new_net_1847),
		.dout(new_net_1846)
	);

	bfr new_net_1848_bfr_before (
		.din(new_net_1848),
		.dout(new_net_1847)
	);

	bfr new_net_1849_bfr_before (
		.din(new_net_1849),
		.dout(new_net_1848)
	);

	bfr new_net_1850_bfr_before (
		.din(new_net_1850),
		.dout(new_net_1849)
	);

	bfr new_net_1851_bfr_before (
		.din(new_net_1851),
		.dout(new_net_1850)
	);

	spl3L _0271__v_fanout (
		.a(_0271_),
		.b(new_net_887),
		.c(new_net_886),
		.d(new_net_1851)
	);

	spl2 _0370__v_fanout (
		.a(_0370_),
		.b(new_net_627),
		.c(new_net_626)
	);

	bfr new_net_1852_bfr_after (
		.din(_0411_),
		.dout(new_net_1852)
	);

	bfr new_net_1853_bfr_after (
		.din(new_net_1852),
		.dout(new_net_1853)
	);

	bfr new_net_1854_bfr_after (
		.din(new_net_1853),
		.dout(new_net_1854)
	);

	spl2 _0411__v_fanout (
		.a(new_net_1854),
		.b(new_net_559),
		.c(new_net_558)
	);

	bfr new_net_1855_bfr_after (
		.din(_0316_),
		.dout(new_net_1855)
	);

	bfr new_net_1856_bfr_after (
		.din(new_net_1855),
		.dout(new_net_1856)
	);

	bfr new_net_1857_bfr_after (
		.din(new_net_1856),
		.dout(new_net_1857)
	);

	spl2 _0316__v_fanout (
		.a(new_net_1857),
		.b(new_net_30),
		.c(new_net_29)
	);

	bfr new_net_1858_bfr_after (
		.din(_0310_),
		.dout(new_net_1858)
	);

	bfr new_net_1859_bfr_after (
		.din(new_net_1858),
		.dout(new_net_1859)
	);

	bfr new_net_1860_bfr_after (
		.din(new_net_1859),
		.dout(new_net_1860)
	);

	spl2 _0310__v_fanout (
		.a(new_net_1860),
		.b(new_net_762),
		.c(new_net_761)
	);

	spl2 _0430__v_fanout (
		.a(_0430_),
		.b(new_net_371),
		.c(new_net_370)
	);

	spl3L _0212__v_fanout (
		.a(_0212_),
		.b(new_net_50),
		.c(new_net_51),
		.d(new_net_49)
	);

	spl3L _0150__v_fanout (
		.a(_0150_),
		.b(new_net_12),
		.c(new_net_13),
		.d(new_net_11)
	);

	spl2 new_net_1239_v_fanout (
		.a(new_net_1239),
		.b(new_net_72),
		.c(new_net_70)
	);

	spl2 new_net_1238_v_fanout (
		.a(new_net_1238),
		.b(new_net_1047),
		.c(new_net_1045)
	);

	spl3L _0260__v_fanout (
		.a(_0260_),
		.b(new_net_366),
		.c(new_net_367),
		.d(new_net_365)
	);

	spl3L _0236__v_fanout (
		.a(_0236_),
		.b(new_net_109),
		.c(new_net_110),
		.d(new_net_108)
	);

	spl3L new_net_1222_v_fanout (
		.a(new_net_1222),
		.b(new_net_482),
		.c(new_net_477),
		.d(new_net_473)
	);

	bfr new_net_1861_bfr_before (
		.din(new_net_1861),
		.dout(new_net_1224)
	);

	bfr new_net_1862_bfr_before (
		.din(new_net_1862),
		.dout(new_net_1223)
	);

	spl4L new_net_1225_v_fanout (
		.a(new_net_1225),
		.b(new_net_476),
		.c(new_net_475),
		.d(new_net_1861),
		.e(new_net_1862)
	);

	spl3L _0183__v_fanout (
		.a(_0183_),
		.b(new_net_834),
		.c(new_net_835),
		.d(new_net_833)
	);

	spl2 new_net_1237_v_fanout (
		.a(new_net_1237),
		.b(new_net_535),
		.c(new_net_533)
	);

	spl4L _0223__v_fanout (
		.a(_0223_),
		.b(new_net_611),
		.c(new_net_612),
		.d(new_net_609),
		.e(new_net_610)
	);

	spl2 _0473__v_fanout (
		.a(_0473_),
		.b(new_net_488),
		.c(new_net_487)
	);

	spl4L new_net_1152_v_fanout (
		.a(new_net_1152),
		.b(new_net_1032),
		.c(new_net_1034),
		.d(new_net_1031),
		.e(new_net_1036)
	);

	spl2 _0100__v_fanout (
		.a(_0100_),
		.b(new_net_1237),
		.c(new_net_534)
	);

	spl3L _0245__v_fanout (
		.a(_0245_),
		.b(new_net_683),
		.c(new_net_684),
		.d(new_net_682)
	);

	spl3L new_net_1151_v_fanout (
		.a(new_net_1151),
		.b(new_net_1033),
		.c(new_net_1038),
		.d(new_net_1037)
	);

	spl2 _0160__v_fanout (
		.a(_0160_),
		.b(new_net_388),
		.c(new_net_387)
	);

	spl2 _0109__v_fanout (
		.a(_0109_),
		.b(new_net_1040),
		.c(new_net_1039)
	);

	spl2 new_net_1232_v_fanout (
		.a(new_net_1232),
		.b(new_net_695),
		.c(new_net_696)
	);

	spl2 _0126__v_fanout (
		.a(_0126_),
		.b(new_net_1046),
		.c(new_net_1238)
	);

	spl2 _0135__v_fanout (
		.a(_0135_),
		.b(new_net_392),
		.c(new_net_391)
	);

	spl4L new_net_1229_v_fanout (
		.a(new_net_1229),
		.b(new_net_571),
		.c(new_net_570),
		.d(new_net_568),
		.e(new_net_569)
	);

	spl3L _0269__v_fanout (
		.a(_0269_),
		.b(new_net_926),
		.c(new_net_927),
		.d(new_net_925)
	);

	spl4L new_net_1157_v_fanout (
		.a(new_net_1157),
		.b(new_net_144),
		.c(new_net_147),
		.d(new_net_142),
		.e(new_net_148)
	);

	bfr new_net_1863_bfr_after (
		.din(_0407_),
		.dout(new_net_1863)
	);

	bfr new_net_1864_bfr_after (
		.din(new_net_1863),
		.dout(new_net_1864)
	);

	bfr new_net_1865_bfr_after (
		.din(new_net_1864),
		.dout(new_net_1865)
	);

	bfr new_net_1866_bfr_after (
		.din(new_net_1865),
		.dout(new_net_1866)
	);

	spl2 _0407__v_fanout (
		.a(new_net_1866),
		.b(new_net_1235),
		.c(new_net_1236)
	);

	spl4L new_net_1230_v_fanout (
		.a(new_net_1230),
		.b(new_net_562),
		.c(new_net_563),
		.d(new_net_573),
		.e(new_net_572)
	);

	spl3L new_net_1156_v_fanout (
		.a(new_net_1156),
		.b(new_net_141),
		.c(new_net_140),
		.d(new_net_146)
	);

	spl4L new_net_1231_v_fanout (
		.a(new_net_1231),
		.b(new_net_566),
		.c(new_net_567),
		.d(new_net_564),
		.e(new_net_565)
	);

	spl2 _0065__v_fanout (
		.a(_0065_),
		.b(new_net_1239),
		.c(new_net_71)
	);

	spl2 _0082__v_fanout (
		.a(_0082_),
		.b(new_net_317),
		.c(new_net_316)
	);

	bfr new_net_1867_bfr_before (
		.din(new_net_1867),
		.dout(new_net_787)
	);

	bfr new_net_1868_bfr_before (
		.din(new_net_1868),
		.dout(new_net_1867)
	);

	spl2 _0395__v_fanout (
		.a(_0395_),
		.b(new_net_788),
		.c(new_net_1868)
	);

	spl2 _0442__v_fanout (
		.a(_0442_),
		.b(new_net_1232),
		.c(new_net_694)
	);

	spl3L _0369__v_fanout (
		.a(_0369_),
		.b(new_net_1230),
		.c(new_net_1229),
		.d(new_net_1231)
	);

	spl2 _0524__v_fanout (
		.a(_0524_),
		.b(new_net_934),
		.c(new_net_933)
	);

	spl4L _0072__v_fanout (
		.a(_0072_),
		.b(new_net_430),
		.c(new_net_428),
		.d(new_net_427),
		.e(new_net_429)
	);

	spl3L _0214__v_fanout (
		.a(_0214_),
		.b(new_net_590),
		.c(new_net_589),
		.d(new_net_588)
	);

	spl2 _0375__v_fanout (
		.a(_0375_),
		.b(new_net_866),
		.c(new_net_865)
	);

	spl2 _0436__v_fanout (
		.a(_0436_),
		.b(new_net_809),
		.c(new_net_808)
	);

	spl2 _0244__v_fanout (
		.a(_0244_),
		.b(new_net_625),
		.c(new_net_624)
	);

	bfr new_net_1869_bfr_after (
		.din(_0337_),
		.dout(new_net_1869)
	);

	bfr new_net_1870_bfr_after (
		.din(new_net_1869),
		.dout(new_net_1870)
	);

	bfr new_net_1871_bfr_after (
		.din(new_net_1870),
		.dout(new_net_1871)
	);

	bfr new_net_1872_bfr_after (
		.din(new_net_1871),
		.dout(new_net_1872)
	);

	bfr new_net_1873_bfr_after (
		.din(new_net_1872),
		.dout(new_net_1873)
	);

	bfr new_net_1874_bfr_after (
		.din(new_net_1873),
		.dout(new_net_1874)
	);

	bfr new_net_1875_bfr_after (
		.din(new_net_1874),
		.dout(new_net_1875)
	);

	bfr new_net_1876_bfr_after (
		.din(new_net_1875),
		.dout(new_net_1876)
	);

	bfr new_net_1877_bfr_after (
		.din(new_net_1876),
		.dout(new_net_1877)
	);

	bfr new_net_1878_bfr_after (
		.din(new_net_1877),
		.dout(new_net_1878)
	);

	bfr new_net_1879_bfr_after (
		.din(new_net_1878),
		.dout(new_net_1879)
	);

	bfr new_net_1880_bfr_after (
		.din(new_net_1879),
		.dout(new_net_1880)
	);

	bfr new_net_1881_bfr_after (
		.din(new_net_1880),
		.dout(new_net_1881)
	);

	bfr new_net_1882_bfr_after (
		.din(new_net_1881),
		.dout(new_net_1882)
	);

	bfr new_net_1883_bfr_after (
		.din(new_net_1882),
		.dout(new_net_1883)
	);

	bfr new_net_1884_bfr_after (
		.din(new_net_1883),
		.dout(new_net_1884)
	);

	bfr new_net_1885_bfr_after (
		.din(new_net_1884),
		.dout(new_net_1885)
	);

	bfr new_net_1886_bfr_after (
		.din(new_net_1885),
		.dout(new_net_1886)
	);

	spl2 _0337__v_fanout (
		.a(new_net_1886),
		.b(new_net_1226),
		.c(new_net_24)
	);

	spl2 _0268__v_fanout (
		.a(_0268_),
		.b(new_net_760),
		.c(new_net_759)
	);

	spl2 _0142__v_fanout (
		.a(_0142_),
		.b(new_net_764),
		.c(new_net_763)
	);

	bfr new_net_1887_bfr_before (
		.din(new_net_1887),
		.dout(new_net_268)
	);

	bfr new_net_1888_bfr_before (
		.din(new_net_1888),
		.dout(new_net_1887)
	);

	bfr new_net_1889_bfr_before (
		.din(new_net_1889),
		.dout(new_net_1888)
	);

	bfr new_net_1890_bfr_before (
		.din(new_net_1890),
		.dout(new_net_1889)
	);

	spl2 _0384__v_fanout (
		.a(_0384_),
		.b(new_net_1890),
		.c(new_net_267)
	);

	spl4L _0195__v_fanout (
		.a(_0195_),
		.b(new_net_101),
		.c(new_net_102),
		.d(new_net_99),
		.e(new_net_100)
	);

	bfr new_net_1891_bfr_before (
		.din(new_net_1891),
		.dout(new_net_1221)
	);

	bfr new_net_1892_bfr_before (
		.din(new_net_1892),
		.dout(new_net_1891)
	);

	bfr new_net_1893_bfr_before (
		.din(new_net_1893),
		.dout(new_net_1892)
	);

	bfr new_net_1894_bfr_before (
		.din(new_net_1894),
		.dout(new_net_1893)
	);

	bfr new_net_1895_bfr_before (
		.din(new_net_1895),
		.dout(new_net_1894)
	);

	bfr new_net_1896_bfr_before (
		.din(new_net_1896),
		.dout(new_net_1895)
	);

	bfr new_net_1897_bfr_before (
		.din(new_net_1897),
		.dout(new_net_1896)
	);

	bfr new_net_1898_bfr_before (
		.din(new_net_1898),
		.dout(new_net_1897)
	);

	bfr new_net_1899_bfr_before (
		.din(new_net_1899),
		.dout(new_net_1898)
	);

	bfr new_net_1900_bfr_before (
		.din(new_net_1900),
		.dout(new_net_1899)
	);

	spl2 _0406__v_fanout (
		.a(_0406_),
		.b(new_net_1900),
		.c(new_net_342)
	);

	bfr new_net_1901_bfr_after (
		.din(_0287_),
		.dout(new_net_1901)
	);

	bfr new_net_1902_bfr_after (
		.din(new_net_1901),
		.dout(new_net_1902)
	);

	spl3L _0287__v_fanout (
		.a(new_net_1902),
		.b(new_net_1222),
		.c(new_net_1225),
		.d(new_net_472)
	);

	bfr new_net_1903_bfr_before (
		.din(new_net_1903),
		.dout(new_net_1157)
	);

	bfr new_net_1904_bfr_before (
		.din(new_net_1904),
		.dout(new_net_1156)
	);

	spl3L new_net_1155_v_fanout (
		.a(new_net_1155),
		.b(new_net_145),
		.c(new_net_1904),
		.d(new_net_1903)
	);

	spl4L new_net_1212_v_fanout (
		.a(new_net_1212),
		.b(new_net_512),
		.c(new_net_511),
		.d(new_net_509),
		.e(new_net_513)
	);

	spl4L new_net_1199_v_fanout (
		.a(new_net_1199),
		.b(new_net_298),
		.c(new_net_308),
		.d(new_net_312),
		.e(new_net_310)
	);

	spl3L new_net_1198_v_fanout (
		.a(new_net_1198),
		.b(new_net_315),
		.c(new_net_301),
		.d(new_net_305)
	);

	bfr new_net_1905_bfr_before (
		.din(new_net_1905),
		.dout(new_net_914)
	);

	bfr new_net_1906_bfr_before (
		.din(new_net_1906),
		.dout(new_net_1905)
	);

	spl2 new_net_1154_v_fanout (
		.a(new_net_1154),
		.b(new_net_1906),
		.c(new_net_911)
	);

	spl3L new_net_1193_v_fanout (
		.a(new_net_1193),
		.b(new_net_398),
		.c(new_net_400),
		.d(new_net_394)
	);

	spl4L new_net_1202_v_fanout (
		.a(new_net_1202),
		.b(new_net_299),
		.c(new_net_311),
		.d(new_net_307),
		.e(new_net_309)
	);

	spl4L new_net_1210_v_fanout (
		.a(new_net_1210),
		.b(new_net_517),
		.c(new_net_518),
		.d(new_net_520),
		.e(new_net_522)
	);

	spl4L new_net_1201_v_fanout (
		.a(new_net_1201),
		.b(new_net_297),
		.c(new_net_313),
		.d(new_net_314),
		.e(new_net_303)
	);

	spl3L new_net_1213_v_fanout (
		.a(new_net_1213),
		.b(new_net_516),
		.c(new_net_515),
		.d(new_net_514)
	);

	spl2 _0033__v_fanout (
		.a(_0033_),
		.b(new_net_273),
		.c(new_net_272)
	);

	spl2 new_net_1209_v_fanout (
		.a(new_net_1209),
		.b(new_net_521),
		.c(new_net_519)
	);

	spl4L _0179__v_fanout (
		.a(_0179_),
		.b(new_net_484),
		.c(new_net_485),
		.d(new_net_483),
		.e(new_net_486)
	);

	bfr new_net_1907_bfr_before (
		.din(new_net_1907),
		.dout(new_net_505)
	);

	bfr new_net_1908_bfr_before (
		.din(new_net_1908),
		.dout(new_net_1907)
	);

	bfr new_net_1909_bfr_before (
		.din(new_net_1909),
		.dout(new_net_1908)
	);

	spl2 new_net_1170_v_fanout (
		.a(new_net_1170),
		.b(new_net_1909),
		.c(new_net_502)
	);

	spl4L new_net_1200_v_fanout (
		.a(new_net_1200),
		.b(new_net_304),
		.c(new_net_302),
		.d(new_net_300),
		.e(new_net_306)
	);

	spl4L new_net_1211_v_fanout (
		.a(new_net_1211),
		.b(new_net_508),
		.c(new_net_507),
		.d(new_net_506),
		.e(new_net_510)
	);

	spl2 new_net_1119_v_fanout (
		.a(new_net_1119),
		.b(new_net_422),
		.c(new_net_420)
	);

	bfr new_net_1910_bfr_before (
		.din(new_net_1910),
		.dout(new_net_180)
	);

	bfr new_net_1911_bfr_before (
		.din(new_net_1911),
		.dout(new_net_171)
	);

	bfr new_net_1912_bfr_before (
		.din(new_net_1912),
		.dout(new_net_1911)
	);

	bfr new_net_1913_bfr_before (
		.din(new_net_1913),
		.dout(new_net_1912)
	);

	bfr new_net_1914_bfr_before (
		.din(new_net_1914),
		.dout(new_net_1913)
	);

	bfr new_net_1915_bfr_before (
		.din(new_net_1915),
		.dout(new_net_1914)
	);

	bfr new_net_1916_bfr_before (
		.din(new_net_1916),
		.dout(new_net_154)
	);

	spl4L new_net_1092_v_fanout (
		.a(new_net_1092),
		.b(new_net_1916),
		.c(new_net_1915),
		.d(new_net_167),
		.e(new_net_1910)
	);

	bfr new_net_1917_bfr_after (
		.din(_0513_),
		.dout(new_net_1917)
	);

	bfr new_net_1918_bfr_before (
		.din(new_net_1918),
		.dout(new_net_780)
	);

	bfr new_net_1919_bfr_before (
		.din(new_net_1919),
		.dout(new_net_1918)
	);

	spl2 _0513__v_fanout (
		.a(new_net_1917),
		.b(new_net_1919),
		.c(new_net_779)
	);

	bfr new_net_1920_bfr_before (
		.din(new_net_1920),
		.dout(new_net_577)
	);

	spl4L _0117__v_fanout (
		.a(_0117_),
		.b(new_net_575),
		.c(new_net_576),
		.d(new_net_574),
		.e(new_net_1920)
	);

	bfr new_net_1921_bfr_after (
		.din(_0575_),
		.dout(new_net_1921)
	);

	bfr new_net_1922_bfr_after (
		.din(new_net_1921),
		.dout(new_net_1922)
	);

	bfr new_net_1923_bfr_after (
		.din(new_net_1922),
		.dout(new_net_1923)
	);

	bfr new_net_1924_bfr_after (
		.din(new_net_1923),
		.dout(new_net_1924)
	);

	bfr new_net_1925_bfr_after (
		.din(new_net_1924),
		.dout(new_net_1925)
	);

	bfr new_net_1926_bfr_after (
		.din(new_net_1925),
		.dout(new_net_1926)
	);

	bfr new_net_1927_bfr_after (
		.din(new_net_1926),
		.dout(new_net_1927)
	);

	bfr new_net_1928_bfr_after (
		.din(new_net_1927),
		.dout(new_net_1928)
	);

	bfr new_net_1929_bfr_after (
		.din(new_net_1928),
		.dout(new_net_1929)
	);

	bfr new_net_1930_bfr_after (
		.din(new_net_1929),
		.dout(new_net_1930)
	);

	bfr new_net_1931_bfr_after (
		.din(new_net_1930),
		.dout(new_net_1931)
	);

	bfr new_net_1932_bfr_after (
		.din(new_net_1931),
		.dout(new_net_1932)
	);

	spl4L _0575__v_fanout (
		.a(new_net_1932),
		.b(new_net_223),
		.c(new_net_225),
		.d(new_net_222),
		.e(new_net_224)
	);

	spl2 new_net_1214_v_fanout (
		.a(new_net_1214),
		.b(new_net_1209),
		.c(new_net_1210)
	);

	spl4L new_net_1216_v_fanout (
		.a(new_net_1216),
		.b(new_net_737),
		.c(new_net_745),
		.d(new_net_735),
		.e(new_net_736)
	);

	spl2 _0071__v_fanout (
		.a(_0071_),
		.b(new_net_724),
		.c(new_net_723)
	);

	bfr new_net_1933_bfr_before (
		.din(new_net_1933),
		.dout(new_net_192)
	);

	bfr new_net_1934_bfr_before (
		.din(new_net_1934),
		.dout(new_net_1933)
	);

	bfr new_net_1935_bfr_before (
		.din(new_net_1935),
		.dout(new_net_1934)
	);

	spl2 new_net_1160_v_fanout (
		.a(new_net_1160),
		.b(new_net_1935),
		.c(new_net_190)
	);

	spl3L new_net_1204_v_fanout (
		.a(new_net_1204),
		.b(new_net_1201),
		.c(new_net_1200),
		.d(new_net_1198)
	);

	bfr new_net_1936_bfr_before (
		.din(new_net_1936),
		.dout(new_net_798)
	);

	bfr new_net_1937_bfr_before (
		.din(new_net_1937),
		.dout(new_net_1936)
	);

	bfr new_net_1938_bfr_before (
		.din(new_net_1938),
		.dout(new_net_1937)
	);

	bfr new_net_1939_bfr_before (
		.din(new_net_1939),
		.dout(new_net_1938)
	);

	spl2 new_net_1149_v_fanout (
		.a(new_net_1149),
		.b(new_net_802),
		.c(new_net_1939)
	);

	spl4L new_net_1208_v_fanout (
		.a(new_net_1208),
		.b(new_net_821),
		.c(new_net_820),
		.d(new_net_818),
		.e(new_net_822)
	);

	spl4L new_net_1189_v_fanout (
		.a(new_net_1189),
		.b(new_net_337),
		.c(new_net_336),
		.d(new_net_334),
		.e(new_net_335)
	);

	bfr new_net_1940_bfr_after (
		.din(_0315_),
		.dout(new_net_1940)
	);

	bfr new_net_1941_bfr_after (
		.din(new_net_1940),
		.dout(new_net_1941)
	);

	bfr new_net_1942_bfr_after (
		.din(new_net_1941),
		.dout(new_net_1942)
	);

	bfr new_net_1943_bfr_after (
		.din(new_net_1942),
		.dout(new_net_1943)
	);

	bfr new_net_1944_bfr_before (
		.din(new_net_1944),
		.dout(new_net_990)
	);

	bfr new_net_1945_bfr_before (
		.din(new_net_1945),
		.dout(new_net_1944)
	);

	bfr new_net_1946_bfr_before (
		.din(new_net_1946),
		.dout(new_net_1945)
	);

	spl3L _0315__v_fanout (
		.a(new_net_1943),
		.b(new_net_991),
		.c(new_net_1946),
		.d(new_net_989)
	);

	spl4L new_net_1217_v_fanout (
		.a(new_net_1217),
		.b(new_net_739),
		.c(new_net_740),
		.d(new_net_738),
		.e(new_net_741)
	);

	spl4L new_net_1206_v_fanout (
		.a(new_net_1206),
		.b(new_net_827),
		.c(new_net_829),
		.d(new_net_830),
		.e(new_net_826)
	);

	spl4L new_net_1205_v_fanout (
		.a(new_net_1205),
		.b(new_net_828),
		.c(new_net_825),
		.d(new_net_823),
		.e(new_net_824)
	);

	spl3L _0336__v_fanout (
		.a(_0336_),
		.b(new_net_1011),
		.c(new_net_1012),
		.d(new_net_1010)
	);

	bfr new_net_1947_bfr_before (
		.din(new_net_1947),
		.dout(new_net_904)
	);

	bfr new_net_1948_bfr_before (
		.din(new_net_1948),
		.dout(new_net_1947)
	);

	bfr new_net_1949_bfr_before (
		.din(new_net_1949),
		.dout(new_net_1948)
	);

	bfr new_net_1950_bfr_before (
		.din(new_net_1950),
		.dout(new_net_1949)
	);

	spl2 new_net_1165_v_fanout (
		.a(new_net_1165),
		.b(new_net_907),
		.c(new_net_1950)
	);

	spl4L new_net_1190_v_fanout (
		.a(new_net_1190),
		.b(new_net_330),
		.c(new_net_331),
		.d(new_net_329),
		.e(new_net_333)
	);

	spl2 new_net_1203_v_fanout (
		.a(new_net_1203),
		.b(new_net_1199),
		.c(new_net_1202)
	);

	bfr new_net_1951_bfr_before (
		.din(new_net_1951),
		.dout(new_net_202)
	);

	spl2 new_net_1174_v_fanout (
		.a(new_net_1174),
		.b(new_net_1951),
		.c(new_net_197)
	);

	bfr new_net_1952_bfr_after (
		.din(_0378_),
		.dout(new_net_1952)
	);

	bfr new_net_1953_bfr_before (
		.din(new_net_1953),
		.dout(new_net_781)
	);

	spl2 _0378__v_fanout (
		.a(new_net_1952),
		.b(new_net_782),
		.c(new_net_1953)
	);

	bfr new_net_1954_bfr_before (
		.din(new_net_1954),
		.dout(new_net_600)
	);

	spl2 new_net_1080_v_fanout (
		.a(new_net_1080),
		.b(new_net_1954),
		.c(new_net_593)
	);

	bfr new_net_1955_bfr_after (
		.din(_0432_),
		.dout(new_net_1955)
	);

	bfr new_net_1956_bfr_after (
		.din(new_net_1955),
		.dout(new_net_1956)
	);

	bfr new_net_1957_bfr_before (
		.din(new_net_1957),
		.dout(new_net_548)
	);

	bfr new_net_1958_bfr_before (
		.din(new_net_1958),
		.dout(new_net_1957)
	);

	bfr new_net_1959_bfr_before (
		.din(new_net_1959),
		.dout(new_net_1958)
	);

	spl2 _0432__v_fanout (
		.a(new_net_1956),
		.b(new_net_1959),
		.c(new_net_547)
	);

	spl3L new_net_1192_v_fanout (
		.a(new_net_1192),
		.b(new_net_1193),
		.c(new_net_396),
		.d(new_net_399)
	);

	spl4L _0052__v_fanout (
		.a(_0052_),
		.b(new_net_448),
		.c(new_net_449),
		.d(new_net_447),
		.e(new_net_450)
	);

	bfr new_net_1960_bfr_after (
		.din(_0481_),
		.dout(new_net_1960)
	);

	bfr new_net_1961_bfr_before (
		.din(new_net_1961),
		.dout(new_net_882)
	);

	bfr new_net_1962_bfr_before (
		.din(new_net_1962),
		.dout(new_net_1961)
	);

	bfr new_net_1963_bfr_before (
		.din(new_net_1963),
		.dout(new_net_1962)
	);

	spl2 _0481__v_fanout (
		.a(new_net_1960),
		.b(new_net_1963),
		.c(new_net_881)
	);

	spl4L new_net_1207_v_fanout (
		.a(new_net_1207),
		.b(new_net_817),
		.c(new_net_819),
		.d(new_net_815),
		.e(new_net_816)
	);

	bfr new_net_1964_bfr_before (
		.din(new_net_1964),
		.dout(new_net_1220)
	);

	bfr new_net_1965_bfr_before (
		.din(new_net_1965),
		.dout(new_net_1964)
	);

	bfr new_net_1966_bfr_before (
		.din(new_net_1966),
		.dout(new_net_1965)
	);

	bfr new_net_1967_bfr_before (
		.din(new_net_1967),
		.dout(new_net_1966)
	);

	bfr new_net_1968_bfr_before (
		.din(new_net_1968),
		.dout(new_net_1967)
	);

	bfr new_net_1969_bfr_before (
		.din(new_net_1969),
		.dout(new_net_1968)
	);

	spl2 _0286__v_fanout (
		.a(_0286_),
		.b(new_net_1969),
		.c(new_net_628)
	);

	spl3L new_net_1215_v_fanout (
		.a(new_net_1215),
		.b(new_net_1213),
		.c(new_net_1212),
		.d(new_net_1211)
	);

	spl4L new_net_1219_v_fanout (
		.a(new_net_1219),
		.b(new_net_732),
		.c(new_net_734),
		.d(new_net_730),
		.e(new_net_731)
	);

	spl4L new_net_1218_v_fanout (
		.a(new_net_1218),
		.b(new_net_743),
		.c(new_net_733),
		.d(new_net_742),
		.e(new_net_744)
	);

	bfr new_net_1970_bfr_before (
		.din(new_net_1970),
		.dout(new_net_196)
	);

	bfr new_net_1971_bfr_before (
		.din(new_net_1971),
		.dout(new_net_200)
	);

	spl3L new_net_1175_v_fanout (
		.a(new_net_1175),
		.b(new_net_199),
		.c(new_net_1971),
		.d(new_net_1970)
	);

	spl4L _0374__v_fanout (
		.a(_0374_),
		.b(new_net_1207),
		.c(new_net_1205),
		.d(new_net_1206),
		.e(new_net_1208)
	);

	bfr new_net_1972_bfr_before (
		.din(new_net_1972),
		.dout(new_net_799)
	);

	bfr new_net_1973_bfr_before (
		.din(new_net_1973),
		.dout(new_net_803)
	);

	bfr new_net_1974_bfr_before (
		.din(new_net_1974),
		.dout(new_net_1973)
	);

	bfr new_net_1975_bfr_before (
		.din(new_net_1975),
		.dout(new_net_797)
	);

	spl4L new_net_1148_v_fanout (
		.a(new_net_1148),
		.b(new_net_1149),
		.c(new_net_1975),
		.d(new_net_1972),
		.e(new_net_1974)
	);

	bfr new_net_1976_bfr_before (
		.din(new_net_1976),
		.dout(new_net_504)
	);

	spl2 new_net_1169_v_fanout (
		.a(new_net_1169),
		.b(new_net_1170),
		.c(new_net_1976)
	);

	bfr new_net_1977_bfr_after (
		.din(_0042_),
		.dout(new_net_1977)
	);

	bfr new_net_1978_bfr_after (
		.din(new_net_1977),
		.dout(new_net_1978)
	);

	spl2 _0042__v_fanout (
		.a(new_net_1978),
		.b(new_net_1021),
		.c(new_net_1020)
	);

	bfr new_net_1979_bfr_before (
		.din(new_net_1979),
		.dout(new_net_720)
	);

	bfr new_net_1980_bfr_before (
		.din(new_net_1980),
		.dout(new_net_1979)
	);

	bfr new_net_1981_bfr_before (
		.din(new_net_1981),
		.dout(new_net_1980)
	);

	spl2 new_net_1168_v_fanout (
		.a(new_net_1168),
		.b(new_net_1981),
		.c(new_net_719)
	);

	spl2 new_net_1130_v_fanout (
		.a(new_net_1130),
		.b(new_net_464),
		.c(new_net_462)
	);

	bfr new_net_1982_bfr_before (
		.din(new_net_1982),
		.dout(new_net_974)
	);

	bfr new_net_1983_bfr_before (
		.din(new_net_1983),
		.dout(new_net_1982)
	);

	bfr new_net_1984_bfr_before (
		.din(new_net_1984),
		.dout(new_net_1983)
	);

	bfr new_net_1985_bfr_before (
		.din(new_net_1985),
		.dout(new_net_1984)
	);

	spl3L new_net_1166_v_fanout (
		.a(new_net_1166),
		.b(new_net_1985),
		.c(new_net_973),
		.d(new_net_971)
	);

	bfr new_net_1986_bfr_before (
		.din(new_net_1986),
		.dout(new_net_671)
	);

	bfr new_net_1987_bfr_before (
		.din(new_net_1987),
		.dout(new_net_672)
	);

	spl3L new_net_1127_v_fanout (
		.a(new_net_1127),
		.b(new_net_1987),
		.c(new_net_676),
		.d(new_net_1986)
	);

	bfr new_net_1988_bfr_before (
		.din(new_net_1988),
		.dout(new_net_852)
	);

	spl2 new_net_1111_v_fanout (
		.a(new_net_1111),
		.b(new_net_853),
		.c(new_net_1988)
	);

	spl4L _0372__v_fanout (
		.a(_0372_),
		.b(new_net_1217),
		.c(new_net_1216),
		.d(new_net_1218),
		.e(new_net_1219)
	);

	bfr new_net_1989_bfr_before (
		.din(new_net_1989),
		.dout(new_net_906)
	);

	bfr new_net_1990_bfr_before (
		.din(new_net_1990),
		.dout(new_net_905)
	);

	bfr new_net_1991_bfr_before (
		.din(new_net_1991),
		.dout(new_net_1990)
	);

	spl3L new_net_1164_v_fanout (
		.a(new_net_1164),
		.b(new_net_1991),
		.c(new_net_1165),
		.d(new_net_1989)
	);

	bfr new_net_1992_bfr_after (
		.din(_0334_),
		.dout(new_net_1992)
	);

	bfr new_net_1993_bfr_after (
		.din(new_net_1992),
		.dout(new_net_1993)
	);

	bfr new_net_1994_bfr_after (
		.din(new_net_1993),
		.dout(new_net_1994)
	);

	bfr new_net_1995_bfr_after (
		.din(new_net_1994),
		.dout(new_net_1995)
	);

	bfr new_net_1996_bfr_after (
		.din(new_net_1995),
		.dout(new_net_1996)
	);

	bfr new_net_1997_bfr_after (
		.din(new_net_1996),
		.dout(new_net_1997)
	);

	bfr new_net_1998_bfr_after (
		.din(new_net_1997),
		.dout(new_net_1998)
	);

	bfr new_net_1999_bfr_after (
		.din(new_net_1998),
		.dout(new_net_1999)
	);

	bfr new_net_2000_bfr_after (
		.din(new_net_1999),
		.dout(new_net_2000)
	);

	bfr new_net_2001_bfr_after (
		.din(new_net_2000),
		.dout(new_net_2001)
	);

	bfr new_net_2002_bfr_after (
		.din(new_net_2001),
		.dout(new_net_2002)
	);

	bfr new_net_2003_bfr_after (
		.din(new_net_2002),
		.dout(new_net_2003)
	);

	bfr new_net_2004_bfr_after (
		.din(new_net_2003),
		.dout(new_net_2004)
	);

	bfr new_net_2005_bfr_after (
		.din(new_net_2004),
		.dout(new_net_2005)
	);

	bfr new_net_2006_bfr_after (
		.din(new_net_2005),
		.dout(new_net_2006)
	);

	bfr new_net_2007_bfr_after (
		.din(new_net_2006),
		.dout(new_net_2007)
	);

	bfr new_net_2008_bfr_after (
		.din(new_net_2007),
		.dout(new_net_2008)
	);

	bfr new_net_2009_bfr_after (
		.din(new_net_2008),
		.dout(new_net_2009)
	);

	bfr new_net_2010_bfr_after (
		.din(new_net_2009),
		.dout(new_net_2010)
	);

	bfr new_net_2011_bfr_after (
		.din(new_net_2010),
		.dout(new_net_2011)
	);

	bfr new_net_2012_bfr_before (
		.din(new_net_2012),
		.dout(new_net_1194)
	);

	bfr new_net_2013_bfr_before (
		.din(new_net_2013),
		.dout(new_net_2012)
	);

	spl2 _0334__v_fanout (
		.a(new_net_2011),
		.b(new_net_2013),
		.c(new_net_924)
	);

	spl2 _0363__v_fanout (
		.a(_0363_),
		.b(new_net_1204),
		.c(new_net_1203)
	);

	bfr new_net_2014_bfr_before (
		.din(new_net_2014),
		.dout(new_net_385)
	);

	bfr new_net_2015_bfr_before (
		.din(new_net_2015),
		.dout(new_net_2014)
	);

	bfr new_net_2016_bfr_before (
		.din(new_net_2016),
		.dout(new_net_2015)
	);

	bfr new_net_2017_bfr_before (
		.din(new_net_2017),
		.dout(new_net_2016)
	);

	bfr new_net_2018_bfr_before (
		.din(new_net_2018),
		.dout(new_net_382)
	);

	spl3L new_net_1142_v_fanout (
		.a(new_net_1142),
		.b(new_net_383),
		.c(new_net_2018),
		.d(new_net_2017)
	);

	bfr new_net_2019_bfr_before (
		.din(new_net_2019),
		.dout(new_net_1154)
	);

	bfr new_net_2020_bfr_before (
		.din(new_net_2020),
		.dout(new_net_909)
	);

	spl3L new_net_1153_v_fanout (
		.a(new_net_1153),
		.b(new_net_2020),
		.c(new_net_913),
		.d(new_net_2019)
	);

	spl2 new_net_1070_v_fanout (
		.a(new_net_1070),
		.b(new_net_288),
		.c(new_net_286)
	);

	bfr new_net_2021_bfr_before (
		.din(new_net_2021),
		.dout(new_net_461)
	);

	bfr new_net_2022_bfr_before (
		.din(new_net_2022),
		.dout(new_net_2021)
	);

	bfr new_net_2023_bfr_before (
		.din(new_net_2023),
		.dout(new_net_2022)
	);

	spl3L new_net_1131_v_fanout (
		.a(new_net_1131),
		.b(new_net_460),
		.c(new_net_2023),
		.d(new_net_463)
	);

	spl2 new_net_1159_v_fanout (
		.a(new_net_1159),
		.b(new_net_189),
		.c(new_net_1160)
	);

	spl2 _0023__v_fanout (
		.a(_0023_),
		.b(new_net_90),
		.c(new_net_89)
	);

	spl2 new_net_1191_v_fanout (
		.a(new_net_1191),
		.b(new_net_1192),
		.c(new_net_397)
	);

	bfr new_net_2024_bfr_before (
		.din(new_net_2024),
		.dout(new_net_444)
	);

	spl2 new_net_1121_v_fanout (
		.a(new_net_1121),
		.b(new_net_442),
		.c(new_net_2024)
	);

	spl2 _0014__v_fanout (
		.a(_0014_),
		.b(new_net_713),
		.c(new_net_712)
	);

	spl2 _0368__v_fanout (
		.a(_0368_),
		.b(new_net_1214),
		.c(new_net_1215)
	);

	spl4L new_net_1181_v_fanout (
		.a(new_net_1181),
		.b(new_net_654),
		.c(new_net_656),
		.d(new_net_652),
		.e(new_net_653)
	);

	spl4L new_net_1188_v_fanout (
		.a(new_net_1188),
		.b(new_net_960),
		.c(new_net_957),
		.d(new_net_959),
		.e(new_net_961)
	);

	bfr new_net_2025_bfr_before (
		.din(new_net_2025),
		.dout(new_net_634)
	);

	spl2 new_net_1058_v_fanout (
		.a(new_net_1058),
		.b(new_net_636),
		.c(new_net_2025)
	);

	bfr new_net_2026_bfr_before (
		.din(new_net_2026),
		.dout(new_net_756)
	);

	spl2 new_net_1089_v_fanout (
		.a(new_net_1089),
		.b(new_net_2026),
		.c(new_net_757)
	);

	spl4L _0000__v_fanout (
		.a(_0000_),
		.b(new_net_1018),
		.c(new_net_1019),
		.d(new_net_1016),
		.e(new_net_1017)
	);

	spl4L new_net_1184_v_fanout (
		.a(new_net_1184),
		.b(new_net_95),
		.c(new_net_93),
		.d(new_net_91),
		.e(new_net_92)
	);

	bfr new_net_2027_bfr_before (
		.din(new_net_2027),
		.dout(new_net_62)
	);

	spl2 new_net_1102_v_fanout (
		.a(new_net_1102),
		.b(new_net_63),
		.c(new_net_2027)
	);

	bfr new_net_2028_bfr_before (
		.din(new_net_2028),
		.dout(new_net_1174)
	);

	bfr new_net_2029_bfr_before (
		.din(new_net_2029),
		.dout(new_net_1175)
	);

	spl3L new_net_1173_v_fanout (
		.a(new_net_1173),
		.b(new_net_2029),
		.c(new_net_2028),
		.d(new_net_201)
	);

	spl3L _0051__v_fanout (
		.a(_0051_),
		.b(new_net_1191),
		.c(new_net_395),
		.d(new_net_393)
	);

	bfr new_net_2030_bfr_before (
		.din(new_net_2030),
		.dout(new_net_690)
	);

	bfr new_net_2031_bfr_before (
		.din(new_net_2031),
		.dout(new_net_2030)
	);

	bfr new_net_2032_bfr_before (
		.din(new_net_2032),
		.dout(new_net_2031)
	);

	spl2 new_net_1163_v_fanout (
		.a(new_net_1163),
		.b(new_net_687),
		.c(new_net_2032)
	);

	spl2 _0030__v_fanout (
		.a(_0030_),
		.b(new_net_553),
		.c(new_net_552)
	);

	spl4L new_net_1187_v_fanout (
		.a(new_net_1187),
		.b(new_net_967),
		.c(new_net_956),
		.d(new_net_966),
		.e(new_net_958)
	);

	bfr new_net_2033_bfr_before (
		.din(new_net_2033),
		.dout(new_net_541)
	);

	bfr new_net_2034_bfr_before (
		.din(new_net_2034),
		.dout(new_net_538)
	);

	bfr new_net_2035_bfr_before (
		.din(new_net_2035),
		.dout(new_net_2034)
	);

	bfr new_net_2036_bfr_before (
		.din(new_net_2036),
		.dout(new_net_2035)
	);

	bfr new_net_2037_bfr_before (
		.din(new_net_2037),
		.dout(new_net_2036)
	);

	spl3L new_net_1074_v_fanout (
		.a(new_net_1074),
		.b(new_net_2037),
		.c(new_net_2033),
		.d(new_net_540)
	);

	bfr new_net_2038_bfr_before (
		.din(new_net_2038),
		.dout(new_net_458)
	);

	bfr new_net_2039_bfr_before (
		.din(new_net_2039),
		.dout(new_net_2038)
	);

	spl2 _0205__v_fanout (
		.a(_0205_),
		.b(new_net_459),
		.c(new_net_2039)
	);

	spl2 new_net_1180_v_fanout (
		.a(new_net_1180),
		.b(new_net_657),
		.c(new_net_655)
	);

	bfr new_net_2040_bfr_before (
		.din(new_net_2040),
		.dout(new_net_402)
	);

	spl2 new_net_1061_v_fanout (
		.a(new_net_1061),
		.b(new_net_2040),
		.c(new_net_401)
	);

	bfr new_net_2041_bfr_before (
		.din(new_net_2041),
		.dout(new_net_615)
	);

	bfr new_net_2042_bfr_before (
		.din(new_net_2042),
		.dout(new_net_2041)
	);

	bfr new_net_2043_bfr_before (
		.din(new_net_2043),
		.dout(new_net_2042)
	);

	bfr new_net_2044_bfr_before (
		.din(new_net_2044),
		.dout(new_net_2043)
	);

	bfr new_net_2045_bfr_before (
		.din(new_net_2045),
		.dout(new_net_616)
	);

	bfr new_net_2046_bfr_before (
		.din(new_net_2046),
		.dout(new_net_618)
	);

	spl4L new_net_1057_v_fanout (
		.a(new_net_1057),
		.b(new_net_619),
		.c(new_net_2046),
		.d(new_net_2044),
		.e(new_net_2045)
	);

	spl3L new_net_1185_v_fanout (
		.a(new_net_1185),
		.b(new_net_277),
		.c(new_net_275),
		.d(new_net_274)
	);

	spl4L new_net_1186_v_fanout (
		.a(new_net_1186),
		.b(new_net_964),
		.c(new_net_965),
		.d(new_net_962),
		.e(new_net_963)
	);

	spl4L new_net_1183_v_fanout (
		.a(new_net_1183),
		.b(new_net_98),
		.c(new_net_97),
		.d(new_net_94),
		.e(new_net_96)
	);

	spl2 new_net_1182_v_fanout (
		.a(new_net_1182),
		.b(new_net_951),
		.c(new_net_950)
	);

	bfr new_net_2047_bfr_before (
		.din(new_net_2047),
		.dout(new_net_1190)
	);

	bfr new_net_2048_bfr_before (
		.din(new_net_2048),
		.dout(new_net_1189)
	);

	spl3L _0070__v_fanout (
		.a(_0070_),
		.b(new_net_2048),
		.c(new_net_2047),
		.d(new_net_332)
	);

	spl4L new_net_1176_v_fanout (
		.a(new_net_1176),
		.b(new_net_417),
		.c(new_net_416),
		.d(new_net_412),
		.e(new_net_415)
	);

	bfr new_net_2049_bfr_before (
		.din(new_net_2049),
		.dout(new_net_1127)
	);

	spl2 new_net_1126_v_fanout (
		.a(new_net_1126),
		.b(new_net_675),
		.c(new_net_2049)
	);

	bfr new_net_2050_bfr_before (
		.din(new_net_2050),
		.dout(new_net_524)
	);

	bfr new_net_2051_bfr_before (
		.din(new_net_2051),
		.dout(new_net_2050)
	);

	bfr new_net_2052_bfr_before (
		.din(new_net_2052),
		.dout(new_net_2051)
	);

	bfr new_net_2053_bfr_before (
		.din(new_net_2053),
		.dout(new_net_2052)
	);

	bfr new_net_2054_bfr_before (
		.din(new_net_2054),
		.dout(new_net_2053)
	);

	bfr new_net_2055_bfr_before (
		.din(new_net_2055),
		.dout(new_net_2054)
	);

	spl3L new_net_1150_v_fanout (
		.a(new_net_1150),
		.b(new_net_525),
		.c(new_net_2055),
		.d(new_net_526)
	);

	bfr new_net_2056_bfr_before (
		.din(new_net_2056),
		.dout(new_net_1074)
	);

	spl2 new_net_1073_v_fanout (
		.a(new_net_1073),
		.b(new_net_2056),
		.c(new_net_543)
	);

	spl3L _0377__v_fanout (
		.a(_0377_),
		.b(new_net_1187),
		.c(new_net_1188),
		.d(new_net_1186)
	);

	spl4L _0057__v_fanout (
		.a(_0057_),
		.b(new_net_940),
		.c(new_net_938),
		.d(new_net_937),
		.e(new_net_939)
	);

	bfr new_net_2057_bfr_before (
		.din(new_net_2057),
		.dout(new_net_1142)
	);

	spl2 new_net_1141_v_fanout (
		.a(new_net_1141),
		.b(new_net_384),
		.c(new_net_2057)
	);

	spl2 _0045__v_fanout (
		.a(_0045_),
		.b(new_net_1183),
		.c(new_net_1184)
	);

	spl2 _0367__v_fanout (
		.a(_0367_),
		.b(new_net_186),
		.c(new_net_185)
	);

	spl2 new_net_1162_v_fanout (
		.a(new_net_1162),
		.b(new_net_1163),
		.c(new_net_689)
	);

	bfr new_net_2058_bfr_before (
		.din(new_net_2058),
		.dout(new_net_114)
	);

	bfr new_net_2059_bfr_before (
		.din(new_net_2059),
		.dout(new_net_2058)
	);

	bfr new_net_2060_bfr_before (
		.din(new_net_2060),
		.dout(new_net_2059)
	);

	spl4L _0213__v_fanout (
		.a(_0213_),
		.b(new_net_116),
		.c(new_net_117),
		.d(new_net_2060),
		.e(new_net_115)
	);

	spl2 _0154__v_fanout (
		.a(_0154_),
		.b(new_net_341),
		.c(new_net_340)
	);

	spl2 _0207__v_fanout (
		.a(_0207_),
		.b(new_net_1182),
		.c(new_net_952)
	);

	spl2 _0793__v_fanout (
		.a(_0793_),
		.b(new_net_771),
		.c(new_net_770)
	);

	bfr new_net_2061_bfr_before (
		.din(new_net_2061),
		.dout(new_net_1057)
	);

	spl2 new_net_1056_v_fanout (
		.a(new_net_1056),
		.b(new_net_2061),
		.c(new_net_614)
	);

	bfr new_net_2062_bfr_before (
		.din(new_net_2062),
		.dout(new_net_61)
	);

	bfr new_net_2063_bfr_before (
		.din(new_net_2063),
		.dout(new_net_2062)
	);

	bfr new_net_2064_bfr_before (
		.din(new_net_2064),
		.dout(new_net_2063)
	);

	spl2 new_net_1115_v_fanout (
		.a(new_net_1115),
		.b(new_net_2064),
		.c(new_net_55)
	);

	bfr new_net_2065_bfr_before (
		.din(new_net_2065),
		.dout(new_net_1070)
	);

	spl2 new_net_1069_v_fanout (
		.a(new_net_1069),
		.b(new_net_2065),
		.c(new_net_279)
	);

	spl2 _0362__v_fanout (
		.a(_0362_),
		.b(new_net_1030),
		.c(new_net_1029)
	);

	spl2 _0076__v_fanout (
		.a(_0076_),
		.b(new_net_632),
		.c(new_net_631)
	);

	spl2 _0060__v_fanout (
		.a(_0060_),
		.b(new_net_1181),
		.c(new_net_1180)
	);

	spl4L new_net_1177_v_fanout (
		.a(new_net_1177),
		.b(new_net_414),
		.c(new_net_411),
		.d(new_net_410),
		.e(new_net_413)
	);

	spl2 new_net_1171_v_fanout (
		.a(new_net_1171),
		.b(new_net_254),
		.c(new_net_252)
	);

	bfr new_net_2066_bfr_after (
		.din(_0359_),
		.dout(new_net_2066)
	);

	bfr new_net_2067_bfr_after (
		.din(new_net_2066),
		.dout(new_net_2067)
	);

	bfr new_net_2068_bfr_after (
		.din(new_net_2067),
		.dout(new_net_2068)
	);

	bfr new_net_2069_bfr_after (
		.din(new_net_2068),
		.dout(new_net_2069)
	);

	bfr new_net_2070_bfr_after (
		.din(new_net_2069),
		.dout(new_net_2070)
	);

	bfr new_net_2071_bfr_after (
		.din(new_net_2070),
		.dout(new_net_2071)
	);

	bfr new_net_2072_bfr_after (
		.din(new_net_2071),
		.dout(new_net_2072)
	);

	bfr new_net_2073_bfr_after (
		.din(new_net_2072),
		.dout(new_net_2073)
	);

	bfr new_net_2074_bfr_after (
		.din(new_net_2073),
		.dout(new_net_2074)
	);

	bfr new_net_2075_bfr_after (
		.din(new_net_2074),
		.dout(new_net_2075)
	);

	bfr new_net_2076_bfr_before (
		.din(new_net_2076),
		.dout(new_net_79)
	);

	bfr new_net_2077_bfr_before (
		.din(new_net_2077),
		.dout(new_net_2076)
	);

	bfr new_net_2078_bfr_before (
		.din(new_net_2078),
		.dout(new_net_80)
	);

	spl4L _0359__v_fanout (
		.a(new_net_2075),
		.b(new_net_1179),
		.c(new_net_1178),
		.d(new_net_2077),
		.e(new_net_2078)
	);

	bfr new_net_2079_bfr_before (
		.din(new_net_2079),
		.dout(new_net_716)
	);

	bfr new_net_2080_bfr_before (
		.din(new_net_2080),
		.dout(new_net_1168)
	);

	bfr new_net_2081_bfr_before (
		.din(new_net_2081),
		.dout(new_net_2080)
	);

	bfr new_net_2082_bfr_before (
		.din(new_net_2082),
		.dout(new_net_2081)
	);

	spl3L new_net_1167_v_fanout (
		.a(new_net_1167),
		.b(new_net_718),
		.c(new_net_2082),
		.d(new_net_2079)
	);

	bfr new_net_2083_bfr_before (
		.din(new_net_2083),
		.dout(new_net_250)
	);

	bfr new_net_2084_bfr_before (
		.din(new_net_2084),
		.dout(new_net_2083)
	);

	bfr new_net_2085_bfr_before (
		.din(new_net_2085),
		.dout(new_net_2084)
	);

	spl3L new_net_1172_v_fanout (
		.a(new_net_1172),
		.b(new_net_253),
		.c(new_net_251),
		.d(new_net_2085)
	);

	spl2 _0027__v_fanout (
		.a(_0027_),
		.b(new_net_1185),
		.c(new_net_276)
	);

	bfr new_net_2086_bfr_before (
		.din(new_net_2086),
		.dout(new_net_184)
	);

	bfr new_net_2087_bfr_before (
		.din(new_net_2087),
		.dout(new_net_2086)
	);

	bfr new_net_2088_bfr_before (
		.din(new_net_2088),
		.dout(new_net_2087)
	);

	spl2 _0796__v_fanout (
		.a(_0796_),
		.b(new_net_2088),
		.c(new_net_183)
	);

	bfr new_net_2089_bfr_before (
		.din(new_net_2089),
		.dout(new_net_1092)
	);

	bfr new_net_2090_bfr_before (
		.din(new_net_2090),
		.dout(new_net_2089)
	);

	bfr new_net_2091_bfr_before (
		.din(new_net_2091),
		.dout(new_net_2090)
	);

	bfr new_net_2092_bfr_before (
		.din(new_net_2092),
		.dout(new_net_2091)
	);

	spl2 new_net_1091_v_fanout (
		.a(new_net_1091),
		.b(new_net_2092),
		.c(new_net_157)
	);

	spl2 new_net_1144_v_fanout (
		.a(new_net_1144),
		.b(new_net_87),
		.c(new_net_85)
	);

	bfr new_net_2093_bfr_before (
		.din(new_net_2093),
		.dout(new_net_113)
	);

	bfr new_net_2094_bfr_before (
		.din(new_net_2094),
		.dout(new_net_2093)
	);

	bfr new_net_2095_bfr_before (
		.din(new_net_2095),
		.dout(new_net_2094)
	);

	bfr new_net_2096_bfr_before (
		.din(new_net_2096),
		.dout(new_net_2095)
	);

	bfr new_net_2097_bfr_before (
		.din(new_net_2097),
		.dout(new_net_2096)
	);

	bfr new_net_2098_bfr_before (
		.din(new_net_2098),
		.dout(new_net_2097)
	);

	bfr new_net_2099_bfr_before (
		.din(new_net_2099),
		.dout(new_net_2098)
	);

	bfr new_net_2100_bfr_before (
		.din(new_net_2100),
		.dout(new_net_2099)
	);

	bfr new_net_2101_bfr_before (
		.din(new_net_2101),
		.dout(new_net_2100)
	);

	bfr new_net_2102_bfr_before (
		.din(new_net_2102),
		.dout(new_net_2101)
	);

	bfr new_net_2103_bfr_before (
		.din(new_net_2103),
		.dout(new_net_2102)
	);

	bfr new_net_2104_bfr_before (
		.din(new_net_2104),
		.dout(new_net_2103)
	);

	bfr new_net_2105_bfr_before (
		.din(new_net_2105),
		.dout(new_net_2104)
	);

	bfr new_net_2106_bfr_before (
		.din(new_net_2106),
		.dout(new_net_2105)
	);

	bfr new_net_2107_bfr_before (
		.din(new_net_2107),
		.dout(new_net_2106)
	);

	bfr new_net_2108_bfr_before (
		.din(new_net_2108),
		.dout(new_net_2107)
	);

	bfr new_net_2109_bfr_before (
		.din(new_net_2109),
		.dout(new_net_2108)
	);

	bfr new_net_2110_bfr_before (
		.din(new_net_2110),
		.dout(new_net_2109)
	);

	bfr new_net_2111_bfr_before (
		.din(new_net_2111),
		.dout(new_net_2110)
	);

	bfr new_net_2112_bfr_before (
		.din(new_net_2112),
		.dout(new_net_2111)
	);

	bfr new_net_2113_bfr_before (
		.din(new_net_2113),
		.dout(new_net_2112)
	);

	bfr new_net_2114_bfr_before (
		.din(new_net_2114),
		.dout(new_net_2113)
	);

	bfr new_net_2115_bfr_before (
		.din(new_net_2115),
		.dout(new_net_2114)
	);

	bfr new_net_2116_bfr_before (
		.din(new_net_2116),
		.dout(new_net_2115)
	);

	bfr new_net_2117_bfr_before (
		.din(new_net_2117),
		.dout(new_net_2116)
	);

	bfr new_net_2118_bfr_before (
		.din(new_net_2118),
		.dout(new_net_2117)
	);

	bfr new_net_2119_bfr_before (
		.din(new_net_2119),
		.dout(new_net_2118)
	);

	bfr new_net_2120_bfr_before (
		.din(new_net_2120),
		.dout(new_net_2119)
	);

	bfr new_net_2121_bfr_before (
		.din(new_net_2121),
		.dout(new_net_2120)
	);

	bfr new_net_2122_bfr_before (
		.din(new_net_2122),
		.dout(new_net_2121)
	);

	bfr new_net_2123_bfr_before (
		.din(new_net_2123),
		.dout(new_net_2122)
	);

	bfr new_net_2124_bfr_before (
		.din(new_net_2124),
		.dout(new_net_2123)
	);

	bfr new_net_2125_bfr_before (
		.din(new_net_2125),
		.dout(new_net_2124)
	);

	bfr new_net_2126_bfr_before (
		.din(new_net_2126),
		.dout(new_net_2125)
	);

	bfr new_net_2127_bfr_before (
		.din(new_net_2127),
		.dout(new_net_2126)
	);

	bfr new_net_2128_bfr_before (
		.din(new_net_2128),
		.dout(new_net_2127)
	);

	bfr new_net_2129_bfr_before (
		.din(new_net_2129),
		.dout(new_net_2128)
	);

	bfr new_net_2130_bfr_before (
		.din(new_net_2130),
		.dout(new_net_2129)
	);

	bfr new_net_2131_bfr_before (
		.din(new_net_2131),
		.dout(new_net_2130)
	);

	bfr new_net_2132_bfr_before (
		.din(new_net_2132),
		.dout(new_net_2131)
	);

	bfr new_net_2133_bfr_before (
		.din(new_net_2133),
		.dout(new_net_2132)
	);

	bfr new_net_2134_bfr_before (
		.din(new_net_2134),
		.dout(new_net_2133)
	);

	spl2 new_net_1086_v_fanout (
		.a(new_net_1086),
		.b(new_net_112),
		.c(new_net_2134)
	);

	spl2 _0103__v_fanout (
		.a(_0103_),
		.b(new_net_884),
		.c(new_net_883)
	);

	bfr new_net_2135_bfr_before (
		.din(new_net_2135),
		.dout(new_net_1173)
	);

	bfr new_net_2136_bfr_before (
		.din(new_net_2136),
		.dout(new_net_2135)
	);

	spl2 _0382__v_fanout (
		.a(_0382_),
		.b(new_net_2136),
		.c(new_net_198)
	);

	bfr new_net_2137_bfr_before (
		.din(new_net_2137),
		.dout(new_net_68)
	);

	spl3L _0028__v_fanout (
		.a(_0028_),
		.b(new_net_2137),
		.c(new_net_69),
		.d(new_net_67)
	);

	spl2 _0039__v_fanout (
		.a(_0039_),
		.b(new_net_700),
		.c(new_net_699)
	);

	bfr new_net_2138_bfr_after (
		.din(_0356_),
		.dout(new_net_2138)
	);

	bfr new_net_2139_bfr_after (
		.din(new_net_2138),
		.dout(new_net_2139)
	);

	bfr new_net_2140_bfr_after (
		.din(new_net_2139),
		.dout(new_net_2140)
	);

	bfr new_net_2141_bfr_after (
		.din(new_net_2140),
		.dout(new_net_2141)
	);

	bfr new_net_2142_bfr_after (
		.din(new_net_2141),
		.dout(new_net_2142)
	);

	bfr new_net_2143_bfr_after (
		.din(new_net_2142),
		.dout(new_net_2143)
	);

	bfr new_net_2144_bfr_after (
		.din(new_net_2143),
		.dout(new_net_2144)
	);

	bfr new_net_2145_bfr_after (
		.din(new_net_2144),
		.dout(new_net_2145)
	);

	bfr new_net_2146_bfr_after (
		.din(new_net_2145),
		.dout(new_net_2146)
	);

	bfr new_net_2147_bfr_after (
		.din(new_net_2146),
		.dout(new_net_2147)
	);

	bfr new_net_2148_bfr_after (
		.din(new_net_2147),
		.dout(new_net_2148)
	);

	bfr new_net_2149_bfr_after (
		.din(new_net_2148),
		.dout(new_net_2149)
	);

	bfr new_net_2150_bfr_after (
		.din(new_net_2149),
		.dout(new_net_2150)
	);

	bfr new_net_2151_bfr_after (
		.din(new_net_2150),
		.dout(new_net_2151)
	);

	bfr new_net_2152_bfr_after (
		.din(new_net_2151),
		.dout(new_net_2152)
	);

	bfr new_net_2153_bfr_after (
		.din(new_net_2152),
		.dout(new_net_2153)
	);

	spl4L _0356__v_fanout (
		.a(new_net_2153),
		.b(new_net_238),
		.c(new_net_239),
		.d(new_net_236),
		.e(new_net_237)
	);

	spl2 _0068__v_fanout (
		.a(_0068_),
		.b(new_net_1172),
		.c(new_net_1171)
	);

	spl2 _0074__v_fanout (
		.a(_0074_),
		.b(new_net_1176),
		.c(new_net_1177)
	);

	spl2 _0020__v_fanout (
		.a(_0020_),
		.b(new_net_104),
		.c(new_net_103)
	);

	spl2 new_net_1158_v_fanout (
		.a(new_net_1158),
		.b(new_net_270),
		.c(new_net_269)
	);

	spl2 _0017__v_fanout (
		.a(_0017_),
		.b(new_net_390),
		.c(new_net_389)
	);

	bfr new_net_2154_bfr_before (
		.din(new_net_2154),
		.dout(new_net_46)
	);

	bfr new_net_2155_bfr_before (
		.din(new_net_2155),
		.dout(new_net_2154)
	);

	spl3L _0652__v_fanout (
		.a(_0652_),
		.b(new_net_47),
		.c(new_net_48),
		.d(new_net_2155)
	);

	bfr new_net_2156_bfr_before (
		.din(new_net_2156),
		.dout(new_net_578)
	);

	bfr new_net_2157_bfr_before (
		.din(new_net_2157),
		.dout(new_net_2156)
	);

	spl2 _0047__v_fanout (
		.a(_0047_),
		.b(new_net_579),
		.c(new_net_2157)
	);

	spl3L _0631__v_fanout (
		.a(_0631_),
		.b(new_net_773),
		.c(new_net_774),
		.d(new_net_772)
	);

	bfr new_net_2158_bfr_after (
		.din(_0365_),
		.dout(new_net_2158)
	);

	bfr new_net_2159_bfr_after (
		.din(new_net_2158),
		.dout(new_net_2159)
	);

	bfr new_net_2160_bfr_after (
		.din(new_net_2159),
		.dout(new_net_2160)
	);

	bfr new_net_2161_bfr_after (
		.din(new_net_2160),
		.dout(new_net_2161)
	);

	bfr new_net_2162_bfr_before (
		.din(new_net_2162),
		.dout(new_net_721)
	);

	spl2 _0365__v_fanout (
		.a(new_net_2161),
		.b(new_net_722),
		.c(new_net_2162)
	);

	bfr new_net_2163_bfr_before (
		.din(new_net_2163),
		.dout(new_net_493)
	);

	bfr new_net_2164_bfr_before (
		.din(new_net_2164),
		.dout(new_net_2163)
	);

	spl2 new_net_1138_v_fanout (
		.a(new_net_1138),
		.b(new_net_495),
		.c(new_net_2164)
	);

	bfr new_net_2165_bfr_before (
		.din(new_net_2165),
		.dout(new_net_235)
	);

	bfr new_net_2166_bfr_before (
		.din(new_net_2166),
		.dout(new_net_2165)
	);

	bfr new_net_2167_bfr_before (
		.din(new_net_2167),
		.dout(new_net_2166)
	);

	spl2 _0069__v_fanout (
		.a(_0069_),
		.b(new_net_2167),
		.c(new_net_234)
	);

	bfr new_net_2168_bfr_after (
		.din(_0517_),
		.dout(new_net_2168)
	);

	bfr new_net_2169_bfr_after (
		.din(new_net_2168),
		.dout(new_net_2169)
	);

	bfr new_net_2170_bfr_after (
		.din(new_net_2169),
		.dout(new_net_2170)
	);

	bfr new_net_2171_bfr_after (
		.din(new_net_2170),
		.dout(new_net_2171)
	);

	bfr new_net_2172_bfr_before (
		.din(new_net_2172),
		.dout(new_net_746)
	);

	spl2 _0517__v_fanout (
		.a(new_net_2171),
		.b(new_net_747),
		.c(new_net_2172)
	);

	spl2 new_net_1124_v_fanout (
		.a(new_net_1124),
		.b(new_net_791),
		.c(new_net_792)
	);

	spl2 _0008__v_fanout (
		.a(_0008_),
		.b(new_net_361),
		.c(new_net_360)
	);

	bfr new_net_2173_bfr_before (
		.din(new_net_2173),
		.dout(new_net_1115)
	);

	spl2 new_net_1114_v_fanout (
		.a(new_net_1114),
		.b(new_net_2173),
		.c(new_net_54)
	);

	spl2 _0011__v_fanout (
		.a(_0011_),
		.b(new_net_490),
		.c(new_net_489)
	);

	spl2 new_net_1161_v_fanout (
		.a(new_net_1161),
		.b(new_net_1162),
		.c(new_net_686)
	);

	spl2 _0036__v_fanout (
		.a(_0036_),
		.b(new_net_1002),
		.c(new_net_1001)
	);

	bfr new_net_2174_bfr_after (
		.din(_0151_),
		.dout(new_net_2174)
	);

	bfr new_net_2175_bfr_after (
		.din(new_net_2174),
		.dout(new_net_2175)
	);

	spl2 _0151__v_fanout (
		.a(new_net_2175),
		.b(new_net_259),
		.c(new_net_258)
	);

	bfr new_net_2176_bfr_before (
		.din(new_net_2176),
		.dout(new_net_949)
	);

	spl4L _0795__v_fanout (
		.a(_0795_),
		.b(new_net_2176),
		.c(new_net_947),
		.d(new_net_946),
		.e(new_net_948)
	);

	bfr new_net_2177_bfr_after (
		.din(_0360_),
		.dout(new_net_2177)
	);

	bfr new_net_2178_bfr_after (
		.din(new_net_2177),
		.dout(new_net_2178)
	);

	spl4L _0360__v_fanout (
		.a(new_net_2178),
		.b(new_net_133),
		.c(new_net_131),
		.d(new_net_130),
		.e(new_net_132)
	);

	bfr new_net_2179_bfr_before (
		.din(new_net_2179),
		.dout(new_net_667)
	);

	bfr new_net_2180_bfr_before (
		.din(new_net_2180),
		.dout(new_net_2179)
	);

	bfr new_net_2181_bfr_before (
		.din(new_net_2181),
		.dout(new_net_2180)
	);

	bfr new_net_2182_bfr_before (
		.din(new_net_2182),
		.dout(new_net_2181)
	);

	bfr new_net_2183_bfr_before (
		.din(new_net_2183),
		.dout(new_net_2182)
	);

	bfr new_net_2184_bfr_before (
		.din(new_net_2184),
		.dout(new_net_2183)
	);

	bfr new_net_2185_bfr_before (
		.din(new_net_2185),
		.dout(new_net_2184)
	);

	bfr new_net_2186_bfr_before (
		.din(new_net_2186),
		.dout(new_net_2185)
	);

	bfr new_net_2187_bfr_before (
		.din(new_net_2187),
		.dout(new_net_2186)
	);

	bfr new_net_2188_bfr_before (
		.din(new_net_2188),
		.dout(new_net_2187)
	);

	bfr new_net_2189_bfr_before (
		.din(new_net_2189),
		.dout(new_net_2188)
	);

	bfr new_net_2190_bfr_before (
		.din(new_net_2190),
		.dout(new_net_2189)
	);

	bfr new_net_2191_bfr_before (
		.din(new_net_2191),
		.dout(new_net_2190)
	);

	bfr new_net_2192_bfr_before (
		.din(new_net_2192),
		.dout(new_net_2191)
	);

	bfr new_net_2193_bfr_before (
		.din(new_net_2193),
		.dout(new_net_2192)
	);

	bfr new_net_2194_bfr_before (
		.din(new_net_2194),
		.dout(new_net_2193)
	);

	bfr new_net_2195_bfr_before (
		.din(new_net_2195),
		.dout(new_net_2194)
	);

	bfr new_net_2196_bfr_before (
		.din(new_net_2196),
		.dout(new_net_2195)
	);

	bfr new_net_2197_bfr_before (
		.din(new_net_2197),
		.dout(new_net_2196)
	);

	bfr new_net_2198_bfr_before (
		.din(new_net_2198),
		.dout(new_net_2197)
	);

	bfr new_net_2199_bfr_before (
		.din(new_net_2199),
		.dout(new_net_2198)
	);

	bfr new_net_2200_bfr_before (
		.din(new_net_2200),
		.dout(new_net_2199)
	);

	bfr new_net_2201_bfr_before (
		.din(new_net_2201),
		.dout(new_net_2200)
	);

	bfr new_net_2202_bfr_before (
		.din(new_net_2202),
		.dout(new_net_2201)
	);

	spl2 new_net_1133_v_fanout (
		.a(new_net_1133),
		.b(new_net_2202),
		.c(new_net_660)
	);

	bfr new_net_2203_bfr_before (
		.din(new_net_2203),
		.dout(new_net_233)
	);

	bfr new_net_2204_bfr_before (
		.din(new_net_2204),
		.dout(new_net_2203)
	);

	spl4L _0792__v_fanout (
		.a(_0792_),
		.b(new_net_2204),
		.c(new_net_231),
		.d(new_net_230),
		.e(new_net_232)
	);

	spl2 _0048__v_fanout (
		.a(_0048_),
		.b(new_net_271),
		.c(new_net_1158)
	);

	spl2 _0001__v_fanout (
		.a(_0001_),
		.b(new_net_26),
		.c(new_net_25)
	);

	bfr new_net_2205_bfr_before (
		.din(new_net_2205),
		.dout(new_net_74)
	);

	spl2 _0191__v_fanout (
		.a(_0191_),
		.b(new_net_2205),
		.c(new_net_73)
	);

	spl4L new_net_1093_v_fanout (
		.a(new_net_1093),
		.b(new_net_151),
		.c(new_net_175),
		.d(new_net_155),
		.e(new_net_1091)
	);

	spl4L new_net_1094_v_fanout (
		.a(new_net_1094),
		.b(new_net_158),
		.c(new_net_173),
		.d(new_net_177),
		.e(new_net_168)
	);

	spl3L new_net_1090_v_fanout (
		.a(new_net_1090),
		.b(new_net_169),
		.c(new_net_153),
		.d(new_net_176)
	);

	bfr new_net_2206_bfr_after (
		.din(_0093_),
		.dout(new_net_2206)
	);

	bfr new_net_2207_bfr_after (
		.din(new_net_2206),
		.dout(new_net_2207)
	);

	bfr new_net_2208_bfr_before (
		.din(new_net_2208),
		.dout(new_net_1164)
	);

	bfr new_net_2209_bfr_before (
		.din(new_net_2209),
		.dout(new_net_902)
	);

	bfr new_net_2210_bfr_before (
		.din(new_net_2210),
		.dout(new_net_908)
	);

	spl4L _0093__v_fanout (
		.a(new_net_2207),
		.b(new_net_2210),
		.c(new_net_903),
		.d(new_net_2208),
		.e(new_net_2209)
	);

	bfr new_net_2211_bfr_before (
		.din(new_net_2211),
		.dout(new_net_33)
	);

	bfr new_net_2212_bfr_before (
		.din(new_net_2212),
		.dout(new_net_2211)
	);

	bfr new_net_2213_bfr_before (
		.din(new_net_2213),
		.dout(new_net_2212)
	);

	spl4L new_net_1104_v_fanout (
		.a(new_net_1104),
		.b(new_net_40),
		.c(new_net_32),
		.d(new_net_2213),
		.e(new_net_37)
	);

	spl2 _0361__v_fanout (
		.a(_0361_),
		.b(new_net_776),
		.c(new_net_775)
	);

	bfr new_net_2214_bfr_before (
		.din(new_net_2214),
		.dout(new_net_1069)
	);

	bfr new_net_2215_bfr_before (
		.din(new_net_2215),
		.dout(new_net_2214)
	);

	spl2 new_net_1068_v_fanout (
		.a(new_net_1068),
		.b(new_net_2215),
		.c(new_net_287)
	);

	bfr new_net_2216_bfr_after (
		.din(_0672_),
		.dout(new_net_2216)
	);

	bfr new_net_2217_bfr_after (
		.din(new_net_2216),
		.dout(new_net_2217)
	);

	bfr new_net_2218_bfr_after (
		.din(new_net_2217),
		.dout(new_net_2218)
	);

	bfr new_net_2219_bfr_after (
		.din(new_net_2218),
		.dout(new_net_2219)
	);

	bfr new_net_2220_bfr_after (
		.din(new_net_2219),
		.dout(new_net_2220)
	);

	bfr new_net_2221_bfr_after (
		.din(new_net_2220),
		.dout(new_net_2221)
	);

	spl2 _0672__v_fanout (
		.a(new_net_2221),
		.b(new_net_784),
		.c(new_net_783)
	);

	bfr new_net_2222_bfr_before (
		.din(new_net_2222),
		.dout(new_net_1167)
	);

	spl2 _0794__v_fanout (
		.a(_0794_),
		.b(new_net_2222),
		.c(new_net_717)
	);

	spl2 _0189__v_fanout (
		.a(_0189_),
		.b(new_net_227),
		.c(new_net_226)
	);

	bfr new_net_2223_bfr_after (
		.din(_0116_),
		.dout(new_net_2223)
	);

	bfr new_net_2224_bfr_after (
		.din(new_net_2223),
		.dout(new_net_2224)
	);

	bfr new_net_2225_bfr_after (
		.din(new_net_2224),
		.dout(new_net_2225)
	);

	bfr new_net_2226_bfr_before (
		.din(new_net_2226),
		.dout(new_net_1169)
	);

	spl2 _0116__v_fanout (
		.a(new_net_2225),
		.b(new_net_503),
		.c(new_net_2226)
	);

	bfr new_net_2227_bfr_after (
		.din(_0770_),
		.dout(new_net_2227)
	);

	bfr new_net_2228_bfr_before (
		.din(new_net_2228),
		.dout(new_net_715)
	);

	bfr new_net_2229_bfr_before (
		.din(new_net_2229),
		.dout(new_net_2228)
	);

	bfr new_net_2230_bfr_before (
		.din(new_net_2230),
		.dout(new_net_2229)
	);

	spl2 _0770__v_fanout (
		.a(new_net_2227),
		.b(new_net_2230),
		.c(new_net_714)
	);

	bfr new_net_2231_bfr_after (
		.din(_0095_),
		.dout(new_net_2231)
	);

	bfr new_net_2232_bfr_before (
		.din(new_net_2232),
		.dout(new_net_1044)
	);

	bfr new_net_2233_bfr_before (
		.din(new_net_2233),
		.dout(new_net_2232)
	);

	bfr new_net_2234_bfr_before (
		.din(new_net_2234),
		.dout(new_net_2233)
	);

	bfr new_net_2235_bfr_before (
		.din(new_net_2235),
		.dout(new_net_2234)
	);

	bfr new_net_2236_bfr_before (
		.din(new_net_2236),
		.dout(new_net_2235)
	);

	bfr new_net_2237_bfr_before (
		.din(new_net_2237),
		.dout(new_net_2236)
	);

	spl2 _0095__v_fanout (
		.a(new_net_2231),
		.b(new_net_2237),
		.c(new_net_1043)
	);

	bfr new_net_2238_bfr_after (
		.din(_0644_),
		.dout(new_net_2238)
	);

	bfr new_net_2239_bfr_after (
		.din(new_net_2238),
		.dout(new_net_2239)
	);

	bfr new_net_2240_bfr_after (
		.din(new_net_2239),
		.dout(new_net_2240)
	);

	bfr new_net_2241_bfr_after (
		.din(new_net_2240),
		.dout(new_net_2241)
	);

	bfr new_net_2242_bfr_after (
		.din(new_net_2241),
		.dout(new_net_2242)
	);

	bfr new_net_2243_bfr_before (
		.din(new_net_2243),
		.dout(new_net_840)
	);

	spl2 _0644__v_fanout (
		.a(new_net_2242),
		.b(new_net_841),
		.c(new_net_2243)
	);

	bfr new_net_2244_bfr_after (
		.din(_0398_),
		.dout(new_net_2244)
	);

	bfr new_net_2245_bfr_after (
		.din(new_net_2244),
		.dout(new_net_2245)
	);

	bfr new_net_2246_bfr_after (
		.din(new_net_2245),
		.dout(new_net_2246)
	);

	bfr new_net_2247_bfr_after (
		.din(new_net_2246),
		.dout(new_net_2247)
	);

	bfr new_net_2248_bfr_after (
		.din(new_net_2247),
		.dout(new_net_2248)
	);

	bfr new_net_2249_bfr_before (
		.din(new_net_2249),
		.dout(new_net_470)
	);

	spl2 _0398__v_fanout (
		.a(new_net_2248),
		.b(new_net_2249),
		.c(new_net_469)
	);

	bfr new_net_2250_bfr_after (
		.din(_0383_),
		.dout(new_net_2250)
	);

	bfr new_net_2251_bfr_after (
		.din(new_net_2250),
		.dout(new_net_2251)
	);

	bfr new_net_2252_bfr_after (
		.din(new_net_2251),
		.dout(new_net_2252)
	);

	bfr new_net_2253_bfr_before (
		.din(new_net_2253),
		.dout(new_net_1166)
	);

	spl2 _0383__v_fanout (
		.a(new_net_2252),
		.b(new_net_2253),
		.c(new_net_972)
	);

	bfr new_net_2254_bfr_after (
		.din(_0172_),
		.dout(new_net_2254)
	);

	bfr new_net_2255_bfr_after (
		.din(new_net_2254),
		.dout(new_net_2255)
	);

	bfr new_net_2256_bfr_after (
		.din(new_net_2255),
		.dout(new_net_2256)
	);

	bfr new_net_2257_bfr_before (
		.din(new_net_2257),
		.dout(new_net_1159)
	);

	spl4L _0172__v_fanout (
		.a(new_net_2256),
		.b(new_net_2257),
		.c(new_net_191),
		.d(new_net_187),
		.e(new_net_188)
	);

	spl4L _0791__v_fanout (
		.a(_0791_),
		.b(new_net_1161),
		.c(new_net_691),
		.d(new_net_685),
		.e(new_net_688)
	);

	bfr new_net_2258_bfr_after (
		.din(_0439_),
		.dout(new_net_2258)
	);

	bfr new_net_2259_bfr_after (
		.din(new_net_2258),
		.dout(new_net_2259)
	);

	bfr new_net_2260_bfr_after (
		.din(new_net_2259),
		.dout(new_net_2260)
	);

	bfr new_net_2261_bfr_after (
		.din(new_net_2260),
		.dout(new_net_2261)
	);

	bfr new_net_2262_bfr_after (
		.din(new_net_2261),
		.dout(new_net_2262)
	);

	bfr new_net_2263_bfr_before (
		.din(new_net_2263),
		.dout(new_net_888)
	);

	spl2 _0439__v_fanout (
		.a(new_net_2262),
		.b(new_net_889),
		.c(new_net_2263)
	);

	bfr new_net_2264_bfr_before (
		.din(new_net_2264),
		.dout(new_net_1114)
	);

	spl2 new_net_1113_v_fanout (
		.a(new_net_1113),
		.b(new_net_58),
		.c(new_net_2264)
	);

	bfr new_net_2265_bfr_after (
		.din(_0416_),
		.dout(new_net_2265)
	);

	bfr new_net_2266_bfr_after (
		.din(new_net_2265),
		.dout(new_net_2266)
	);

	bfr new_net_2267_bfr_after (
		.din(new_net_2266),
		.dout(new_net_2267)
	);

	bfr new_net_2268_bfr_after (
		.din(new_net_2267),
		.dout(new_net_2268)
	);

	bfr new_net_2269_bfr_after (
		.din(new_net_2268),
		.dout(new_net_2269)
	);

	bfr new_net_2270_bfr_after (
		.din(new_net_2269),
		.dout(new_net_2270)
	);

	bfr new_net_2271_bfr_before (
		.din(new_net_2271),
		.dout(new_net_811)
	);

	spl2 _0416__v_fanout (
		.a(new_net_2270),
		.b(new_net_2271),
		.c(new_net_810)
	);

	bfr new_net_2272_bfr_before (
		.din(new_net_2272),
		.dout(new_net_352)
	);

	spl3L new_net_1108_v_fanout (
		.a(new_net_1108),
		.b(new_net_2272),
		.c(new_net_354),
		.d(new_net_350)
	);

	spl2 new_net_1063_v_fanout (
		.a(new_net_1063),
		.b(new_net_897),
		.c(new_net_894)
	);

	spl2 new_net_1078_v_fanout (
		.a(new_net_1078),
		.b(new_net_242),
		.c(new_net_245)
	);

	bfr new_net_2273_bfr_before (
		.din(new_net_2273),
		.dout(new_net_125)
	);

	bfr new_net_2274_bfr_before (
		.din(new_net_2274),
		.dout(new_net_2273)
	);

	bfr new_net_2275_bfr_before (
		.din(new_net_2275),
		.dout(new_net_2274)
	);

	bfr new_net_2276_bfr_before (
		.din(new_net_2276),
		.dout(new_net_2275)
	);

	bfr new_net_2277_bfr_before (
		.din(new_net_2277),
		.dout(new_net_2276)
	);

	bfr new_net_2278_bfr_before (
		.din(new_net_2278),
		.dout(new_net_2277)
	);

	bfr new_net_2279_bfr_before (
		.din(new_net_2279),
		.dout(new_net_2278)
	);

	bfr new_net_2280_bfr_before (
		.din(new_net_2280),
		.dout(new_net_2279)
	);

	bfr new_net_2281_bfr_before (
		.din(new_net_2281),
		.dout(new_net_2280)
	);

	bfr new_net_2282_bfr_before (
		.din(new_net_2282),
		.dout(new_net_2281)
	);

	bfr new_net_2283_bfr_before (
		.din(new_net_2283),
		.dout(new_net_2282)
	);

	spl2 new_net_1087_v_fanout (
		.a(new_net_1087),
		.b(new_net_126),
		.c(new_net_2283)
	);

	spl3L new_net_1067_v_fanout (
		.a(new_net_1067),
		.b(new_net_284),
		.c(new_net_278),
		.d(new_net_1068)
	);

	bfr new_net_2284_bfr_before (
		.din(new_net_2284),
		.dout(new_net_1141)
	);

	bfr new_net_2285_bfr_before (
		.din(new_net_2285),
		.dout(new_net_2284)
	);

	bfr new_net_2286_bfr_before (
		.din(new_net_2286),
		.dout(new_net_2285)
	);

	spl2 new_net_1140_v_fanout (
		.a(new_net_1140),
		.b(new_net_2286),
		.c(new_net_380)
	);

	bfr new_net_2287_bfr_after (
		.din(_0085_),
		.dout(new_net_2287)
	);

	bfr new_net_2288_bfr_after (
		.din(new_net_2287),
		.dout(new_net_2288)
	);

	bfr new_net_2289_bfr_after (
		.din(new_net_2288),
		.dout(new_net_2289)
	);

	bfr new_net_2290_bfr_after (
		.din(new_net_2289),
		.dout(new_net_2290)
	);

	bfr new_net_2291_bfr_after (
		.din(new_net_2290),
		.dout(new_net_2291)
	);

	bfr new_net_2292_bfr_after (
		.din(new_net_2291),
		.dout(new_net_2292)
	);

	bfr new_net_2293_bfr_after (
		.din(new_net_2292),
		.dout(new_net_2293)
	);

	bfr new_net_2294_bfr_after (
		.din(new_net_2293),
		.dout(new_net_2294)
	);

	bfr new_net_2295_bfr_before (
		.din(new_net_2295),
		.dout(new_net_1152)
	);

	bfr new_net_2296_bfr_before (
		.din(new_net_2296),
		.dout(new_net_1151)
	);

	spl3L _0085__v_fanout (
		.a(new_net_2294),
		.b(new_net_2296),
		.c(new_net_2295),
		.d(new_net_1035)
	);

	spl3L new_net_1134_v_fanout (
		.a(new_net_1134),
		.b(new_net_659),
		.c(new_net_664),
		.d(new_net_665)
	);

	spl4L new_net_1096_v_fanout (
		.a(new_net_1096),
		.b(new_net_170),
		.c(new_net_1090),
		.d(new_net_164),
		.e(new_net_160)
	);

	spl2 new_net_1050_v_fanout (
		.a(new_net_1050),
		.b(new_net_139),
		.c(new_net_137)
	);

	bfr new_net_2297_bfr_before (
		.din(new_net_2297),
		.dout(new_net_845)
	);

	bfr new_net_2298_bfr_before (
		.din(new_net_2298),
		.dout(new_net_2297)
	);

	bfr new_net_2299_bfr_before (
		.din(new_net_2299),
		.dout(new_net_2298)
	);

	bfr new_net_2300_bfr_before (
		.din(new_net_2300),
		.dout(new_net_2299)
	);

	spl3L new_net_1129_v_fanout (
		.a(new_net_1129),
		.b(new_net_847),
		.c(new_net_2300),
		.d(new_net_844)
	);

	bfr new_net_2301_bfr_before (
		.din(new_net_2301),
		.dout(new_net_159)
	);

	bfr new_net_2302_bfr_before (
		.din(new_net_2302),
		.dout(new_net_165)
	);

	spl4L new_net_1099_v_fanout (
		.a(new_net_1099),
		.b(new_net_2302),
		.c(new_net_166),
		.d(new_net_163),
		.e(new_net_2301)
	);

	bfr new_net_2303_bfr_before (
		.din(new_net_2303),
		.dout(new_net_1138)
	);

	spl2 new_net_1137_v_fanout (
		.a(new_net_1137),
		.b(new_net_2303),
		.c(new_net_492)
	);

	bfr new_net_2304_bfr_after (
		.din(_0489_),
		.dout(new_net_2304)
	);

	bfr new_net_2305_bfr_after (
		.din(new_net_2304),
		.dout(new_net_2305)
	);

	bfr new_net_2306_bfr_after (
		.din(new_net_2305),
		.dout(new_net_2306)
	);

	bfr new_net_2307_bfr_after (
		.din(new_net_2306),
		.dout(new_net_2307)
	);

	bfr new_net_2308_bfr_after (
		.din(new_net_2307),
		.dout(new_net_2308)
	);

	bfr new_net_2309_bfr_after (
		.din(new_net_2308),
		.dout(new_net_2309)
	);

	bfr new_net_2310_bfr_before (
		.din(new_net_2310),
		.dout(new_net_295)
	);

	spl2 _0489__v_fanout (
		.a(new_net_2309),
		.b(new_net_296),
		.c(new_net_2310)
	);

	spl4L new_net_1097_v_fanout (
		.a(new_net_1097),
		.b(new_net_162),
		.c(new_net_1094),
		.d(new_net_1093),
		.e(new_net_178)
	);

	bfr new_net_2311_bfr_before (
		.din(new_net_2311),
		.dout(new_net_1080)
	);

	bfr new_net_2312_bfr_before (
		.din(new_net_2312),
		.dout(new_net_2311)
	);

	bfr new_net_2313_bfr_before (
		.din(new_net_2313),
		.dout(new_net_2312)
	);

	bfr new_net_2314_bfr_before (
		.din(new_net_2314),
		.dout(new_net_2313)
	);

	bfr new_net_2315_bfr_before (
		.din(new_net_2315),
		.dout(new_net_2314)
	);

	bfr new_net_2316_bfr_before (
		.din(new_net_2316),
		.dout(new_net_2315)
	);

	spl3L new_net_1079_v_fanout (
		.a(new_net_1079),
		.b(new_net_597),
		.c(new_net_594),
		.d(new_net_2316)
	);

	spl2 new_net_1055_v_fanout (
		.a(new_net_1055),
		.b(new_net_1056),
		.c(new_net_613)
	);

	bfr new_net_2317_bfr_before (
		.din(new_net_2317),
		.dout(new_net_1144)
	);

	bfr new_net_2318_bfr_before (
		.din(new_net_2318),
		.dout(new_net_2317)
	);

	spl2 new_net_1143_v_fanout (
		.a(new_net_1143),
		.b(new_net_2318),
		.c(new_net_84)
	);

	bfr new_net_2319_bfr_before (
		.din(new_net_2319),
		.dout(new_net_149)
	);

	spl4L new_net_1095_v_fanout (
		.a(new_net_1095),
		.b(new_net_179),
		.c(new_net_174),
		.d(new_net_2319),
		.e(new_net_156)
	);

	spl2 new_net_1103_v_fanout (
		.a(new_net_1103),
		.b(new_net_1104),
		.c(new_net_43)
	);

	spl2 new_net_1132_v_fanout (
		.a(new_net_1132),
		.b(new_net_1133),
		.c(new_net_663)
	);

	bfr new_net_2320_bfr_after (
		.din(_0252_),
		.dout(new_net_2320)
	);

	bfr new_net_2321_bfr_after (
		.din(new_net_2320),
		.dout(new_net_2321)
	);

	bfr new_net_2322_bfr_after (
		.din(new_net_2321),
		.dout(new_net_2322)
	);

	bfr new_net_2323_bfr_before (
		.din(new_net_2323),
		.dout(new_net_912)
	);

	bfr new_net_2324_bfr_before (
		.din(new_net_2324),
		.dout(new_net_1153)
	);

	bfr new_net_2325_bfr_before (
		.din(new_net_2325),
		.dout(new_net_2324)
	);

	spl3L _0252__v_fanout (
		.a(new_net_2322),
		.b(new_net_2325),
		.c(new_net_2323),
		.d(new_net_910)
	);

	bfr new_net_2326_bfr_before (
		.din(new_net_2326),
		.dout(new_net_291)
	);

	bfr new_net_2327_bfr_before (
		.din(new_net_2327),
		.dout(new_net_2326)
	);

	bfr new_net_2328_bfr_before (
		.din(new_net_2328),
		.dout(new_net_2327)
	);

	spl2 new_net_1145_v_fanout (
		.a(new_net_1145),
		.b(new_net_294),
		.c(new_net_2328)
	);

	bfr new_net_2329_bfr_before (
		.din(new_net_2329),
		.dout(new_net_262)
	);

	bfr new_net_2330_bfr_before (
		.din(new_net_2330),
		.dout(new_net_2329)
	);

	bfr new_net_2331_bfr_before (
		.din(new_net_2331),
		.dout(new_net_2330)
	);

	bfr new_net_2332_bfr_before (
		.din(new_net_2332),
		.dout(new_net_2331)
	);

	bfr new_net_2333_bfr_before (
		.din(new_net_2333),
		.dout(new_net_2332)
	);

	bfr new_net_2334_bfr_before (
		.din(new_net_2334),
		.dout(new_net_2333)
	);

	bfr new_net_2335_bfr_before (
		.din(new_net_2335),
		.dout(new_net_2334)
	);

	bfr new_net_2336_bfr_before (
		.din(new_net_2336),
		.dout(new_net_2335)
	);

	spl3L new_net_1083_v_fanout (
		.a(new_net_1083),
		.b(new_net_2336),
		.c(new_net_263),
		.d(new_net_260)
	);

	bfr new_net_2337_bfr_after (
		.din(_0059_),
		.dout(new_net_2337)
	);

	bfr new_net_2338_bfr_after (
		.din(new_net_2337),
		.dout(new_net_2338)
	);

	bfr new_net_2339_bfr_after (
		.din(new_net_2338),
		.dout(new_net_2339)
	);

	bfr new_net_2340_bfr_after (
		.din(new_net_2339),
		.dout(new_net_2340)
	);

	spl4L _0059__v_fanout (
		.a(new_net_2340),
		.b(new_net_1148),
		.c(new_net_801),
		.d(new_net_796),
		.e(new_net_800)
	);

	bfr new_net_2341_bfr_before (
		.din(new_net_2341),
		.dout(new_net_1124)
	);

	bfr new_net_2342_bfr_before (
		.din(new_net_2342),
		.dout(new_net_2341)
	);

	spl2 new_net_1123_v_fanout (
		.a(new_net_1123),
		.b(new_net_795),
		.c(new_net_2342)
	);

	bfr new_net_2343_bfr_before (
		.din(new_net_2343),
		.dout(new_net_1119)
	);

	bfr new_net_2344_bfr_before (
		.din(new_net_2344),
		.dout(new_net_2343)
	);

	bfr new_net_2345_bfr_before (
		.din(new_net_2345),
		.dout(new_net_2344)
	);

	bfr new_net_2346_bfr_before (
		.din(new_net_2346),
		.dout(new_net_2345)
	);

	bfr new_net_2347_bfr_before (
		.din(new_net_2347),
		.dout(new_net_2346)
	);

	bfr new_net_2348_bfr_before (
		.din(new_net_2348),
		.dout(new_net_2347)
	);

	bfr new_net_2349_bfr_before (
		.din(new_net_2349),
		.dout(new_net_2348)
	);

	spl2 new_net_1118_v_fanout (
		.a(new_net_1118),
		.b(new_net_2349),
		.c(new_net_418)
	);

	bfr new_net_2350_bfr_after (
		.din(_0620_),
		.dout(new_net_2350)
	);

	bfr new_net_2351_bfr_after (
		.din(new_net_2350),
		.dout(new_net_2351)
	);

	bfr new_net_2352_bfr_before (
		.din(new_net_2352),
		.dout(new_net_1150)
	);

	spl2 _0620__v_fanout (
		.a(new_net_2351),
		.b(new_net_523),
		.c(new_net_2352)
	);

	spl2 new_net_1088_v_fanout (
		.a(new_net_1088),
		.b(new_net_861),
		.c(new_net_860)
	);

	bfr new_net_2353_bfr_after (
		.din(_0285_),
		.dout(new_net_2353)
	);

	bfr new_net_2354_bfr_after (
		.din(new_net_2353),
		.dout(new_net_2354)
	);

	bfr new_net_2355_bfr_after (
		.din(new_net_2354),
		.dout(new_net_2355)
	);

	bfr new_net_2356_bfr_after (
		.din(new_net_2355),
		.dout(new_net_2356)
	);

	bfr new_net_2357_bfr_before (
		.din(new_net_2357),
		.dout(new_net_10)
	);

	bfr new_net_2358_bfr_before (
		.din(new_net_2358),
		.dout(new_net_2357)
	);

	bfr new_net_2359_bfr_before (
		.din(new_net_2359),
		.dout(new_net_2358)
	);

	bfr new_net_2360_bfr_before (
		.din(new_net_2360),
		.dout(new_net_2359)
	);

	bfr new_net_2361_bfr_before (
		.din(new_net_2361),
		.dout(new_net_2360)
	);

	bfr new_net_2362_bfr_before (
		.din(new_net_2362),
		.dout(new_net_2361)
	);

	bfr new_net_2363_bfr_before (
		.din(new_net_2363),
		.dout(new_net_2362)
	);

	bfr new_net_2364_bfr_before (
		.din(new_net_2364),
		.dout(new_net_2363)
	);

	bfr new_net_2365_bfr_before (
		.din(new_net_2365),
		.dout(new_net_2364)
	);

	bfr new_net_2366_bfr_before (
		.din(new_net_2366),
		.dout(new_net_2365)
	);

	bfr new_net_2367_bfr_before (
		.din(new_net_2367),
		.dout(new_net_2366)
	);

	bfr new_net_2368_bfr_before (
		.din(new_net_2368),
		.dout(new_net_2367)
	);

	bfr new_net_2369_bfr_before (
		.din(new_net_2369),
		.dout(new_net_2368)
	);

	bfr new_net_2370_bfr_before (
		.din(new_net_2370),
		.dout(new_net_2369)
	);

	bfr new_net_2371_bfr_before (
		.din(new_net_2371),
		.dout(new_net_2370)
	);

	bfr new_net_2372_bfr_before (
		.din(new_net_2372),
		.dout(new_net_2371)
	);

	bfr new_net_2373_bfr_before (
		.din(new_net_2373),
		.dout(new_net_2372)
	);

	bfr new_net_2374_bfr_before (
		.din(new_net_2374),
		.dout(new_net_2373)
	);

	bfr new_net_2375_bfr_before (
		.din(new_net_2375),
		.dout(new_net_2374)
	);

	bfr new_net_2376_bfr_before (
		.din(new_net_2376),
		.dout(new_net_2375)
	);

	bfr new_net_2377_bfr_before (
		.din(new_net_2377),
		.dout(new_net_2376)
	);

	bfr new_net_2378_bfr_before (
		.din(new_net_2378),
		.dout(new_net_2377)
	);

	bfr new_net_2379_bfr_before (
		.din(new_net_2379),
		.dout(new_net_2378)
	);

	bfr new_net_2380_bfr_before (
		.din(new_net_2380),
		.dout(new_net_2379)
	);

	bfr new_net_2381_bfr_before (
		.din(new_net_2381),
		.dout(new_net_2380)
	);

	bfr new_net_2382_bfr_before (
		.din(new_net_2382),
		.dout(new_net_2381)
	);

	bfr new_net_2383_bfr_before (
		.din(new_net_2383),
		.dout(new_net_2382)
	);

	bfr new_net_2384_bfr_before (
		.din(new_net_2384),
		.dout(new_net_2383)
	);

	bfr new_net_2385_bfr_before (
		.din(new_net_2385),
		.dout(new_net_2384)
	);

	bfr new_net_2386_bfr_before (
		.din(new_net_2386),
		.dout(new_net_2385)
	);

	bfr new_net_2387_bfr_before (
		.din(new_net_2387),
		.dout(new_net_2386)
	);

	bfr new_net_2388_bfr_before (
		.din(new_net_2388),
		.dout(new_net_2387)
	);

	bfr new_net_2389_bfr_before (
		.din(new_net_2389),
		.dout(new_net_2388)
	);

	bfr new_net_2390_bfr_before (
		.din(new_net_2390),
		.dout(new_net_2389)
	);

	bfr new_net_2391_bfr_before (
		.din(new_net_2391),
		.dout(new_net_2390)
	);

	bfr new_net_2392_bfr_before (
		.din(new_net_2392),
		.dout(new_net_2391)
	);

	bfr new_net_2393_bfr_before (
		.din(new_net_2393),
		.dout(new_net_2392)
	);

	bfr new_net_2394_bfr_before (
		.din(new_net_2394),
		.dout(new_net_2393)
	);

	bfr new_net_2395_bfr_before (
		.din(new_net_2395),
		.dout(new_net_2394)
	);

	bfr new_net_2396_bfr_before (
		.din(new_net_2396),
		.dout(new_net_2395)
	);

	bfr new_net_2397_bfr_before (
		.din(new_net_2397),
		.dout(new_net_2396)
	);

	bfr new_net_2398_bfr_before (
		.din(new_net_2398),
		.dout(new_net_2397)
	);

	bfr new_net_2399_bfr_before (
		.din(new_net_2399),
		.dout(new_net_2398)
	);

	spl2 _0285__v_fanout (
		.a(new_net_2356),
		.b(new_net_2399),
		.c(new_net_9)
	);

	bfr new_net_2400_bfr_before (
		.din(new_net_2400),
		.dout(new_net_152)
	);

	spl4L new_net_1098_v_fanout (
		.a(new_net_1098),
		.b(new_net_150),
		.c(new_net_2400),
		.d(new_net_172),
		.e(new_net_161)
	);

	bfr new_net_2401_bfr_before (
		.din(new_net_2401),
		.dout(new_net_1155)
	);

	bfr new_net_2402_bfr_before (
		.din(new_net_2402),
		.dout(new_net_2401)
	);

	bfr new_net_2403_bfr_before (
		.din(new_net_2403),
		.dout(new_net_2402)
	);

	bfr new_net_2404_bfr_before (
		.din(new_net_2404),
		.dout(new_net_2403)
	);

	bfr new_net_2405_bfr_before (
		.din(new_net_2405),
		.dout(new_net_2404)
	);

	bfr new_net_2406_bfr_before (
		.din(new_net_2406),
		.dout(new_net_2405)
	);

	bfr new_net_2407_bfr_before (
		.din(new_net_2407),
		.dout(new_net_2406)
	);

	spl2 _0066__v_fanout (
		.a(_0066_),
		.b(new_net_2407),
		.c(new_net_143)
	);

	spl2 new_net_1112_v_fanout (
		.a(new_net_1112),
		.b(new_net_1113),
		.c(new_net_60)
	);

	spl2 new_net_1146_v_fanout (
		.a(new_net_1146),
		.b(new_net_290),
		.c(new_net_293)
	);

	spl2 new_net_1100_v_fanout (
		.a(new_net_1100),
		.b(new_net_1099),
		.c(new_net_1098)
	);

	spl3L new_net_1101_v_fanout (
		.a(new_net_1101),
		.b(new_net_1095),
		.c(new_net_1097),
		.d(new_net_1096)
	);

	bfr new_net_2408_bfr_before (
		.din(new_net_2408),
		.dout(new_net_409)
	);

	bfr new_net_2409_bfr_before (
		.din(new_net_2409),
		.dout(new_net_2408)
	);

	spl2 new_net_1053_v_fanout (
		.a(new_net_1053),
		.b(new_net_2409),
		.c(new_net_405)
	);

	bfr new_net_2410_bfr_before (
		.din(new_net_2410),
		.dout(new_net_39)
	);

	spl3L new_net_1107_v_fanout (
		.a(new_net_1107),
		.b(new_net_2410),
		.c(new_net_42),
		.d(new_net_34)
	);

	bfr new_net_2411_bfr_before (
		.din(new_net_2411),
		.dout(new_net_1073)
	);

	bfr new_net_2412_bfr_before (
		.din(new_net_2412),
		.dout(new_net_2411)
	);

	bfr new_net_2413_bfr_before (
		.din(new_net_2413),
		.dout(new_net_2412)
	);

	bfr new_net_2414_bfr_before (
		.din(new_net_2414),
		.dout(new_net_2413)
	);

	spl3L new_net_1076_v_fanout (
		.a(new_net_1076),
		.b(new_net_539),
		.c(new_net_537),
		.d(new_net_2414)
	);

	spl2 new_net_1075_v_fanout (
		.a(new_net_1075),
		.b(new_net_536),
		.c(new_net_542)
	);

	spl2 new_net_1109_v_fanout (
		.a(new_net_1109),
		.b(new_net_1108),
		.c(new_net_353)
	);

	bfr new_net_2415_bfr_before (
		.din(new_net_2415),
		.dout(new_net_217)
	);

	bfr new_net_2416_bfr_before (
		.din(new_net_2416),
		.dout(new_net_221)
	);

	bfr new_net_2417_bfr_before (
		.din(new_net_2417),
		.dout(new_net_2416)
	);

	spl3L new_net_1049_v_fanout (
		.a(new_net_1049),
		.b(new_net_219),
		.c(new_net_2417),
		.d(new_net_2415)
	);

	spl2 new_net_1051_v_fanout (
		.a(new_net_1051),
		.b(new_net_136),
		.c(new_net_138)
	);

	bfr new_net_2418_bfr_before (
		.din(new_net_2418),
		.dout(new_net_896)
	);

	bfr new_net_2419_bfr_before (
		.din(new_net_2419),
		.dout(new_net_1063)
	);

	bfr new_net_2420_bfr_before (
		.din(new_net_2420),
		.dout(new_net_2419)
	);

	bfr new_net_2421_bfr_before (
		.din(new_net_2421),
		.dout(new_net_2420)
	);

	bfr new_net_2422_bfr_before (
		.din(new_net_2422),
		.dout(new_net_2421)
	);

	spl4L new_net_1064_v_fanout (
		.a(new_net_1064),
		.b(new_net_2422),
		.c(new_net_898),
		.d(new_net_893),
		.e(new_net_2418)
	);

	spl2 new_net_1071_v_fanout (
		.a(new_net_1071),
		.b(new_net_280),
		.c(new_net_1067)
	);

	bfr new_net_2423_bfr_before (
		.din(new_net_2423),
		.dout(new_net_282)
	);

	spl4L new_net_1072_v_fanout (
		.a(new_net_1072),
		.b(new_net_285),
		.c(new_net_2423),
		.d(new_net_283),
		.e(new_net_281)
	);

	bfr new_net_2424_bfr_before (
		.din(new_net_2424),
		.dout(new_net_1121)
	);

	bfr new_net_2425_bfr_before (
		.din(new_net_2425),
		.dout(new_net_2424)
	);

	bfr new_net_2426_bfr_before (
		.din(new_net_2426),
		.dout(new_net_2425)
	);

	bfr new_net_2427_bfr_before (
		.din(new_net_2427),
		.dout(new_net_2426)
	);

	bfr new_net_2428_bfr_before (
		.din(new_net_2428),
		.dout(new_net_2427)
	);

	bfr new_net_2429_bfr_before (
		.din(new_net_2429),
		.dout(new_net_2428)
	);

	spl2 new_net_1120_v_fanout (
		.a(new_net_1120),
		.b(new_net_2429),
		.c(new_net_441)
	);

	bfr new_net_2430_bfr_before (
		.din(new_net_2430),
		.dout(new_net_15)
	);

	bfr new_net_2431_bfr_before (
		.din(new_net_2431),
		.dout(new_net_2430)
	);

	bfr new_net_2432_bfr_before (
		.din(new_net_2432),
		.dout(new_net_2431)
	);

	bfr new_net_2433_bfr_before (
		.din(new_net_2433),
		.dout(new_net_2432)
	);

	spl2 new_net_1062_v_fanout (
		.a(new_net_1062),
		.b(new_net_2433),
		.c(new_net_16)
	);

	bfr new_net_2434_bfr_before (
		.din(new_net_2434),
		.dout(new_net_36)
	);

	bfr new_net_2435_bfr_before (
		.din(new_net_2435),
		.dout(new_net_38)
	);

	spl4L new_net_1106_v_fanout (
		.a(new_net_1106),
		.b(new_net_2435),
		.c(new_net_35),
		.d(new_net_31),
		.e(new_net_2434)
	);

	spl2 new_net_1084_v_fanout (
		.a(new_net_1084),
		.b(new_net_261),
		.c(new_net_265)
	);

	bfr new_net_2436_bfr_before (
		.din(new_net_2436),
		.dout(new_net_891)
	);

	bfr new_net_2437_bfr_before (
		.din(new_net_2437),
		.dout(new_net_2436)
	);

	bfr new_net_2438_bfr_before (
		.din(new_net_2438),
		.dout(new_net_892)
	);

	spl4L new_net_1065_v_fanout (
		.a(new_net_1065),
		.b(new_net_2438),
		.c(new_net_895),
		.d(new_net_890),
		.e(new_net_2437)
	);

	bfr new_net_2439_bfr_before (
		.din(new_net_2439),
		.dout(new_net_633)
	);

	spl3L new_net_1060_v_fanout (
		.a(new_net_1060),
		.b(new_net_635),
		.c(new_net_637),
		.d(new_net_2439)
	);

	bfr new_net_2440_bfr_before (
		.din(new_net_2440),
		.dout(new_net_1078)
	);

	bfr new_net_2441_bfr_before (
		.din(new_net_2441),
		.dout(new_net_2440)
	);

	bfr new_net_2442_bfr_before (
		.din(new_net_2442),
		.dout(new_net_2441)
	);

	spl4L new_net_1077_v_fanout (
		.a(new_net_1077),
		.b(new_net_2442),
		.c(new_net_244),
		.d(new_net_240),
		.e(new_net_241)
	);

	bfr new_net_2443_bfr_before (
		.din(new_net_2443),
		.dout(new_net_1058)
	);

	bfr new_net_2444_bfr_before (
		.din(new_net_2444),
		.dout(new_net_2443)
	);

	bfr new_net_2445_bfr_before (
		.din(new_net_2445),
		.dout(new_net_2444)
	);

	bfr new_net_2446_bfr_before (
		.din(new_net_2446),
		.dout(new_net_2445)
	);

	bfr new_net_2447_bfr_before (
		.din(new_net_2447),
		.dout(new_net_2446)
	);

	bfr new_net_2448_bfr_before (
		.din(new_net_2448),
		.dout(new_net_2447)
	);

	spl2 new_net_1059_v_fanout (
		.a(new_net_1059),
		.b(new_net_2448),
		.c(new_net_638)
	);

	bfr new_net_2449_bfr_before (
		.din(new_net_2449),
		.dout(new_net_599)
	);

	bfr new_net_2450_bfr_before (
		.din(new_net_2450),
		.dout(new_net_2449)
	);

	bfr new_net_2451_bfr_before (
		.din(new_net_2451),
		.dout(new_net_595)
	);

	spl4L new_net_1082_v_fanout (
		.a(new_net_1082),
		.b(new_net_1079),
		.c(new_net_2451),
		.d(new_net_2450),
		.e(new_net_601)
	);

	spl4L new_net_1136_v_fanout (
		.a(new_net_1136),
		.b(new_net_666),
		.c(new_net_662),
		.d(new_net_668),
		.e(new_net_658)
	);

	spl3L new_net_1116_v_fanout (
		.a(new_net_1116),
		.b(new_net_53),
		.c(new_net_57),
		.d(new_net_56)
	);

	spl2 new_net_1105_v_fanout (
		.a(new_net_1105),
		.b(new_net_41),
		.c(new_net_1103)
	);

	spl2 new_net_1139_v_fanout (
		.a(new_net_1139),
		.b(new_net_1140),
		.c(new_net_381)
	);

	spl2 new_net_1117_v_fanout (
		.a(new_net_1117),
		.b(new_net_421),
		.c(new_net_1118)
	);

	spl3L new_net_1085_v_fanout (
		.a(new_net_1085),
		.b(new_net_266),
		.c(new_net_264),
		.d(new_net_1083)
	);

	spl4L new_net_1110_v_fanout (
		.a(new_net_1110),
		.b(new_net_351),
		.c(new_net_347),
		.d(new_net_348),
		.e(new_net_349)
	);

	spl4L new_net_1128_v_fanout (
		.a(new_net_1128),
		.b(new_net_1129),
		.c(new_net_846),
		.d(new_net_848),
		.e(new_net_843)
	);

	bfr new_net_2452_bfr_before (
		.din(new_net_2452),
		.dout(new_net_591)
	);

	bfr new_net_2453_bfr_before (
		.din(new_net_2453),
		.dout(new_net_2452)
	);

	bfr new_net_2454_bfr_before (
		.din(new_net_2454),
		.dout(new_net_598)
	);

	spl4L new_net_1081_v_fanout (
		.a(new_net_1081),
		.b(new_net_2454),
		.c(new_net_592),
		.d(new_net_2453),
		.e(new_net_596)
	);

	spl2 new_net_1048_v_fanout (
		.a(new_net_1048),
		.b(new_net_220),
		.c(new_net_218)
	);

	bfr new_net_2455_bfr_before (
		.din(new_net_2455),
		.dout(new_net_1050)
	);

	bfr new_net_2456_bfr_before (
		.din(new_net_2456),
		.dout(new_net_2455)
	);

	bfr new_net_2457_bfr_before (
		.din(new_net_2457),
		.dout(new_net_2456)
	);

	bfr new_net_2458_bfr_before (
		.din(new_net_2458),
		.dout(new_net_135)
	);

	bfr new_net_2459_bfr_before (
		.din(new_net_2459),
		.dout(new_net_2458)
	);

	spl3L new_net_1052_v_fanout (
		.a(new_net_1052),
		.b(new_net_134),
		.c(new_net_2459),
		.d(new_net_2457)
	);

	bfr new_net_2460_bfr_before (
		.din(new_net_2460),
		.dout(new_net_1126)
	);

	bfr new_net_2461_bfr_before (
		.din(new_net_2461),
		.dout(new_net_2460)
	);

	bfr new_net_2462_bfr_before (
		.din(new_net_2462),
		.dout(new_net_2461)
	);

	bfr new_net_2463_bfr_before (
		.din(new_net_2463),
		.dout(new_net_2462)
	);

	spl3L new_net_1125_v_fanout (
		.a(new_net_1125),
		.b(new_net_2463),
		.c(new_net_677),
		.d(new_net_673)
	);

	bfr new_net_2464_bfr_before (
		.din(new_net_2464),
		.dout(new_net_404)
	);

	bfr new_net_2465_bfr_before (
		.din(new_net_2465),
		.dout(new_net_2464)
	);

	bfr new_net_2466_bfr_before (
		.din(new_net_2466),
		.dout(new_net_2465)
	);

	bfr new_net_2467_bfr_before (
		.din(new_net_2467),
		.dout(new_net_2466)
	);

	bfr new_net_2468_bfr_before (
		.din(new_net_2468),
		.dout(new_net_406)
	);

	spl4L new_net_1054_v_fanout (
		.a(new_net_1054),
		.b(new_net_408),
		.c(new_net_407),
		.d(new_net_2467),
		.e(new_net_2468)
	);

	spl3L new_net_1147_v_fanout (
		.a(new_net_1147),
		.b(new_net_1145),
		.c(new_net_292),
		.d(new_net_289)
	);

	spl3L new_net_1122_v_fanout (
		.a(new_net_1122),
		.b(new_net_1123),
		.c(new_net_793),
		.d(new_net_789)
	);

	spl3L new_net_1135_v_fanout (
		.a(new_net_1135),
		.b(new_net_1132),
		.c(new_net_1134),
		.d(new_net_661)
	);

	bfr new_net_2469_bfr_before (
		.din(new_net_2469),
		.dout(new_net_436)
	);

	bfr new_net_2470_bfr_before (
		.din(new_net_2470),
		.dout(new_net_438)
	);

	bfr new_net_2471_bfr_before (
		.din(new_net_2471),
		.dout(new_net_437)
	);

	bfr new_net_2472_bfr_before (
		.din(new_net_2472),
		.dout(new_net_2471)
	);

	bfr new_net_2473_bfr_before (
		.din(new_net_2473),
		.dout(new_net_2472)
	);

	bfr new_net_2474_bfr_before (
		.din(new_net_2474),
		.dout(new_net_2473)
	);

	bfr new_net_2475_bfr_before (
		.din(new_net_2475),
		.dout(new_net_2474)
	);

	spl4L G37_v_fanout (
		.a(G37),
		.b(new_net_2475),
		.c(new_net_2470),
		.d(new_net_435),
		.e(new_net_2469)
	);

	bfr new_net_2476_bfr_after (
		.din(G16),
		.dout(new_net_2476)
	);

	bfr new_net_2477_bfr_after (
		.din(new_net_2476),
		.dout(new_net_2477)
	);

	bfr new_net_2478_bfr_after (
		.din(new_net_2477),
		.dout(new_net_2478)
	);

	bfr new_net_2479_bfr_after (
		.din(new_net_2478),
		.dout(new_net_2479)
	);

	bfr new_net_2480_bfr_after (
		.din(new_net_2479),
		.dout(new_net_2480)
	);

	bfr new_net_2481_bfr_after (
		.din(new_net_2480),
		.dout(new_net_2481)
	);

	bfr new_net_2482_bfr_after (
		.din(new_net_2481),
		.dout(new_net_2482)
	);

	bfr new_net_2483_bfr_after (
		.din(new_net_2482),
		.dout(new_net_2483)
	);

	bfr new_net_2484_bfr_after (
		.din(new_net_2483),
		.dout(new_net_2484)
	);

	spl2 G16_v_fanout (
		.a(new_net_2484),
		.b(new_net_319),
		.c(new_net_318)
	);

	bfr new_net_2485_bfr_after (
		.din(G38),
		.dout(new_net_2485)
	);

	bfr new_net_2486_bfr_after (
		.din(new_net_2485),
		.dout(new_net_2486)
	);

	bfr new_net_2487_bfr_after (
		.din(new_net_2486),
		.dout(new_net_2487)
	);

	bfr new_net_2488_bfr_before (
		.din(new_net_2488),
		.dout(new_net_692)
	);

	bfr new_net_2489_bfr_before (
		.din(new_net_2489),
		.dout(new_net_2488)
	);

	bfr new_net_2490_bfr_before (
		.din(new_net_2490),
		.dout(new_net_2489)
	);

	spl2 G38_v_fanout (
		.a(new_net_2487),
		.b(new_net_693),
		.c(new_net_2490)
	);

	spl2 G10_v_fanout (
		.a(G10),
		.b(new_net_1065),
		.c(new_net_1064)
	);

	bfr new_net_2491_bfr_after (
		.din(G50),
		.dout(new_net_2491)
	);

	bfr new_net_2492_bfr_after (
		.din(new_net_2491),
		.dout(new_net_2492)
	);

	bfr new_net_2493_bfr_after (
		.din(new_net_2492),
		.dout(new_net_2493)
	);

	bfr new_net_2494_bfr_after (
		.din(new_net_2493),
		.dout(new_net_2494)
	);

	bfr new_net_2495_bfr_after (
		.din(new_net_2494),
		.dout(new_net_2495)
	);

	bfr new_net_2496_bfr_after (
		.din(new_net_2495),
		.dout(new_net_2496)
	);

	bfr new_net_2497_bfr_after (
		.din(new_net_2496),
		.dout(new_net_2497)
	);

	bfr new_net_2498_bfr_after (
		.din(new_net_2497),
		.dout(new_net_2498)
	);

	bfr new_net_2499_bfr_after (
		.din(new_net_2498),
		.dout(new_net_2499)
	);

	bfr new_net_2500_bfr_after (
		.din(new_net_2499),
		.dout(new_net_2500)
	);

	bfr new_net_2501_bfr_after (
		.din(new_net_2500),
		.dout(new_net_2501)
	);

	bfr new_net_2502_bfr_after (
		.din(new_net_2501),
		.dout(new_net_2502)
	);

	bfr new_net_2503_bfr_after (
		.din(new_net_2502),
		.dout(new_net_2503)
	);

	bfr new_net_2504_bfr_after (
		.din(new_net_2503),
		.dout(new_net_2504)
	);

	bfr new_net_2505_bfr_after (
		.din(new_net_2504),
		.dout(new_net_2505)
	);

	bfr new_net_2506_bfr_after (
		.din(new_net_2505),
		.dout(new_net_2506)
	);

	bfr new_net_2507_bfr_after (
		.din(new_net_2506),
		.dout(new_net_2507)
	);

	bfr new_net_2508_bfr_after (
		.din(new_net_2507),
		.dout(new_net_2508)
	);

	bfr new_net_2509_bfr_after (
		.din(new_net_2508),
		.dout(new_net_2509)
	);

	bfr new_net_2510_bfr_after (
		.din(new_net_2509),
		.dout(new_net_2510)
	);

	bfr new_net_2511_bfr_after (
		.din(new_net_2510),
		.dout(new_net_2511)
	);

	bfr new_net_2512_bfr_after (
		.din(new_net_2511),
		.dout(new_net_2512)
	);

	bfr new_net_2513_bfr_after (
		.din(new_net_2512),
		.dout(new_net_2513)
	);

	bfr new_net_2514_bfr_after (
		.din(new_net_2513),
		.dout(new_net_2514)
	);

	bfr new_net_2515_bfr_after (
		.din(new_net_2514),
		.dout(new_net_2515)
	);

	bfr new_net_2516_bfr_after (
		.din(new_net_2515),
		.dout(new_net_2516)
	);

	bfr new_net_2517_bfr_after (
		.din(new_net_2516),
		.dout(new_net_2517)
	);

	bfr new_net_2518_bfr_after (
		.din(new_net_2517),
		.dout(new_net_2518)
	);

	bfr new_net_2519_bfr_after (
		.din(new_net_2518),
		.dout(new_net_2519)
	);

	bfr new_net_2520_bfr_after (
		.din(new_net_2519),
		.dout(new_net_2520)
	);

	bfr new_net_2521_bfr_after (
		.din(new_net_2520),
		.dout(new_net_2521)
	);

	bfr new_net_2522_bfr_after (
		.din(new_net_2521),
		.dout(new_net_2522)
	);

	bfr new_net_2523_bfr_after (
		.din(new_net_2522),
		.dout(new_net_2523)
	);

	bfr new_net_2524_bfr_after (
		.din(new_net_2523),
		.dout(new_net_2524)
	);

	bfr new_net_2525_bfr_after (
		.din(new_net_2524),
		.dout(new_net_2525)
	);

	bfr new_net_2526_bfr_after (
		.din(new_net_2525),
		.dout(new_net_2526)
	);

	bfr new_net_2527_bfr_after (
		.din(new_net_2526),
		.dout(new_net_2527)
	);

	bfr new_net_2528_bfr_after (
		.din(new_net_2527),
		.dout(new_net_2528)
	);

	bfr new_net_2529_bfr_after (
		.din(new_net_2528),
		.dout(new_net_2529)
	);

	bfr new_net_2530_bfr_after (
		.din(new_net_2529),
		.dout(new_net_2530)
	);

	bfr new_net_2531_bfr_after (
		.din(new_net_2530),
		.dout(new_net_2531)
	);

	bfr new_net_2532_bfr_after (
		.din(new_net_2531),
		.dout(new_net_2532)
	);

	bfr new_net_2533_bfr_after (
		.din(new_net_2532),
		.dout(new_net_2533)
	);

	bfr new_net_2534_bfr_after (
		.din(new_net_2533),
		.dout(new_net_2534)
	);

	bfr new_net_2535_bfr_after (
		.din(new_net_2534),
		.dout(new_net_2535)
	);

	bfr new_net_2536_bfr_after (
		.din(new_net_2535),
		.dout(new_net_2536)
	);

	bfr new_net_2537_bfr_after (
		.din(new_net_2536),
		.dout(new_net_2537)
	);

	bfr new_net_2538_bfr_after (
		.din(new_net_2537),
		.dout(new_net_2538)
	);

	spl2 G50_v_fanout (
		.a(new_net_2538),
		.b(new_net_209),
		.c(new_net_208)
	);

	spl2 G4_v_fanout (
		.a(G4),
		.b(new_net_1101),
		.c(new_net_1100)
	);

	spl4L G14_v_fanout (
		.a(G14),
		.b(new_net_1128),
		.c(new_net_850),
		.d(new_net_842),
		.e(new_net_849)
	);

	bfr new_net_2539_bfr_after (
		.din(G30),
		.dout(new_net_2539)
	);

	spl4L G30_v_fanout (
		.a(new_net_2539),
		.b(new_net_1143),
		.c(new_net_88),
		.d(new_net_83),
		.e(new_net_86)
	);

	bfr new_net_2540_bfr_after (
		.din(G21),
		.dout(new_net_2540)
	);

	bfr new_net_2541_bfr_before (
		.din(new_net_2541),
		.dout(new_net_1055)
	);

	bfr new_net_2542_bfr_before (
		.din(new_net_2542),
		.dout(new_net_2541)
	);

	bfr new_net_2543_bfr_before (
		.din(new_net_2543),
		.dout(new_net_2542)
	);

	spl2 G21_v_fanout (
		.a(new_net_2540),
		.b(new_net_2543),
		.c(new_net_617)
	);

	bfr new_net_2544_bfr_before (
		.din(new_net_2544),
		.dout(new_net_1060)
	);

	spl2 G41_v_fanout (
		.a(G41),
		.b(new_net_1059),
		.c(new_net_2544)
	);

	bfr new_net_2545_bfr_before (
		.din(new_net_2545),
		.dout(new_net_1066)
	);

	bfr new_net_2546_bfr_before (
		.din(new_net_2546),
		.dout(new_net_2545)
	);

	bfr new_net_2547_bfr_before (
		.din(new_net_2547),
		.dout(new_net_2546)
	);

	bfr new_net_2548_bfr_before (
		.din(new_net_2548),
		.dout(new_net_2547)
	);

	bfr new_net_2549_bfr_before (
		.din(new_net_2549),
		.dout(new_net_2548)
	);

	bfr new_net_2550_bfr_before (
		.din(new_net_2550),
		.dout(new_net_2549)
	);

	bfr new_net_2551_bfr_before (
		.din(new_net_2551),
		.dout(new_net_2550)
	);

	bfr new_net_2552_bfr_before (
		.din(new_net_2552),
		.dout(new_net_2551)
	);

	bfr new_net_2553_bfr_before (
		.din(new_net_2553),
		.dout(new_net_2552)
	);

	bfr new_net_2554_bfr_before (
		.din(new_net_2554),
		.dout(new_net_2553)
	);

	bfr new_net_2555_bfr_before (
		.din(new_net_2555),
		.dout(new_net_2554)
	);

	bfr new_net_2556_bfr_before (
		.din(new_net_2556),
		.dout(new_net_2555)
	);

	bfr new_net_2557_bfr_before (
		.din(new_net_2557),
		.dout(new_net_2556)
	);

	bfr new_net_2558_bfr_before (
		.din(new_net_2558),
		.dout(new_net_2557)
	);

	bfr new_net_2559_bfr_before (
		.din(new_net_2559),
		.dout(new_net_2558)
	);

	bfr new_net_2560_bfr_before (
		.din(new_net_2560),
		.dout(new_net_2559)
	);

	bfr new_net_2561_bfr_before (
		.din(new_net_2561),
		.dout(new_net_2560)
	);

	bfr new_net_2562_bfr_before (
		.din(new_net_2562),
		.dout(new_net_2561)
	);

	bfr new_net_2563_bfr_before (
		.din(new_net_2563),
		.dout(new_net_2562)
	);

	spl2 G47_v_fanout (
		.a(G47),
		.b(new_net_2563),
		.c(new_net_994)
	);

	spl2 G7_v_fanout (
		.a(G7),
		.b(new_net_1071),
		.c(new_net_1072)
	);

	bfr new_net_2564_bfr_before (
		.din(new_net_2564),
		.dout(new_net_1075)
	);

	bfr new_net_2565_bfr_before (
		.din(new_net_2565),
		.dout(new_net_2564)
	);

	spl2 G39_v_fanout (
		.a(G39),
		.b(new_net_1076),
		.c(new_net_2565)
	);

	bfr new_net_2566_bfr_before (
		.din(new_net_2566),
		.dout(new_net_243)
	);

	bfr new_net_2567_bfr_before (
		.din(new_net_2567),
		.dout(new_net_2566)
	);

	spl2 G33_v_fanout (
		.a(G33),
		.b(new_net_1077),
		.c(new_net_2567)
	);

	bfr new_net_2568_bfr_before (
		.din(new_net_2568),
		.dout(new_net_45)
	);

	bfr new_net_2569_bfr_before (
		.din(new_net_2569),
		.dout(new_net_2568)
	);

	bfr new_net_2570_bfr_before (
		.din(new_net_2570),
		.dout(new_net_2569)
	);

	bfr new_net_2571_bfr_before (
		.din(new_net_2571),
		.dout(new_net_2570)
	);

	bfr new_net_2572_bfr_before (
		.din(new_net_2572),
		.dout(new_net_2571)
	);

	bfr new_net_2573_bfr_before (
		.din(new_net_2573),
		.dout(new_net_2572)
	);

	bfr new_net_2574_bfr_before (
		.din(new_net_2574),
		.dout(new_net_2573)
	);

	bfr new_net_2575_bfr_before (
		.din(new_net_2575),
		.dout(new_net_2574)
	);

	bfr new_net_2576_bfr_before (
		.din(new_net_2576),
		.dout(new_net_2575)
	);

	bfr new_net_2577_bfr_before (
		.din(new_net_2577),
		.dout(new_net_2576)
	);

	bfr new_net_2578_bfr_before (
		.din(new_net_2578),
		.dout(new_net_2577)
	);

	bfr new_net_2579_bfr_before (
		.din(new_net_2579),
		.dout(new_net_2578)
	);

	bfr new_net_2580_bfr_before (
		.din(new_net_2580),
		.dout(new_net_2579)
	);

	bfr new_net_2581_bfr_before (
		.din(new_net_2581),
		.dout(new_net_2580)
	);

	bfr new_net_2582_bfr_before (
		.din(new_net_2582),
		.dout(new_net_2581)
	);

	bfr new_net_2583_bfr_before (
		.din(new_net_2583),
		.dout(new_net_2582)
	);

	bfr new_net_2584_bfr_before (
		.din(new_net_2584),
		.dout(new_net_2583)
	);

	bfr new_net_2585_bfr_before (
		.din(new_net_2585),
		.dout(new_net_2584)
	);

	bfr new_net_2586_bfr_before (
		.din(new_net_2586),
		.dout(new_net_2585)
	);

	bfr new_net_2587_bfr_before (
		.din(new_net_2587),
		.dout(new_net_2586)
	);

	bfr new_net_2588_bfr_before (
		.din(new_net_2588),
		.dout(new_net_2587)
	);

	bfr new_net_2589_bfr_before (
		.din(new_net_2589),
		.dout(new_net_2588)
	);

	bfr new_net_2590_bfr_before (
		.din(new_net_2590),
		.dout(new_net_2589)
	);

	bfr new_net_2591_bfr_before (
		.din(new_net_2591),
		.dout(new_net_2590)
	);

	bfr new_net_2592_bfr_before (
		.din(new_net_2592),
		.dout(new_net_2591)
	);

	bfr new_net_2593_bfr_before (
		.din(new_net_2593),
		.dout(new_net_2592)
	);

	bfr new_net_2594_bfr_before (
		.din(new_net_2594),
		.dout(new_net_2593)
	);

	bfr new_net_2595_bfr_before (
		.din(new_net_2595),
		.dout(new_net_2594)
	);

	bfr new_net_2596_bfr_before (
		.din(new_net_2596),
		.dout(new_net_2595)
	);

	bfr new_net_2597_bfr_before (
		.din(new_net_2597),
		.dout(new_net_2596)
	);

	bfr new_net_2598_bfr_before (
		.din(new_net_2598),
		.dout(new_net_2597)
	);

	bfr new_net_2599_bfr_before (
		.din(new_net_2599),
		.dout(new_net_2598)
	);

	bfr new_net_2600_bfr_before (
		.din(new_net_2600),
		.dout(new_net_2599)
	);

	bfr new_net_2601_bfr_before (
		.din(new_net_2601),
		.dout(new_net_2600)
	);

	bfr new_net_2602_bfr_before (
		.din(new_net_2602),
		.dout(new_net_2601)
	);

	bfr new_net_2603_bfr_before (
		.din(new_net_2603),
		.dout(new_net_2602)
	);

	bfr new_net_2604_bfr_before (
		.din(new_net_2604),
		.dout(new_net_2603)
	);

	bfr new_net_2605_bfr_before (
		.din(new_net_2605),
		.dout(new_net_2604)
	);

	bfr new_net_2606_bfr_before (
		.din(new_net_2606),
		.dout(new_net_2605)
	);

	bfr new_net_2607_bfr_before (
		.din(new_net_2607),
		.dout(new_net_2606)
	);

	bfr new_net_2608_bfr_before (
		.din(new_net_2608),
		.dout(new_net_2607)
	);

	bfr new_net_2609_bfr_before (
		.din(new_net_2609),
		.dout(new_net_2608)
	);

	bfr new_net_2610_bfr_before (
		.din(new_net_2610),
		.dout(new_net_2609)
	);

	bfr new_net_2611_bfr_before (
		.din(new_net_2611),
		.dout(new_net_2610)
	);

	bfr new_net_2612_bfr_before (
		.din(new_net_2612),
		.dout(new_net_2611)
	);

	bfr new_net_2613_bfr_before (
		.din(new_net_2613),
		.dout(new_net_2612)
	);

	spl2 G48_v_fanout (
		.a(G48),
		.b(new_net_2613),
		.c(new_net_44)
	);

	bfr new_net_2614_bfr_before (
		.din(new_net_2614),
		.dout(new_net_1086)
	);

	bfr new_net_2615_bfr_before (
		.din(new_net_2615),
		.dout(new_net_2614)
	);

	bfr new_net_2616_bfr_before (
		.din(new_net_2616),
		.dout(new_net_2615)
	);

	bfr new_net_2617_bfr_before (
		.din(new_net_2617),
		.dout(new_net_2616)
	);

	bfr new_net_2618_bfr_before (
		.din(new_net_2618),
		.dout(new_net_2617)
	);

	spl2 G27_v_fanout (
		.a(G27),
		.b(new_net_2618),
		.c(new_net_111)
	);

	bfr new_net_2619_bfr_before (
		.din(new_net_2619),
		.dout(new_net_1089)
	);

	bfr new_net_2620_bfr_before (
		.din(new_net_2620),
		.dout(new_net_2619)
	);

	bfr new_net_2621_bfr_before (
		.din(new_net_2621),
		.dout(new_net_2620)
	);

	bfr new_net_2622_bfr_before (
		.din(new_net_2622),
		.dout(new_net_2621)
	);

	bfr new_net_2623_bfr_before (
		.din(new_net_2623),
		.dout(new_net_2622)
	);

	bfr new_net_2624_bfr_before (
		.din(new_net_2624),
		.dout(new_net_2623)
	);

	bfr new_net_2625_bfr_before (
		.din(new_net_2625),
		.dout(new_net_2624)
	);

	spl3L G42_v_fanout (
		.a(G42),
		.b(new_net_2625),
		.c(new_net_758),
		.d(new_net_755)
	);

	bfr new_net_2626_bfr_after (
		.din(G43),
		.dout(new_net_2626)
	);

	bfr new_net_2627_bfr_before (
		.din(new_net_2627),
		.dout(new_net_1102)
	);

	bfr new_net_2628_bfr_before (
		.din(new_net_2628),
		.dout(new_net_2627)
	);

	bfr new_net_2629_bfr_before (
		.din(new_net_2629),
		.dout(new_net_2628)
	);

	bfr new_net_2630_bfr_before (
		.din(new_net_2630),
		.dout(new_net_2629)
	);

	bfr new_net_2631_bfr_before (
		.din(new_net_2631),
		.dout(new_net_2630)
	);

	bfr new_net_2632_bfr_before (
		.din(new_net_2632),
		.dout(new_net_2631)
	);

	spl2 G43_v_fanout (
		.a(new_net_2626),
		.b(new_net_2632),
		.c(new_net_64)
	);

	bfr new_net_2633_bfr_after (
		.din(G29),
		.dout(new_net_2633)
	);

	bfr new_net_2634_bfr_after (
		.din(new_net_2633),
		.dout(new_net_2634)
	);

	bfr new_net_2635_bfr_before (
		.din(new_net_2635),
		.dout(new_net_603)
	);

	bfr new_net_2636_bfr_before (
		.din(new_net_2636),
		.dout(new_net_2635)
	);

	bfr new_net_2637_bfr_before (
		.din(new_net_2637),
		.dout(new_net_2636)
	);

	spl2 G29_v_fanout (
		.a(new_net_2634),
		.b(new_net_2637),
		.c(new_net_602)
	);

	spl3L G3_v_fanout (
		.a(G3),
		.b(new_net_1106),
		.c(new_net_1105),
		.d(new_net_1107)
	);

	spl2 G24_v_fanout (
		.a(G24),
		.b(new_net_1117),
		.c(new_net_419)
	);

	bfr new_net_2638_bfr_before (
		.din(new_net_2638),
		.dout(new_net_790)
	);

	bfr new_net_2639_bfr_before (
		.din(new_net_2639),
		.dout(new_net_794)
	);

	spl3L G35_v_fanout (
		.a(G35),
		.b(new_net_1122),
		.c(new_net_2639),
		.d(new_net_2638)
	);

	spl2 G34_v_fanout (
		.a(G34),
		.b(new_net_1146),
		.c(new_net_1147)
	);

	spl2 G32_v_fanout (
		.a(G32),
		.b(new_net_1049),
		.c(new_net_1048)
	);

	bfr new_net_2640_bfr_before (
		.din(new_net_2640),
		.dout(new_net_204)
	);

	spl2 G23_v_fanout (
		.a(G23),
		.b(new_net_2640),
		.c(new_net_203)
	);

	bfr new_net_2641_bfr_before (
		.din(new_net_2641),
		.dout(new_net_1061)
	);

	bfr new_net_2642_bfr_before (
		.din(new_net_2642),
		.dout(new_net_2641)
	);

	bfr new_net_2643_bfr_before (
		.din(new_net_2643),
		.dout(new_net_2642)
	);

	bfr new_net_2644_bfr_before (
		.din(new_net_2644),
		.dout(new_net_2643)
	);

	bfr new_net_2645_bfr_before (
		.din(new_net_2645),
		.dout(new_net_2644)
	);

	bfr new_net_2646_bfr_before (
		.din(new_net_2646),
		.dout(new_net_2645)
	);

	bfr new_net_2647_bfr_before (
		.din(new_net_2647),
		.dout(new_net_2646)
	);

	spl2 G18_v_fanout (
		.a(G18),
		.b(new_net_2647),
		.c(new_net_403)
	);

	bfr new_net_2648_bfr_before (
		.din(new_net_2648),
		.dout(new_net_1087)
	);

	bfr new_net_2649_bfr_before (
		.din(new_net_2649),
		.dout(new_net_2648)
	);

	bfr new_net_2650_bfr_before (
		.din(new_net_2650),
		.dout(new_net_128)
	);

	bfr new_net_2651_bfr_before (
		.din(new_net_2651),
		.dout(new_net_2650)
	);

	spl4L G5_v_fanout (
		.a(G5),
		.b(new_net_127),
		.c(new_net_2651),
		.d(new_net_2649),
		.e(new_net_129)
	);

	spl2 G12_v_fanout (
		.a(G12),
		.b(new_net_1109),
		.c(new_net_1110)
	);

	bfr new_net_2652_bfr_before (
		.din(new_net_2652),
		.dout(new_net_1111)
	);

	bfr new_net_2653_bfr_before (
		.din(new_net_2653),
		.dout(new_net_2652)
	);

	bfr new_net_2654_bfr_before (
		.din(new_net_2654),
		.dout(new_net_2653)
	);

	bfr new_net_2655_bfr_before (
		.din(new_net_2655),
		.dout(new_net_2654)
	);

	bfr new_net_2656_bfr_before (
		.din(new_net_2656),
		.dout(new_net_2655)
	);

	bfr new_net_2657_bfr_before (
		.din(new_net_2657),
		.dout(new_net_2656)
	);

	bfr new_net_2658_bfr_before (
		.din(new_net_2658),
		.dout(new_net_2657)
	);

	spl2 G44_v_fanout (
		.a(G44),
		.b(new_net_2658),
		.c(new_net_851)
	);

	bfr new_net_2659_bfr_before (
		.din(new_net_2659),
		.dout(new_net_59)
	);

	spl4L G11_v_fanout (
		.a(G11),
		.b(new_net_1112),
		.c(new_net_1116),
		.d(new_net_52),
		.e(new_net_2659)
	);

	spl2 G19_v_fanout (
		.a(G19),
		.b(new_net_1120),
		.c(new_net_443)
	);

	bfr new_net_2660_bfr_after (
		.din(G20),
		.dout(new_net_2660)
	);

	bfr new_net_2661_bfr_after (
		.din(new_net_2660),
		.dout(new_net_2661)
	);

	bfr new_net_2662_bfr_after (
		.din(new_net_2661),
		.dout(new_net_2662)
	);

	bfr new_net_2663_bfr_after (
		.din(new_net_2662),
		.dout(new_net_2663)
	);

	bfr new_net_2664_bfr_after (
		.din(new_net_2663),
		.dout(new_net_2664)
	);

	bfr new_net_2665_bfr_after (
		.din(new_net_2664),
		.dout(new_net_2665)
	);

	bfr new_net_2666_bfr_after (
		.din(new_net_2665),
		.dout(new_net_2666)
	);

	bfr new_net_2667_bfr_before (
		.din(new_net_2667),
		.dout(new_net_1131)
	);

	spl2 G20_v_fanout (
		.a(new_net_2666),
		.b(new_net_2667),
		.c(new_net_1130)
	);

	spl2 G1_v_fanout (
		.a(G1),
		.b(new_net_1136),
		.c(new_net_1135)
	);

	bfr new_net_2668_bfr_after (
		.din(G2),
		.dout(new_net_2668)
	);

	spl4L G2_v_fanout (
		.a(new_net_2668),
		.b(new_net_1137),
		.c(new_net_496),
		.d(new_net_491),
		.e(new_net_494)
	);

	spl2 G31_v_fanout (
		.a(G31),
		.b(new_net_1051),
		.c(new_net_1052)
	);

	spl2 G36_v_fanout (
		.a(G36),
		.b(new_net_1054),
		.c(new_net_1053)
	);

	bfr new_net_2669_bfr_after (
		.din(G17),
		.dout(new_net_2669)
	);

	bfr new_net_2670_bfr_after (
		.din(new_net_2669),
		.dout(new_net_2670)
	);

	bfr new_net_2671_bfr_after (
		.din(new_net_2670),
		.dout(new_net_2671)
	);

	bfr new_net_2672_bfr_after (
		.din(new_net_2671),
		.dout(new_net_2672)
	);

	bfr new_net_2673_bfr_after (
		.din(new_net_2672),
		.dout(new_net_2673)
	);

	bfr new_net_2674_bfr_after (
		.din(new_net_2673),
		.dout(new_net_2674)
	);

	bfr new_net_2675_bfr_after (
		.din(new_net_2674),
		.dout(new_net_2675)
	);

	bfr new_net_2676_bfr_after (
		.din(new_net_2675),
		.dout(new_net_2676)
	);

	bfr new_net_2677_bfr_before (
		.din(new_net_2677),
		.dout(new_net_355)
	);

	bfr new_net_2678_bfr_before (
		.din(new_net_2678),
		.dout(new_net_356)
	);

	spl3L G17_v_fanout (
		.a(new_net_2676),
		.b(new_net_2678),
		.c(new_net_357),
		.d(new_net_2677)
	);

	bfr new_net_2679_bfr_before (
		.din(new_net_2679),
		.dout(new_net_805)
	);

	spl2 G25_v_fanout (
		.a(G25),
		.b(new_net_2679),
		.c(new_net_804)
	);

	bfr new_net_2680_bfr_before (
		.din(new_net_2680),
		.dout(new_net_14)
	);

	bfr new_net_2681_bfr_before (
		.din(new_net_2681),
		.dout(new_net_18)
	);

	spl4L G8_v_fanout (
		.a(G8),
		.b(new_net_17),
		.c(new_net_2681),
		.d(new_net_1062),
		.e(new_net_2680)
	);

	spl2 G13_v_fanout (
		.a(G13),
		.b(new_net_1082),
		.c(new_net_1081)
	);

	spl2 G9_v_fanout (
		.a(G9),
		.b(new_net_1085),
		.c(new_net_1084)
	);

	bfr new_net_2682_bfr_before (
		.din(new_net_2682),
		.dout(new_net_249)
	);

	bfr new_net_2683_bfr_before (
		.din(new_net_2683),
		.dout(new_net_248)
	);

	bfr new_net_2684_bfr_before (
		.din(new_net_2684),
		.dout(new_net_2683)
	);

	bfr new_net_2685_bfr_before (
		.din(new_net_2685),
		.dout(new_net_2684)
	);

	bfr new_net_2686_bfr_before (
		.din(new_net_2686),
		.dout(new_net_2685)
	);

	bfr new_net_2687_bfr_before (
		.din(new_net_2687),
		.dout(new_net_2686)
	);

	bfr new_net_2688_bfr_before (
		.din(new_net_2688),
		.dout(new_net_2687)
	);

	bfr new_net_2689_bfr_before (
		.din(new_net_2689),
		.dout(new_net_2688)
	);

	bfr new_net_2690_bfr_before (
		.din(new_net_2690),
		.dout(new_net_2689)
	);

	bfr new_net_2691_bfr_before (
		.din(new_net_2691),
		.dout(new_net_247)
	);

	spl4L G6_v_fanout (
		.a(G6),
		.b(new_net_2691),
		.c(new_net_2690),
		.d(new_net_246),
		.e(new_net_2682)
	);

	bfr new_net_2692_bfr_before (
		.din(new_net_2692),
		.dout(new_net_1088)
	);

	bfr new_net_2693_bfr_before (
		.din(new_net_2693),
		.dout(new_net_2692)
	);

	spl2 G26_v_fanout (
		.a(G26),
		.b(new_net_2693),
		.c(new_net_859)
	);

	spl2 G22_v_fanout (
		.a(G22),
		.b(new_net_1125),
		.c(new_net_674)
	);

	spl2 G40_v_fanout (
		.a(G40),
		.b(new_net_386),
		.c(new_net_1139)
	);

	bfr new_net_2694_bfr_after (
		.din(_0557_),
		.dout(new_net_2694)
	);

	bfr new_net_2695_bfr_after (
		.din(new_net_2694),
		.dout(new_net_2695)
	);

	bfr new_net_2696_bfr_after (
		.din(new_net_2695),
		.dout(new_net_2696)
	);

	bfr new_net_2697_bfr_after (
		.din(new_net_2696),
		.dout(new_net_2697)
	);

	bfr new_net_2698_bfr_after (
		.din(new_net_2697),
		.dout(new_net_2698)
	);

	bfr new_net_1391_bfr_after (
		.din(new_net_2698),
		.dout(new_net_1391)
	);

	bfr new_net_2699_bfr_after (
		.din(_0475_),
		.dout(new_net_2699)
	);

	bfr new_net_2700_bfr_after (
		.din(new_net_2699),
		.dout(new_net_2700)
	);

	bfr new_net_2701_bfr_after (
		.din(new_net_2700),
		.dout(new_net_2701)
	);

	bfr new_net_2702_bfr_after (
		.din(new_net_2701),
		.dout(new_net_2702)
	);

	bfr new_net_2703_bfr_after (
		.din(new_net_2702),
		.dout(new_net_2703)
	);

	bfr new_net_1365_bfr_after (
		.din(new_net_2703),
		.dout(new_net_1365)
	);

	bfr new_net_1257_bfr_after (
		.din(_0788_),
		.dout(new_net_1257)
	);

	bfr new_net_1413_bfr_after (
		.din(_0632_),
		.dout(new_net_1413)
	);

	bfr new_net_1387_bfr_after (
		.din(_0534_),
		.dout(new_net_1387)
	);

	bfr new_net_2704_bfr_after (
		.din(new_net_1465),
		.dout(new_net_2704)
	);

	bfr new_net_2705_bfr_after (
		.din(new_net_2704),
		.dout(new_net_2705)
	);

	bfr new_net_2706_bfr_after (
		.din(new_net_2705),
		.dout(new_net_2706)
	);

	bfr new_net_2707_bfr_after (
		.din(new_net_2706),
		.dout(new_net_2707)
	);

	bfr new_net_2708_bfr_after (
		.din(new_net_2707),
		.dout(new_net_2708)
	);

	bfr new_net_2709_bfr_after (
		.din(new_net_2708),
		.dout(new_net_2709)
	);

	bfr new_net_2710_bfr_after (
		.din(new_net_2709),
		.dout(new_net_2710)
	);

	bfr new_net_2711_bfr_after (
		.din(new_net_2710),
		.dout(new_net_2711)
	);

	bfr new_net_2712_bfr_after (
		.din(new_net_2711),
		.dout(new_net_2712)
	);

	bfr new_net_2713_bfr_after (
		.din(new_net_2712),
		.dout(new_net_2713)
	);

	bfr new_net_2714_bfr_after (
		.din(new_net_2713),
		.dout(new_net_2714)
	);

	bfr new_net_2715_bfr_after (
		.din(new_net_2714),
		.dout(new_net_2715)
	);

	bfr new_net_2716_bfr_after (
		.din(new_net_2715),
		.dout(new_net_2716)
	);

	bfr new_net_2717_bfr_after (
		.din(new_net_2716),
		.dout(new_net_2717)
	);

	bfr new_net_2718_bfr_after (
		.din(new_net_2717),
		.dout(new_net_2718)
	);

	bfr new_net_2719_bfr_after (
		.din(new_net_2718),
		.dout(new_net_2719)
	);

	bfr new_net_2720_bfr_after (
		.din(new_net_2719),
		.dout(new_net_2720)
	);

	bfr new_net_2721_bfr_after (
		.din(new_net_2720),
		.dout(new_net_2721)
	);

	bfr new_net_2722_bfr_after (
		.din(new_net_2721),
		.dout(new_net_2722)
	);

	bfr new_net_2723_bfr_after (
		.din(new_net_2722),
		.dout(new_net_2723)
	);

	bfr new_net_2724_bfr_after (
		.din(new_net_2723),
		.dout(new_net_2724)
	);

	bfr new_net_2725_bfr_after (
		.din(new_net_2724),
		.dout(new_net_2725)
	);

	bfr new_net_2726_bfr_after (
		.din(new_net_2725),
		.dout(new_net_2726)
	);

	bfr new_net_2727_bfr_after (
		.din(new_net_2726),
		.dout(new_net_2727)
	);

	bfr new_net_2728_bfr_after (
		.din(new_net_2727),
		.dout(new_net_2728)
	);

	bfr new_net_2729_bfr_after (
		.din(new_net_2728),
		.dout(new_net_2729)
	);

	bfr new_net_2730_bfr_after (
		.din(new_net_2729),
		.dout(new_net_2730)
	);

	bfr G3525_bfr_after (
		.din(new_net_2730),
		.dout(G3525)
	);

	bfr new_net_2731_bfr_after (
		.din(new_net_1477),
		.dout(new_net_2731)
	);

	bfr new_net_2732_bfr_after (
		.din(new_net_2731),
		.dout(new_net_2732)
	);

	bfr new_net_2733_bfr_after (
		.din(new_net_2732),
		.dout(new_net_2733)
	);

	bfr new_net_2734_bfr_after (
		.din(new_net_2733),
		.dout(new_net_2734)
	);

	bfr new_net_2735_bfr_after (
		.din(new_net_2734),
		.dout(new_net_2735)
	);

	bfr new_net_2736_bfr_after (
		.din(new_net_2735),
		.dout(new_net_2736)
	);

	bfr new_net_2737_bfr_after (
		.din(new_net_2736),
		.dout(new_net_2737)
	);

	bfr new_net_2738_bfr_after (
		.din(new_net_2737),
		.dout(new_net_2738)
	);

	bfr new_net_2739_bfr_after (
		.din(new_net_2738),
		.dout(new_net_2739)
	);

	bfr new_net_2740_bfr_after (
		.din(new_net_2739),
		.dout(new_net_2740)
	);

	bfr new_net_2741_bfr_after (
		.din(new_net_2740),
		.dout(new_net_2741)
	);

	bfr new_net_2742_bfr_after (
		.din(new_net_2741),
		.dout(new_net_2742)
	);

	bfr new_net_2743_bfr_after (
		.din(new_net_2742),
		.dout(new_net_2743)
	);

	bfr new_net_2744_bfr_after (
		.din(new_net_2743),
		.dout(new_net_2744)
	);

	bfr new_net_2745_bfr_after (
		.din(new_net_2744),
		.dout(new_net_2745)
	);

	bfr new_net_2746_bfr_after (
		.din(new_net_2745),
		.dout(new_net_2746)
	);

	bfr new_net_2747_bfr_after (
		.din(new_net_2746),
		.dout(new_net_2747)
	);

	bfr new_net_2748_bfr_after (
		.din(new_net_2747),
		.dout(new_net_2748)
	);

	bfr new_net_2749_bfr_after (
		.din(new_net_2748),
		.dout(new_net_2749)
	);

	bfr new_net_2750_bfr_after (
		.din(new_net_2749),
		.dout(new_net_2750)
	);

	bfr new_net_2751_bfr_after (
		.din(new_net_2750),
		.dout(new_net_2751)
	);

	bfr new_net_2752_bfr_after (
		.din(new_net_2751),
		.dout(new_net_2752)
	);

	bfr new_net_2753_bfr_after (
		.din(new_net_2752),
		.dout(new_net_2753)
	);

	bfr new_net_2754_bfr_after (
		.din(new_net_2753),
		.dout(new_net_2754)
	);

	bfr new_net_2755_bfr_after (
		.din(new_net_2754),
		.dout(new_net_2755)
	);

	bfr new_net_2756_bfr_after (
		.din(new_net_2755),
		.dout(new_net_2756)
	);

	bfr new_net_2757_bfr_after (
		.din(new_net_2756),
		.dout(new_net_2757)
	);

	bfr new_net_2758_bfr_after (
		.din(new_net_2757),
		.dout(new_net_2758)
	);

	bfr new_net_2759_bfr_after (
		.din(new_net_2758),
		.dout(new_net_2759)
	);

	bfr new_net_2760_bfr_after (
		.din(new_net_2759),
		.dout(new_net_2760)
	);

	bfr new_net_2761_bfr_after (
		.din(new_net_2760),
		.dout(new_net_2761)
	);

	bfr new_net_2762_bfr_after (
		.din(new_net_2761),
		.dout(new_net_2762)
	);

	bfr new_net_2763_bfr_after (
		.din(new_net_2762),
		.dout(new_net_2763)
	);

	bfr new_net_2764_bfr_after (
		.din(new_net_2763),
		.dout(new_net_2764)
	);

	bfr new_net_2765_bfr_after (
		.din(new_net_2764),
		.dout(new_net_2765)
	);

	bfr new_net_2766_bfr_after (
		.din(new_net_2765),
		.dout(new_net_2766)
	);

	bfr new_net_2767_bfr_after (
		.din(new_net_2766),
		.dout(new_net_2767)
	);

	bfr new_net_2768_bfr_after (
		.din(new_net_2767),
		.dout(new_net_2768)
	);

	bfr new_net_2769_bfr_after (
		.din(new_net_2768),
		.dout(new_net_2769)
	);

	bfr new_net_2770_bfr_after (
		.din(new_net_2769),
		.dout(new_net_2770)
	);

	bfr new_net_2771_bfr_after (
		.din(new_net_2770),
		.dout(new_net_2771)
	);

	bfr new_net_2772_bfr_after (
		.din(new_net_2771),
		.dout(new_net_2772)
	);

	bfr new_net_2773_bfr_after (
		.din(new_net_2772),
		.dout(new_net_2773)
	);

	bfr new_net_2774_bfr_after (
		.din(new_net_2773),
		.dout(new_net_2774)
	);

	bfr G3522_bfr_after (
		.din(new_net_2774),
		.dout(G3522)
	);

	bfr new_net_1351_bfr_after (
		.din(_0421_),
		.dout(new_net_1351)
	);

	bfr new_net_2775_bfr_after (
		.din(_0679_),
		.dout(new_net_2775)
	);

	bfr new_net_2776_bfr_after (
		.din(new_net_2775),
		.dout(new_net_2776)
	);

	bfr new_net_1435_bfr_after (
		.din(new_net_2776),
		.dout(new_net_1435)
	);

	bfr new_net_2777_bfr_after (
		.din(_0409_),
		.dout(new_net_2777)
	);

	bfr new_net_2778_bfr_after (
		.din(new_net_2777),
		.dout(new_net_2778)
	);

	bfr new_net_2779_bfr_after (
		.din(new_net_2778),
		.dout(new_net_2779)
	);

	bfr new_net_2780_bfr_after (
		.din(new_net_2779),
		.dout(new_net_2780)
	);

	bfr new_net_2781_bfr_after (
		.din(new_net_2780),
		.dout(new_net_2781)
	);

	bfr new_net_2782_bfr_after (
		.din(new_net_2781),
		.dout(new_net_2782)
	);

	bfr new_net_2783_bfr_after (
		.din(new_net_2782),
		.dout(new_net_2783)
	);

	bfr new_net_2784_bfr_after (
		.din(new_net_2783),
		.dout(new_net_2784)
	);

	bfr new_net_2785_bfr_after (
		.din(new_net_2784),
		.dout(new_net_2785)
	);

	bfr new_net_2786_bfr_after (
		.din(new_net_2785),
		.dout(new_net_2786)
	);

	bfr new_net_2787_bfr_after (
		.din(new_net_2786),
		.dout(new_net_2787)
	);

	bfr new_net_2788_bfr_after (
		.din(new_net_2787),
		.dout(new_net_2788)
	);

	bfr new_net_2789_bfr_after (
		.din(new_net_2788),
		.dout(new_net_2789)
	);

	bfr new_net_2790_bfr_after (
		.din(new_net_2789),
		.dout(new_net_2790)
	);

	bfr new_net_2791_bfr_after (
		.din(new_net_2790),
		.dout(new_net_2791)
	);

	bfr new_net_2792_bfr_after (
		.din(new_net_2791),
		.dout(new_net_2792)
	);

	bfr new_net_2793_bfr_after (
		.din(new_net_2792),
		.dout(new_net_2793)
	);

	bfr new_net_2794_bfr_after (
		.din(new_net_2793),
		.dout(new_net_2794)
	);

	bfr new_net_1346_bfr_after (
		.din(new_net_2794),
		.dout(new_net_1346)
	);

	bfr new_net_1409_bfr_after (
		.din(_0574_),
		.dout(new_net_1409)
	);

	bfr new_net_2795_bfr_after (
		.din(_0120_),
		.dout(new_net_2795)
	);

	bfr new_net_1282_bfr_after (
		.din(new_net_2795),
		.dout(new_net_1282)
	);

	bfr new_net_2796_bfr_after (
		.din(_0201_),
		.dout(new_net_2796)
	);

	bfr new_net_2797_bfr_after (
		.din(new_net_2796),
		.dout(new_net_2797)
	);

	bfr new_net_1303_bfr_after (
		.din(new_net_2797),
		.dout(new_net_1303)
	);

	bfr new_net_2798_bfr_after (
		.din(_0280_),
		.dout(new_net_2798)
	);

	bfr new_net_1324_bfr_after (
		.din(new_net_2798),
		.dout(new_net_1324)
	);

	bfr new_net_1261_bfr_after (
		.din(_0790_),
		.dout(new_net_1261)
	);

	bfr new_net_2799_bfr_after (
		.din(_0096_),
		.dout(new_net_2799)
	);

	bfr new_net_1274_bfr_after (
		.din(new_net_2799),
		.dout(new_net_1274)
	);

	bfr new_net_1278_bfr_after (
		.din(_0101_),
		.dout(new_net_1278)
	);

	bfr new_net_2800_bfr_after (
		.din(_0170_),
		.dout(new_net_2800)
	);

	bfr new_net_1295_bfr_after (
		.din(new_net_2800),
		.dout(new_net_1295)
	);

	bfr new_net_1316_bfr_after (
		.din(_0237_),
		.dout(new_net_1316)
	);

	bfr new_net_2801_bfr_after (
		.din(_0187_),
		.dout(new_net_2801)
	);

	bfr new_net_1299_bfr_after (
		.din(new_net_2801),
		.dout(new_net_1299)
	);

	bfr new_net_1320_bfr_after (
		.din(_0264_),
		.dout(new_net_1320)
	);

	bfr new_net_2802_bfr_after (
		.din(_0496_),
		.dout(new_net_2802)
	);

	bfr new_net_2803_bfr_after (
		.din(new_net_2802),
		.dout(new_net_2803)
	);

	bfr new_net_1373_bfr_after (
		.din(new_net_2803),
		.dout(new_net_1373)
	);

	bfr new_net_1378_bfr_after (
		.din(_0508_),
		.dout(new_net_1378)
	);

	bfr new_net_2804_bfr_after (
		.din(_0761_),
		.dout(new_net_2804)
	);

	bfr new_net_2805_bfr_after (
		.din(new_net_2804),
		.dout(new_net_2805)
	);

	bfr new_net_1457_bfr_after (
		.din(new_net_2805),
		.dout(new_net_1457)
	);

	bfr new_net_2806_bfr_after (
		.din(_0366_),
		.dout(new_net_2806)
	);

	bfr new_net_2807_bfr_after (
		.din(new_net_2806),
		.dout(new_net_2807)
	);

	bfr new_net_2808_bfr_after (
		.din(new_net_2807),
		.dout(new_net_2808)
	);

	bfr new_net_1337_bfr_after (
		.din(new_net_2808),
		.dout(new_net_1337)
	);

	bfr new_net_2809_bfr_after (
		.din(_0582_),
		.dout(new_net_2809)
	);

	bfr new_net_1400_bfr_after (
		.din(new_net_2809),
		.dout(new_net_1400)
	);

	bfr new_net_2810_bfr_after (
		.din(_0573_),
		.dout(new_net_2810)
	);

	bfr new_net_1395_bfr_after (
		.din(new_net_2810),
		.dout(new_net_1395)
	);

	bfr new_net_2811_bfr_after (
		.din(_0660_),
		.dout(new_net_2811)
	);

	bfr new_net_1422_bfr_after (
		.din(new_net_2811),
		.dout(new_net_1422)
	);

	bfr new_net_1443_bfr_after (
		.din(_0715_),
		.dout(new_net_1443)
	);

	bfr new_net_1260_bfr_after (
		.din(_0797_),
		.dout(new_net_1260)
	);

	bfr new_net_1417_bfr_after (
		.din(_0646_),
		.dout(new_net_1417)
	);

	bfr new_net_1355_bfr_after (
		.din(_0435_),
		.dout(new_net_1355)
	);

	bfr new_net_2812_bfr_after (
		.din(_0702_),
		.dout(new_net_2812)
	);

	bfr new_net_2813_bfr_after (
		.din(new_net_2812),
		.dout(new_net_2813)
	);

	bfr new_net_1439_bfr_after (
		.din(new_net_2813),
		.dout(new_net_1439)
	);

	bfr new_net_2814_bfr_after (
		.din(_0515_),
		.dout(new_net_2814)
	);

	bfr new_net_1382_bfr_after (
		.din(new_net_2814),
		.dout(new_net_1382)
	);

	bfr new_net_2815_bfr_after (
		.din(_0497_),
		.dout(new_net_2815)
	);

	bfr new_net_2816_bfr_after (
		.din(new_net_2815),
		.dout(new_net_2816)
	);

	bfr new_net_2817_bfr_after (
		.din(new_net_2816),
		.dout(new_net_2817)
	);

	bfr new_net_2818_bfr_after (
		.din(new_net_2817),
		.dout(new_net_2818)
	);

	bfr new_net_2819_bfr_after (
		.din(new_net_2818),
		.dout(new_net_2819)
	);

	bfr new_net_2820_bfr_after (
		.din(new_net_2819),
		.dout(new_net_2820)
	);

	bfr new_net_2821_bfr_after (
		.din(new_net_2820),
		.dout(new_net_2821)
	);

	bfr new_net_2822_bfr_after (
		.din(new_net_2821),
		.dout(new_net_2822)
	);

	bfr new_net_2823_bfr_after (
		.din(new_net_2822),
		.dout(new_net_2823)
	);

	bfr new_net_2824_bfr_after (
		.din(new_net_2823),
		.dout(new_net_2824)
	);

	bfr new_net_1377_bfr_after (
		.din(new_net_2824),
		.dout(new_net_1377)
	);

	bfr new_net_2825_bfr_after (
		.din(_0780_),
		.dout(new_net_2825)
	);

	bfr new_net_2826_bfr_after (
		.din(new_net_2825),
		.dout(new_net_2826)
	);

	bfr new_net_2827_bfr_after (
		.din(new_net_2826),
		.dout(new_net_2827)
	);

	bfr new_net_2828_bfr_after (
		.din(new_net_2827),
		.dout(new_net_2828)
	);

	bfr new_net_2829_bfr_after (
		.din(new_net_2828),
		.dout(new_net_2829)
	);

	bfr new_net_2830_bfr_after (
		.din(new_net_2829),
		.dout(new_net_2830)
	);

	bfr new_net_2831_bfr_after (
		.din(new_net_2830),
		.dout(new_net_2831)
	);

	bfr new_net_2832_bfr_after (
		.din(new_net_2831),
		.dout(new_net_2832)
	);

	bfr new_net_2833_bfr_after (
		.din(new_net_2832),
		.dout(new_net_2833)
	);

	bfr new_net_2834_bfr_after (
		.din(new_net_2833),
		.dout(new_net_2834)
	);

	bfr new_net_2835_bfr_after (
		.din(new_net_2834),
		.dout(new_net_2835)
	);

	bfr new_net_2836_bfr_after (
		.din(new_net_2835),
		.dout(new_net_2836)
	);

	bfr new_net_2837_bfr_after (
		.din(new_net_2836),
		.dout(new_net_2837)
	);

	bfr new_net_2838_bfr_after (
		.din(new_net_2837),
		.dout(new_net_2838)
	);

	bfr new_net_2839_bfr_after (
		.din(new_net_2838),
		.dout(new_net_2839)
	);

	bfr new_net_2840_bfr_after (
		.din(new_net_2839),
		.dout(new_net_2840)
	);

	bfr new_net_2841_bfr_after (
		.din(new_net_2840),
		.dout(new_net_2841)
	);

	bfr new_net_2842_bfr_after (
		.din(new_net_2841),
		.dout(new_net_2842)
	);

	bfr new_net_2843_bfr_after (
		.din(new_net_2842),
		.dout(new_net_2843)
	);

	bfr new_net_2844_bfr_after (
		.din(new_net_2843),
		.dout(new_net_2844)
	);

	bfr new_net_2845_bfr_after (
		.din(new_net_2844),
		.dout(new_net_2845)
	);

	bfr new_net_2846_bfr_after (
		.din(new_net_2845),
		.dout(new_net_2846)
	);

	bfr new_net_2847_bfr_after (
		.din(new_net_2846),
		.dout(new_net_2847)
	);

	bfr new_net_2848_bfr_after (
		.din(new_net_2847),
		.dout(new_net_2848)
	);

	bfr new_net_2849_bfr_after (
		.din(new_net_2848),
		.dout(new_net_2849)
	);

	bfr new_net_1461_bfr_after (
		.din(new_net_2849),
		.dout(new_net_1461)
	);

	bfr new_net_1286_bfr_after (
		.din(_0137_),
		.dout(new_net_1286)
	);

	bfr new_net_1307_bfr_after (
		.din(_0211_),
		.dout(new_net_1307)
	);

	bfr new_net_1328_bfr_after (
		.din(_0299_),
		.dout(new_net_1328)
	);

	bfr new_net_2850_bfr_after (
		.din(G28),
		.dout(new_net_2850)
	);

	bfr new_net_2851_bfr_after (
		.din(new_net_2850),
		.dout(new_net_2851)
	);

	bfr new_net_2852_bfr_after (
		.din(new_net_2851),
		.dout(new_net_2852)
	);

	bfr new_net_2853_bfr_after (
		.din(new_net_2852),
		.dout(new_net_2853)
	);

	bfr new_net_2854_bfr_after (
		.din(new_net_2853),
		.dout(new_net_2854)
	);

	bfr new_net_1269_bfr_after (
		.din(new_net_2854),
		.dout(new_net_1269)
	);

	bfr new_net_1290_bfr_after (
		.din(_0155_),
		.dout(new_net_1290)
	);

	bfr new_net_1311_bfr_after (
		.din(_0222_),
		.dout(new_net_1311)
	);

	bfr new_net_1265_bfr_after (
		.din(_0058_),
		.dout(new_net_1265)
	);

	bfr new_net_2855_bfr_after (
		.din(_0324_),
		.dout(new_net_2855)
	);

	bfr new_net_2856_bfr_after (
		.din(new_net_2855),
		.dout(new_net_2856)
	);

	bfr new_net_2857_bfr_after (
		.din(new_net_2856),
		.dout(new_net_2857)
	);

	bfr new_net_2858_bfr_after (
		.din(new_net_2857),
		.dout(new_net_2858)
	);

	bfr new_net_1332_bfr_after (
		.din(new_net_2858),
		.dout(new_net_1332)
	);

	bfr new_net_2859_bfr_after (
		.din(_0391_),
		.dout(new_net_2859)
	);

	bfr new_net_2860_bfr_after (
		.din(new_net_2859),
		.dout(new_net_2860)
	);

	bfr new_net_1341_bfr_after (
		.din(new_net_2860),
		.dout(new_net_1341)
	);

	bfr new_net_1349_bfr_after (
		.din(G15),
		.dout(new_net_1349)
	);

	bfr new_net_2861_bfr_after (
		.din(_0599_),
		.dout(new_net_2861)
	);

	bfr new_net_2862_bfr_after (
		.din(new_net_2861),
		.dout(new_net_2862)
	);

	bfr new_net_1404_bfr_after (
		.din(new_net_2862),
		.dout(new_net_1404)
	);

	bfr new_net_2863_bfr_after (
		.din(_0470_),
		.dout(new_net_2863)
	);

	bfr new_net_1368_bfr_after (
		.din(new_net_2863),
		.dout(new_net_1368)
	);

	bfr new_net_1452_bfr_after (
		.din(_0739_),
		.dout(new_net_1452)
	);

	bfr new_net_2864_bfr_after (
		.din(_0669_),
		.dout(new_net_2864)
	);

	bfr new_net_1426_bfr_after (
		.din(new_net_2864),
		.dout(new_net_1426)
	);

	bfr new_net_2865_bfr_after (
		.din(_0729_),
		.dout(new_net_2865)
	);

	bfr new_net_1447_bfr_after (
		.din(new_net_2865),
		.dout(new_net_1447)
	);

	bfr new_net_2866_bfr_after (
		.din(_0540_),
		.dout(new_net_2866)
	);

	bfr new_net_2867_bfr_after (
		.din(new_net_2866),
		.dout(new_net_2867)
	);

	bfr new_net_1390_bfr_after (
		.din(new_net_2867),
		.dout(new_net_1390)
	);

	bfr new_net_2868_bfr_after (
		.din(new_net_1469),
		.dout(new_net_2868)
	);

	bfr G3540_bfr_after (
		.din(new_net_2868),
		.dout(G3540)
	);

	bfr new_net_2869_bfr_after (
		.din(new_net_1481),
		.dout(new_net_2869)
	);

	bfr new_net_2870_bfr_after (
		.din(new_net_2869),
		.dout(new_net_2870)
	);

	bfr new_net_2871_bfr_after (
		.din(new_net_2870),
		.dout(new_net_2871)
	);

	bfr new_net_2872_bfr_after (
		.din(new_net_2871),
		.dout(new_net_2872)
	);

	bfr new_net_2873_bfr_after (
		.din(new_net_2872),
		.dout(new_net_2873)
	);

	bfr new_net_2874_bfr_after (
		.din(new_net_2873),
		.dout(new_net_2874)
	);

	bfr new_net_2875_bfr_after (
		.din(new_net_2874),
		.dout(new_net_2875)
	);

	bfr new_net_2876_bfr_after (
		.din(new_net_2875),
		.dout(new_net_2876)
	);

	bfr new_net_2877_bfr_after (
		.din(new_net_2876),
		.dout(new_net_2877)
	);

	bfr new_net_2878_bfr_after (
		.din(new_net_2877),
		.dout(new_net_2878)
	);

	bfr new_net_2879_bfr_after (
		.din(new_net_2878),
		.dout(new_net_2879)
	);

	bfr new_net_2880_bfr_after (
		.din(new_net_2879),
		.dout(new_net_2880)
	);

	bfr new_net_2881_bfr_after (
		.din(new_net_2880),
		.dout(new_net_2881)
	);

	bfr new_net_2882_bfr_after (
		.din(new_net_2881),
		.dout(new_net_2882)
	);

	bfr new_net_2883_bfr_after (
		.din(new_net_2882),
		.dout(new_net_2883)
	);

	bfr new_net_2884_bfr_after (
		.din(new_net_2883),
		.dout(new_net_2884)
	);

	bfr new_net_2885_bfr_after (
		.din(new_net_2884),
		.dout(new_net_2885)
	);

	bfr new_net_2886_bfr_after (
		.din(new_net_2885),
		.dout(new_net_2886)
	);

	bfr new_net_2887_bfr_after (
		.din(new_net_2886),
		.dout(new_net_2887)
	);

	bfr new_net_2888_bfr_after (
		.din(new_net_2887),
		.dout(new_net_2888)
	);

	bfr new_net_2889_bfr_after (
		.din(new_net_2888),
		.dout(new_net_2889)
	);

	bfr new_net_2890_bfr_after (
		.din(new_net_2889),
		.dout(new_net_2890)
	);

	bfr new_net_2891_bfr_after (
		.din(new_net_2890),
		.dout(new_net_2891)
	);

	bfr new_net_2892_bfr_after (
		.din(new_net_2891),
		.dout(new_net_2892)
	);

	bfr new_net_2893_bfr_after (
		.din(new_net_2892),
		.dout(new_net_2893)
	);

	bfr new_net_2894_bfr_after (
		.din(new_net_2893),
		.dout(new_net_2894)
	);

	bfr new_net_2895_bfr_after (
		.din(new_net_2894),
		.dout(new_net_2895)
	);

	bfr new_net_2896_bfr_after (
		.din(new_net_2895),
		.dout(new_net_2896)
	);

	bfr new_net_2897_bfr_after (
		.din(new_net_2896),
		.dout(new_net_2897)
	);

	bfr new_net_2898_bfr_after (
		.din(new_net_2897),
		.dout(new_net_2898)
	);

	bfr new_net_2899_bfr_after (
		.din(new_net_2898),
		.dout(new_net_2899)
	);

	bfr new_net_2900_bfr_after (
		.din(new_net_2899),
		.dout(new_net_2900)
	);

	bfr new_net_2901_bfr_after (
		.din(new_net_2900),
		.dout(new_net_2901)
	);

	bfr new_net_2902_bfr_after (
		.din(new_net_2901),
		.dout(new_net_2902)
	);

	bfr new_net_2903_bfr_after (
		.din(new_net_2902),
		.dout(new_net_2903)
	);

	bfr new_net_2904_bfr_after (
		.din(new_net_2903),
		.dout(new_net_2904)
	);

	bfr new_net_2905_bfr_after (
		.din(new_net_2904),
		.dout(new_net_2905)
	);

	bfr new_net_2906_bfr_after (
		.din(new_net_2905),
		.dout(new_net_2906)
	);

	bfr new_net_2907_bfr_after (
		.din(new_net_2906),
		.dout(new_net_2907)
	);

	bfr new_net_2908_bfr_after (
		.din(new_net_2907),
		.dout(new_net_2908)
	);

	bfr new_net_2909_bfr_after (
		.din(new_net_2908),
		.dout(new_net_2909)
	);

	bfr new_net_2910_bfr_after (
		.din(new_net_2909),
		.dout(new_net_2910)
	);

	bfr new_net_2911_bfr_after (
		.din(new_net_2910),
		.dout(new_net_2911)
	);

	bfr new_net_2912_bfr_after (
		.din(new_net_2911),
		.dout(new_net_2912)
	);

	bfr G3521_bfr_after (
		.din(new_net_2912),
		.dout(G3521)
	);

	bfr new_net_2913_bfr_after (
		.din(new_net_1467),
		.dout(new_net_2913)
	);

	bfr new_net_2914_bfr_after (
		.din(new_net_2913),
		.dout(new_net_2914)
	);

	bfr new_net_2915_bfr_after (
		.din(new_net_2914),
		.dout(new_net_2915)
	);

	bfr new_net_2916_bfr_after (
		.din(new_net_2915),
		.dout(new_net_2916)
	);

	bfr new_net_2917_bfr_after (
		.din(new_net_2916),
		.dout(new_net_2917)
	);

	bfr new_net_2918_bfr_after (
		.din(new_net_2917),
		.dout(new_net_2918)
	);

	bfr new_net_2919_bfr_after (
		.din(new_net_2918),
		.dout(new_net_2919)
	);

	bfr new_net_2920_bfr_after (
		.din(new_net_2919),
		.dout(new_net_2920)
	);

	bfr new_net_2921_bfr_after (
		.din(new_net_2920),
		.dout(new_net_2921)
	);

	bfr new_net_2922_bfr_after (
		.din(new_net_2921),
		.dout(new_net_2922)
	);

	bfr new_net_2923_bfr_after (
		.din(new_net_2922),
		.dout(new_net_2923)
	);

	bfr new_net_2924_bfr_after (
		.din(new_net_2923),
		.dout(new_net_2924)
	);

	bfr new_net_2925_bfr_after (
		.din(new_net_2924),
		.dout(new_net_2925)
	);

	bfr new_net_2926_bfr_after (
		.din(new_net_2925),
		.dout(new_net_2926)
	);

	bfr new_net_2927_bfr_after (
		.din(new_net_2926),
		.dout(new_net_2927)
	);

	bfr new_net_2928_bfr_after (
		.din(new_net_2927),
		.dout(new_net_2928)
	);

	bfr new_net_2929_bfr_after (
		.din(new_net_2928),
		.dout(new_net_2929)
	);

	bfr new_net_2930_bfr_after (
		.din(new_net_2929),
		.dout(new_net_2930)
	);

	bfr new_net_2931_bfr_after (
		.din(new_net_2930),
		.dout(new_net_2931)
	);

	bfr new_net_2932_bfr_after (
		.din(new_net_2931),
		.dout(new_net_2932)
	);

	bfr new_net_2933_bfr_after (
		.din(new_net_2932),
		.dout(new_net_2933)
	);

	bfr new_net_2934_bfr_after (
		.din(new_net_2933),
		.dout(new_net_2934)
	);

	bfr new_net_2935_bfr_after (
		.din(new_net_2934),
		.dout(new_net_2935)
	);

	bfr new_net_2936_bfr_after (
		.din(new_net_2935),
		.dout(new_net_2936)
	);

	bfr new_net_2937_bfr_after (
		.din(new_net_2936),
		.dout(new_net_2937)
	);

	bfr new_net_2938_bfr_after (
		.din(new_net_2937),
		.dout(new_net_2938)
	);

	bfr new_net_2939_bfr_after (
		.din(new_net_2938),
		.dout(new_net_2939)
	);

	bfr new_net_2940_bfr_after (
		.din(new_net_2939),
		.dout(new_net_2940)
	);

	bfr new_net_2941_bfr_after (
		.din(new_net_2940),
		.dout(new_net_2941)
	);

	bfr new_net_2942_bfr_after (
		.din(new_net_2941),
		.dout(new_net_2942)
	);

	bfr new_net_2943_bfr_after (
		.din(new_net_2942),
		.dout(new_net_2943)
	);

	bfr new_net_2944_bfr_after (
		.din(new_net_2943),
		.dout(new_net_2944)
	);

	bfr new_net_2945_bfr_after (
		.din(new_net_2944),
		.dout(new_net_2945)
	);

	bfr new_net_2946_bfr_after (
		.din(new_net_2945),
		.dout(new_net_2946)
	);

	bfr new_net_2947_bfr_after (
		.din(new_net_2946),
		.dout(new_net_2947)
	);

	bfr new_net_2948_bfr_after (
		.din(new_net_2947),
		.dout(new_net_2948)
	);

	bfr new_net_2949_bfr_after (
		.din(new_net_2948),
		.dout(new_net_2949)
	);

	bfr new_net_2950_bfr_after (
		.din(new_net_2949),
		.dout(new_net_2950)
	);

	bfr new_net_2951_bfr_after (
		.din(new_net_2950),
		.dout(new_net_2951)
	);

	bfr new_net_2952_bfr_after (
		.din(new_net_2951),
		.dout(new_net_2952)
	);

	bfr new_net_2953_bfr_after (
		.din(new_net_2952),
		.dout(new_net_2953)
	);

	bfr new_net_2954_bfr_after (
		.din(new_net_2953),
		.dout(new_net_2954)
	);

	bfr new_net_2955_bfr_after (
		.din(new_net_2954),
		.dout(new_net_2955)
	);

	bfr new_net_2956_bfr_after (
		.din(new_net_2955),
		.dout(new_net_2956)
	);

	bfr new_net_2957_bfr_after (
		.din(new_net_2956),
		.dout(new_net_2957)
	);

	bfr new_net_2958_bfr_after (
		.din(new_net_2957),
		.dout(new_net_2958)
	);

	bfr new_net_2959_bfr_after (
		.din(new_net_2958),
		.dout(new_net_2959)
	);

	bfr new_net_2960_bfr_after (
		.din(new_net_2959),
		.dout(new_net_2960)
	);

	bfr G3519_bfr_after (
		.din(new_net_2960),
		.dout(G3519)
	);

	bfr new_net_2961_bfr_after (
		.din(new_net_1479),
		.dout(new_net_2961)
	);

	bfr new_net_2962_bfr_after (
		.din(new_net_2961),
		.dout(new_net_2962)
	);

	bfr new_net_2963_bfr_after (
		.din(new_net_2962),
		.dout(new_net_2963)
	);

	bfr new_net_2964_bfr_after (
		.din(new_net_2963),
		.dout(new_net_2964)
	);

	bfr G3537_bfr_after (
		.din(new_net_2964),
		.dout(G3537)
	);

	bfr new_net_1412_bfr_after (
		.din(_0633_),
		.dout(new_net_1412)
	);

	bfr new_net_1386_bfr_after (
		.din(_0531_),
		.dout(new_net_1386)
	);

	bfr new_net_2965_bfr_after (
		.din(_0003_),
		.dout(new_net_2965)
	);

	bfr new_net_1259_bfr_after (
		.din(new_net_2965),
		.dout(new_net_1259)
	);

	bfr new_net_2966_bfr_after (
		.din(_0705_),
		.dout(new_net_2966)
	);

	bfr new_net_1256_bfr_after (
		.din(new_net_2966),
		.dout(new_net_1256)
	);

	bfr new_net_2967_bfr_after (
		.din(_0408_),
		.dout(new_net_2967)
	);

	bfr new_net_1345_bfr_after (
		.din(new_net_2967),
		.dout(new_net_1345)
	);

	bfr new_net_2968_bfr_after (
		.din(_0605_),
		.dout(new_net_2968)
	);

	bfr new_net_2969_bfr_after (
		.din(new_net_2968),
		.dout(new_net_2969)
	);

	bfr new_net_2970_bfr_after (
		.din(new_net_2969),
		.dout(new_net_2970)
	);

	bfr new_net_2971_bfr_after (
		.din(new_net_2970),
		.dout(new_net_2971)
	);

	bfr new_net_2972_bfr_after (
		.din(new_net_2971),
		.dout(new_net_2972)
	);

	bfr new_net_2973_bfr_after (
		.din(new_net_2972),
		.dout(new_net_2973)
	);

	bfr new_net_2974_bfr_after (
		.din(new_net_2973),
		.dout(new_net_2974)
	);

	bfr new_net_2975_bfr_after (
		.din(new_net_2974),
		.dout(new_net_2975)
	);

	bfr new_net_2976_bfr_after (
		.din(new_net_2975),
		.dout(new_net_2976)
	);

	bfr new_net_2977_bfr_after (
		.din(new_net_2976),
		.dout(new_net_2977)
	);

	bfr new_net_1408_bfr_after (
		.din(new_net_2977),
		.dout(new_net_1408)
	);

	bfr new_net_1434_bfr_after (
		.din(_0689_),
		.dout(new_net_1434)
	);

	bfr new_net_2978_bfr_after (
		.din(_0487_),
		.dout(new_net_2978)
	);

	bfr new_net_1372_bfr_after (
		.din(new_net_2978),
		.dout(new_net_1372)
	);

	bfr new_net_2979_bfr_after (
		.din(_0757_),
		.dout(new_net_2979)
	);

	bfr new_net_2980_bfr_after (
		.din(new_net_2979),
		.dout(new_net_2980)
	);

	bfr new_net_2981_bfr_after (
		.din(new_net_2980),
		.dout(new_net_2981)
	);

	bfr new_net_2982_bfr_after (
		.din(new_net_2981),
		.dout(new_net_2982)
	);

	bfr new_net_2983_bfr_after (
		.din(new_net_2982),
		.dout(new_net_2983)
	);

	bfr new_net_2984_bfr_after (
		.din(new_net_2983),
		.dout(new_net_2984)
	);

	bfr new_net_2985_bfr_after (
		.din(new_net_2984),
		.dout(new_net_2985)
	);

	bfr new_net_2986_bfr_after (
		.din(new_net_2985),
		.dout(new_net_2986)
	);

	bfr new_net_2987_bfr_after (
		.din(new_net_2986),
		.dout(new_net_2987)
	);

	bfr new_net_2988_bfr_after (
		.din(new_net_2987),
		.dout(new_net_2988)
	);

	bfr new_net_2989_bfr_after (
		.din(new_net_2988),
		.dout(new_net_2989)
	);

	bfr new_net_2990_bfr_after (
		.din(new_net_2989),
		.dout(new_net_2990)
	);

	bfr new_net_2991_bfr_after (
		.din(new_net_2990),
		.dout(new_net_2991)
	);

	bfr new_net_2992_bfr_after (
		.din(new_net_2991),
		.dout(new_net_2992)
	);

	bfr new_net_2993_bfr_after (
		.din(new_net_2992),
		.dout(new_net_2993)
	);

	bfr new_net_2994_bfr_after (
		.din(new_net_2993),
		.dout(new_net_2994)
	);

	bfr new_net_2995_bfr_after (
		.din(new_net_2994),
		.dout(new_net_2995)
	);

	bfr new_net_2996_bfr_after (
		.din(new_net_2995),
		.dout(new_net_2996)
	);

	bfr new_net_1456_bfr_after (
		.din(new_net_2996),
		.dout(new_net_1456)
	);

	bfr new_net_1430_bfr_after (
		.din(_0671_),
		.dout(new_net_1430)
	);

	bfr new_net_2997_bfr_after (
		.din(_0737_),
		.dout(new_net_2997)
	);

	bfr new_net_1451_bfr_after (
		.din(new_net_2997),
		.dout(new_net_1451)
	);

	bfr new_net_1281_bfr_after (
		.din(_0121_),
		.dout(new_net_1281)
	);

	bfr new_net_2998_bfr_after (
		.din(_0198_),
		.dout(new_net_2998)
	);

	bfr new_net_1302_bfr_after (
		.din(new_net_2998),
		.dout(new_net_1302)
	);

	bfr new_net_1323_bfr_after (
		.din(_0276_),
		.dout(new_net_1323)
	);

	bfr new_net_2999_bfr_after (
		.din(_0090_),
		.dout(new_net_2999)
	);

	bfr new_net_1273_bfr_after (
		.din(new_net_2999),
		.dout(new_net_1273)
	);

	bfr new_net_1277_bfr_after (
		.din(_0105_),
		.dout(new_net_1277)
	);

	bfr new_net_1294_bfr_after (
		.din(_0171_),
		.dout(new_net_1294)
	);

	bfr new_net_3000_bfr_after (
		.din(_0240_),
		.dout(new_net_3000)
	);

	bfr new_net_1315_bfr_after (
		.din(new_net_3000),
		.dout(new_net_1315)
	);

	bfr new_net_1298_bfr_after (
		.din(_0176_),
		.dout(new_net_1298)
	);

	bfr new_net_3001_bfr_after (
		.din(_0259_),
		.dout(new_net_3001)
	);

	bfr new_net_3002_bfr_after (
		.din(new_net_3001),
		.dout(new_net_3002)
	);

	bfr new_net_1319_bfr_after (
		.din(new_net_3002),
		.dout(new_net_1319)
	);

	bfr new_net_1336_bfr_after (
		.din(_0358_),
		.dout(new_net_1336)
	);

	bfr new_net_3003_bfr_after (
		.din(_0567_),
		.dout(new_net_3003)
	);

	bfr new_net_3004_bfr_after (
		.din(new_net_3003),
		.dout(new_net_3004)
	);

	bfr new_net_3005_bfr_after (
		.din(new_net_3004),
		.dout(new_net_3005)
	);

	bfr new_net_1394_bfr_after (
		.din(new_net_3005),
		.dout(new_net_1394)
	);

	bfr new_net_3006_bfr_after (
		.din(_0585_),
		.dout(new_net_3006)
	);

	bfr new_net_1399_bfr_after (
		.din(new_net_3006),
		.dout(new_net_1399)
	);

	bfr new_net_3007_bfr_after (
		.din(new_net_1485),
		.dout(new_net_3007)
	);

	bfr new_net_3008_bfr_after (
		.din(new_net_3007),
		.dout(new_net_3008)
	);

	bfr new_net_3009_bfr_after (
		.din(new_net_3008),
		.dout(new_net_3009)
	);

	bfr new_net_3010_bfr_after (
		.din(new_net_3009),
		.dout(new_net_3010)
	);

	bfr new_net_3011_bfr_after (
		.din(new_net_3010),
		.dout(new_net_3011)
	);

	bfr new_net_3012_bfr_after (
		.din(new_net_3011),
		.dout(new_net_3012)
	);

	bfr new_net_3013_bfr_after (
		.din(new_net_3012),
		.dout(new_net_3013)
	);

	bfr new_net_3014_bfr_after (
		.din(new_net_3013),
		.dout(new_net_3014)
	);

	bfr new_net_3015_bfr_after (
		.din(new_net_3014),
		.dout(new_net_3015)
	);

	bfr new_net_3016_bfr_after (
		.din(new_net_3015),
		.dout(new_net_3016)
	);

	bfr new_net_3017_bfr_after (
		.din(new_net_3016),
		.dout(new_net_3017)
	);

	bfr new_net_3018_bfr_after (
		.din(new_net_3017),
		.dout(new_net_3018)
	);

	bfr new_net_3019_bfr_after (
		.din(new_net_3018),
		.dout(new_net_3019)
	);

	bfr new_net_3020_bfr_after (
		.din(new_net_3019),
		.dout(new_net_3020)
	);

	bfr new_net_3021_bfr_after (
		.din(new_net_3020),
		.dout(new_net_3021)
	);

	bfr new_net_3022_bfr_after (
		.din(new_net_3021),
		.dout(new_net_3022)
	);

	bfr new_net_3023_bfr_after (
		.din(new_net_3022),
		.dout(new_net_3023)
	);

	bfr G3530_bfr_after (
		.din(new_net_3023),
		.dout(G3530)
	);

	bfr new_net_3024_bfr_after (
		.din(_0647_),
		.dout(new_net_3024)
	);

	bfr new_net_3025_bfr_after (
		.din(new_net_3024),
		.dout(new_net_3025)
	);

	bfr new_net_3026_bfr_after (
		.din(new_net_3025),
		.dout(new_net_3026)
	);

	bfr new_net_1421_bfr_after (
		.din(new_net_3026),
		.dout(new_net_1421)
	);

	bfr new_net_3027_bfr_after (
		.din(_0709_),
		.dout(new_net_3027)
	);

	bfr new_net_1442_bfr_after (
		.din(new_net_3027),
		.dout(new_net_1442)
	);

	bfr new_net_3028_bfr_after (
		.din(_0639_),
		.dout(new_net_3028)
	);

	bfr new_net_1416_bfr_after (
		.din(new_net_3028),
		.dout(new_net_1416)
	);

	bfr new_net_3029_bfr_after (
		.din(_0452_),
		.dout(new_net_3029)
	);

	bfr new_net_1359_bfr_after (
		.din(new_net_3029),
		.dout(new_net_1359)
	);

	bfr new_net_3030_bfr_after (
		.din(_0694_),
		.dout(new_net_3030)
	);

	bfr new_net_3031_bfr_after (
		.din(new_net_3030),
		.dout(new_net_3031)
	);

	bfr new_net_1438_bfr_after (
		.din(new_net_3031),
		.dout(new_net_1438)
	);

	bfr new_net_3032_bfr_after (
		.din(_0519_),
		.dout(new_net_3032)
	);

	bfr new_net_1381_bfr_after (
		.din(new_net_3032),
		.dout(new_net_1381)
	);

	bfr new_net_1376_bfr_after (
		.din(_0502_),
		.dout(new_net_1376)
	);

	bfr new_net_1460_bfr_after (
		.din(_0779_),
		.dout(new_net_1460)
	);

	bfr new_net_3033_bfr_after (
		.din(_0730_),
		.dout(new_net_3033)
	);

	bfr new_net_3034_bfr_after (
		.din(new_net_3033),
		.dout(new_net_3034)
	);

	bfr new_net_3035_bfr_after (
		.din(new_net_3034),
		.dout(new_net_3035)
	);

	bfr new_net_3036_bfr_after (
		.din(new_net_3035),
		.dout(new_net_3036)
	);

	bfr new_net_3037_bfr_after (
		.din(new_net_3036),
		.dout(new_net_3037)
	);

	bfr new_net_1448_bfr_after (
		.din(new_net_3037),
		.dout(new_net_1448)
	);

	bfr new_net_3038_bfr_after (
		.din(_0387_),
		.dout(new_net_3038)
	);

	bfr new_net_1340_bfr_after (
		.din(new_net_3038),
		.dout(new_net_1340)
	);

	bfr new_net_3039_bfr_after (
		.din(_0594_),
		.dout(new_net_3039)
	);

	bfr new_net_3040_bfr_after (
		.din(new_net_3039),
		.dout(new_net_3040)
	);

	bfr new_net_1403_bfr_after (
		.din(new_net_3040),
		.dout(new_net_1403)
	);

	bfr new_net_1398_bfr_after (
		.din(_0577_),
		.dout(new_net_1398)
	);

	bfr new_net_1453_bfr_after (
		.din(_0741_),
		.dout(new_net_1453)
	);

	bfr new_net_1289_bfr_after (
		.din(_0149_),
		.dout(new_net_1289)
	);

	bfr new_net_1310_bfr_after (
		.din(_0215_),
		.dout(new_net_1310)
	);

	bfr new_net_1331_bfr_after (
		.din(_0320_),
		.dout(new_net_1331)
	);

	bfr new_net_3041_bfr_after (
		.din(_0210_),
		.dout(new_net_3041)
	);

	bfr new_net_1306_bfr_after (
		.din(new_net_3041),
		.dout(new_net_1306)
	);

	bfr new_net_1272_bfr_after (
		.din(_0081_),
		.dout(new_net_1272)
	);

	bfr new_net_1293_bfr_after (
		.din(_0166_),
		.dout(new_net_1293)
	);

	bfr new_net_3042_bfr_after (
		.din(_0234_),
		.dout(new_net_3042)
	);

	bfr new_net_3043_bfr_after (
		.din(new_net_3042),
		.dout(new_net_3043)
	);

	bfr new_net_3044_bfr_after (
		.din(new_net_3043),
		.dout(new_net_3044)
	);

	bfr new_net_1314_bfr_after (
		.din(new_net_3044),
		.dout(new_net_1314)
	);

	bfr new_net_1327_bfr_after (
		.din(_0291_),
		.dout(new_net_1327)
	);

	bfr new_net_1255_bfr_after (
		.din(_0673_),
		.dout(new_net_1255)
	);

	bfr new_net_1258_bfr_after (
		.din(_0002_),
		.dout(new_net_1258)
	);

	bfr new_net_3045_bfr_after (
		.din(_0667_),
		.dout(new_net_3045)
	);

	bfr new_net_3046_bfr_after (
		.din(new_net_3045),
		.dout(new_net_3046)
	);

	bfr new_net_3047_bfr_after (
		.din(new_net_3046),
		.dout(new_net_3047)
	);

	bfr new_net_1425_bfr_after (
		.din(new_net_3047),
		.dout(new_net_1425)
	);

	bfr new_net_1446_bfr_after (
		.din(_0714_),
		.dout(new_net_1446)
	);

	bfr new_net_3048_bfr_after (
		.din(_0538_),
		.dout(new_net_3048)
	);

	bfr new_net_3049_bfr_after (
		.din(new_net_3048),
		.dout(new_net_3049)
	);

	bfr new_net_3050_bfr_after (
		.din(new_net_3049),
		.dout(new_net_3050)
	);

	bfr new_net_3051_bfr_after (
		.din(new_net_3050),
		.dout(new_net_3051)
	);

	bfr new_net_3052_bfr_after (
		.din(new_net_3051),
		.dout(new_net_3052)
	);

	bfr new_net_3053_bfr_after (
		.din(new_net_3052),
		.dout(new_net_3053)
	);

	bfr new_net_3054_bfr_after (
		.din(new_net_3053),
		.dout(new_net_3054)
	);

	bfr new_net_3055_bfr_after (
		.din(new_net_3054),
		.dout(new_net_3055)
	);

	bfr new_net_3056_bfr_after (
		.din(new_net_3055),
		.dout(new_net_3056)
	);

	bfr new_net_3057_bfr_after (
		.din(new_net_3056),
		.dout(new_net_3057)
	);

	bfr new_net_3058_bfr_after (
		.din(new_net_3057),
		.dout(new_net_3058)
	);

	bfr new_net_3059_bfr_after (
		.din(new_net_3058),
		.dout(new_net_3059)
	);

	bfr new_net_3060_bfr_after (
		.din(new_net_3059),
		.dout(new_net_3060)
	);

	bfr new_net_3061_bfr_after (
		.din(new_net_3060),
		.dout(new_net_3061)
	);

	bfr new_net_1389_bfr_after (
		.din(new_net_3061),
		.dout(new_net_1389)
	);

	bfr new_net_3062_bfr_after (
		.din(_0467_),
		.dout(new_net_3062)
	);

	bfr new_net_3063_bfr_after (
		.din(new_net_3062),
		.dout(new_net_3063)
	);

	bfr new_net_1363_bfr_after (
		.din(new_net_3063),
		.dout(new_net_1363)
	);

	bfr new_net_3064_bfr_after (
		.din(_0628_),
		.dout(new_net_3064)
	);

	bfr new_net_1411_bfr_after (
		.din(new_net_3064),
		.dout(new_net_1411)
	);

	bfr new_net_3065_bfr_after (
		.din(_0529_),
		.dout(new_net_3065)
	);

	bfr new_net_1385_bfr_after (
		.din(new_net_3065),
		.dout(new_net_1385)
	);

	bfr new_net_1433_bfr_after (
		.din(_0687_),
		.dout(new_net_1433)
	);

	bfr new_net_3066_bfr_after (
		.din(_0393_),
		.dout(new_net_3066)
	);

	bfr new_net_3067_bfr_after (
		.din(new_net_3066),
		.dout(new_net_3067)
	);

	bfr new_net_1344_bfr_after (
		.din(new_net_3067),
		.dout(new_net_1344)
	);

	bfr new_net_1407_bfr_after (
		.din(_0607_),
		.dout(new_net_1407)
	);

	bfr new_net_3068_bfr_after (
		.din(_0491_),
		.dout(new_net_3068)
	);

	bfr new_net_1371_bfr_after (
		.din(new_net_3068),
		.dout(new_net_1371)
	);

	bfr new_net_1455_bfr_after (
		.din(_0745_),
		.dout(new_net_1455)
	);

	bfr new_net_3069_bfr_after (
		.din(_0675_),
		.dout(new_net_3069)
	);

	bfr new_net_3070_bfr_after (
		.din(new_net_3069),
		.dout(new_net_3070)
	);

	bfr new_net_3071_bfr_after (
		.din(new_net_3070),
		.dout(new_net_3071)
	);

	bfr new_net_3072_bfr_after (
		.din(new_net_3071),
		.dout(new_net_3072)
	);

	bfr new_net_3073_bfr_after (
		.din(new_net_3072),
		.dout(new_net_3073)
	);

	bfr new_net_3074_bfr_after (
		.din(new_net_3073),
		.dout(new_net_3074)
	);

	bfr new_net_3075_bfr_after (
		.din(new_net_3074),
		.dout(new_net_3075)
	);

	bfr new_net_1429_bfr_after (
		.din(new_net_3075),
		.dout(new_net_1429)
	);

	bfr new_net_3076_bfr_after (
		.din(_0733_),
		.dout(new_net_3076)
	);

	bfr new_net_3077_bfr_after (
		.din(new_net_3076),
		.dout(new_net_3077)
	);

	bfr new_net_3078_bfr_after (
		.din(new_net_3077),
		.dout(new_net_3078)
	);

	bfr new_net_1450_bfr_after (
		.din(new_net_3078),
		.dout(new_net_1450)
	);

	bfr new_net_1393_bfr_after (
		.din(_0562_),
		.dout(new_net_1393)
	);

	bfr new_net_1367_bfr_after (
		.din(_0477_),
		.dout(new_net_1367)
	);

	bfr new_net_1276_bfr_after (
		.din(_0104_),
		.dout(new_net_1276)
	);

	bfr new_net_1280_bfr_after (
		.din(_0111_),
		.dout(new_net_1280)
	);

	bfr new_net_3079_bfr_after (
		.din(_0181_),
		.dout(new_net_3079)
	);

	bfr new_net_3080_bfr_after (
		.din(new_net_3079),
		.dout(new_net_3080)
	);

	bfr new_net_1297_bfr_after (
		.din(new_net_3080),
		.dout(new_net_1297)
	);

	bfr new_net_1318_bfr_after (
		.din(_0256_),
		.dout(new_net_1318)
	);

	bfr new_net_3081_bfr_after (
		.din(_0275_),
		.dout(new_net_3081)
	);

	bfr new_net_3082_bfr_after (
		.din(new_net_3081),
		.dout(new_net_3082)
	);

	bfr new_net_1322_bfr_after (
		.din(new_net_3082),
		.dout(new_net_1322)
	);

	bfr new_net_3083_bfr_after (
		.din(_0196_),
		.dout(new_net_3083)
	);

	bfr new_net_1301_bfr_after (
		.din(new_net_3083),
		.dout(new_net_1301)
	);

	bfr new_net_1339_bfr_after (
		.din(_0381_),
		.dout(new_net_1339)
	);

	bfr new_net_3084_bfr_after (
		.din(_0400_),
		.dout(new_net_3084)
	);

	bfr new_net_3085_bfr_after (
		.din(new_net_3084),
		.dout(new_net_3085)
	);

	bfr new_net_1343_bfr_after (
		.din(new_net_3085),
		.dout(new_net_1343)
	);

	bfr new_net_3086_bfr_after (
		.din(_0455_),
		.dout(new_net_3086)
	);

	bfr new_net_3087_bfr_after (
		.din(new_net_3086),
		.dout(new_net_3087)
	);

	bfr new_net_3088_bfr_after (
		.din(new_net_3087),
		.dout(new_net_3088)
	);

	bfr new_net_3089_bfr_after (
		.din(new_net_3088),
		.dout(new_net_3089)
	);

	bfr new_net_3090_bfr_after (
		.din(new_net_3089),
		.dout(new_net_3090)
	);

	bfr new_net_3091_bfr_after (
		.din(new_net_3090),
		.dout(new_net_3091)
	);

	bfr new_net_3092_bfr_after (
		.din(new_net_3091),
		.dout(new_net_3092)
	);

	bfr new_net_3093_bfr_after (
		.din(new_net_3092),
		.dout(new_net_3093)
	);

	bfr new_net_1360_bfr_after (
		.din(new_net_3093),
		.dout(new_net_1360)
	);

	bfr new_net_3094_bfr_after (
		.din(_0466_),
		.dout(new_net_3094)
	);

	bfr new_net_1364_bfr_after (
		.din(new_net_3094),
		.dout(new_net_1364)
	);

	bfr new_net_3095_bfr_after (
		.din(_0638_),
		.dout(new_net_3095)
	);

	bfr new_net_3096_bfr_after (
		.din(new_net_3095),
		.dout(new_net_3096)
	);

	bfr new_net_1415_bfr_after (
		.din(new_net_3096),
		.dout(new_net_1415)
	);

	bfr new_net_3097_bfr_after (
		.din(_0650_),
		.dout(new_net_3097)
	);

	bfr new_net_3098_bfr_after (
		.din(new_net_3097),
		.dout(new_net_3098)
	);

	bfr new_net_1420_bfr_after (
		.din(new_net_3098),
		.dout(new_net_1420)
	);

	bfr new_net_3099_bfr_after (
		.din(_0712_),
		.dout(new_net_3099)
	);

	bfr new_net_3100_bfr_after (
		.din(new_net_3099),
		.dout(new_net_3100)
	);

	bfr new_net_1441_bfr_after (
		.din(new_net_3100),
		.dout(new_net_1441)
	);

	bfr new_net_3101_bfr_after (
		.din(_0448_),
		.dout(new_net_3101)
	);

	bfr new_net_1358_bfr_after (
		.din(new_net_3101),
		.dout(new_net_1358)
	);

	bfr new_net_3102_bfr_after (
		.din(_0427_),
		.dout(new_net_3102)
	);

	bfr new_net_1353_bfr_after (
		.din(new_net_3102),
		.dout(new_net_1353)
	);

	bfr new_net_3103_bfr_after (
		.din(_0697_),
		.dout(new_net_3103)
	);

	bfr new_net_1437_bfr_after (
		.din(new_net_3103),
		.dout(new_net_1437)
	);

	bfr new_net_1380_bfr_after (
		.din(_0514_),
		.dout(new_net_1380)
	);

	bfr new_net_1375_bfr_after (
		.din(_0500_),
		.dout(new_net_1375)
	);

	bfr new_net_3104_bfr_after (
		.din(_0773_),
		.dout(new_net_3104)
	);

	bfr new_net_3105_bfr_after (
		.din(new_net_3104),
		.dout(new_net_3105)
	);

	bfr new_net_1459_bfr_after (
		.din(new_net_3105),
		.dout(new_net_1459)
	);

	bfr new_net_3106_bfr_after (
		.din(new_net_1463),
		.dout(new_net_3106)
	);

	bfr new_net_3107_bfr_after (
		.din(new_net_3106),
		.dout(new_net_3107)
	);

	bfr new_net_3108_bfr_after (
		.din(new_net_3107),
		.dout(new_net_3108)
	);

	bfr new_net_3109_bfr_after (
		.din(new_net_3108),
		.dout(new_net_3109)
	);

	bfr new_net_3110_bfr_after (
		.din(new_net_3109),
		.dout(new_net_3110)
	);

	bfr new_net_3111_bfr_after (
		.din(new_net_3110),
		.dout(new_net_3111)
	);

	bfr new_net_3112_bfr_after (
		.din(new_net_3111),
		.dout(new_net_3112)
	);

	bfr new_net_3113_bfr_after (
		.din(new_net_3112),
		.dout(new_net_3113)
	);

	bfr new_net_3114_bfr_after (
		.din(new_net_3113),
		.dout(new_net_3114)
	);

	bfr new_net_3115_bfr_after (
		.din(new_net_3114),
		.dout(new_net_3115)
	);

	bfr new_net_3116_bfr_after (
		.din(new_net_3115),
		.dout(new_net_3116)
	);

	bfr new_net_3117_bfr_after (
		.din(new_net_3116),
		.dout(new_net_3117)
	);

	bfr new_net_3118_bfr_after (
		.din(new_net_3117),
		.dout(new_net_3118)
	);

	bfr new_net_3119_bfr_after (
		.din(new_net_3118),
		.dout(new_net_3119)
	);

	bfr new_net_3120_bfr_after (
		.din(new_net_3119),
		.dout(new_net_3120)
	);

	bfr new_net_3121_bfr_after (
		.din(new_net_3120),
		.dout(new_net_3121)
	);

	bfr new_net_3122_bfr_after (
		.din(new_net_3121),
		.dout(new_net_3122)
	);

	bfr new_net_3123_bfr_after (
		.din(new_net_3122),
		.dout(new_net_3123)
	);

	bfr new_net_3124_bfr_after (
		.din(new_net_3123),
		.dout(new_net_3124)
	);

	bfr new_net_3125_bfr_after (
		.din(new_net_3124),
		.dout(new_net_3125)
	);

	bfr new_net_3126_bfr_after (
		.din(new_net_3125),
		.dout(new_net_3126)
	);

	bfr new_net_3127_bfr_after (
		.din(new_net_3126),
		.dout(new_net_3127)
	);

	bfr new_net_3128_bfr_after (
		.din(new_net_3127),
		.dout(new_net_3128)
	);

	bfr new_net_3129_bfr_after (
		.din(new_net_3128),
		.dout(new_net_3129)
	);

	bfr new_net_3130_bfr_after (
		.din(new_net_3129),
		.dout(new_net_3130)
	);

	bfr new_net_3131_bfr_after (
		.din(new_net_3130),
		.dout(new_net_3131)
	);

	bfr new_net_3132_bfr_after (
		.din(new_net_3131),
		.dout(new_net_3132)
	);

	bfr new_net_3133_bfr_after (
		.din(new_net_3132),
		.dout(new_net_3133)
	);

	bfr new_net_3134_bfr_after (
		.din(new_net_3133),
		.dout(new_net_3134)
	);

	bfr new_net_3135_bfr_after (
		.din(new_net_3134),
		.dout(new_net_3135)
	);

	bfr new_net_3136_bfr_after (
		.din(new_net_3135),
		.dout(new_net_3136)
	);

	bfr new_net_3137_bfr_after (
		.din(new_net_3136),
		.dout(new_net_3137)
	);

	bfr new_net_3138_bfr_after (
		.din(new_net_3137),
		.dout(new_net_3138)
	);

	bfr new_net_3139_bfr_after (
		.din(new_net_3138),
		.dout(new_net_3139)
	);

	bfr new_net_3140_bfr_after (
		.din(new_net_3139),
		.dout(new_net_3140)
	);

	bfr new_net_3141_bfr_after (
		.din(new_net_3140),
		.dout(new_net_3141)
	);

	bfr new_net_3142_bfr_after (
		.din(new_net_3141),
		.dout(new_net_3142)
	);

	bfr new_net_3143_bfr_after (
		.din(new_net_3142),
		.dout(new_net_3143)
	);

	bfr new_net_3144_bfr_after (
		.din(new_net_3143),
		.dout(new_net_3144)
	);

	bfr new_net_3145_bfr_after (
		.din(new_net_3144),
		.dout(new_net_3145)
	);

	bfr new_net_3146_bfr_after (
		.din(new_net_3145),
		.dout(new_net_3146)
	);

	bfr new_net_3147_bfr_after (
		.din(new_net_3146),
		.dout(new_net_3147)
	);

	bfr G3523_bfr_after (
		.din(new_net_3147),
		.dout(G3523)
	);

	bfr new_net_3148_bfr_after (
		.din(new_net_1475),
		.dout(new_net_3148)
	);

	bfr new_net_3149_bfr_after (
		.din(new_net_3148),
		.dout(new_net_3149)
	);

	bfr new_net_3150_bfr_after (
		.din(new_net_3149),
		.dout(new_net_3150)
	);

	bfr new_net_3151_bfr_after (
		.din(new_net_3150),
		.dout(new_net_3151)
	);

	bfr new_net_3152_bfr_after (
		.din(new_net_3151),
		.dout(new_net_3152)
	);

	bfr new_net_3153_bfr_after (
		.din(new_net_3152),
		.dout(new_net_3153)
	);

	bfr new_net_3154_bfr_after (
		.din(new_net_3153),
		.dout(new_net_3154)
	);

	bfr new_net_3155_bfr_after (
		.din(new_net_3154),
		.dout(new_net_3155)
	);

	bfr new_net_3156_bfr_after (
		.din(new_net_3155),
		.dout(new_net_3156)
	);

	bfr new_net_3157_bfr_after (
		.din(new_net_3156),
		.dout(new_net_3157)
	);

	bfr new_net_3158_bfr_after (
		.din(new_net_3157),
		.dout(new_net_3158)
	);

	bfr new_net_3159_bfr_after (
		.din(new_net_3158),
		.dout(new_net_3159)
	);

	bfr new_net_3160_bfr_after (
		.din(new_net_3159),
		.dout(new_net_3160)
	);

	bfr new_net_3161_bfr_after (
		.din(new_net_3160),
		.dout(new_net_3161)
	);

	bfr new_net_3162_bfr_after (
		.din(new_net_3161),
		.dout(new_net_3162)
	);

	bfr new_net_3163_bfr_after (
		.din(new_net_3162),
		.dout(new_net_3163)
	);

	bfr new_net_3164_bfr_after (
		.din(new_net_3163),
		.dout(new_net_3164)
	);

	bfr new_net_3165_bfr_after (
		.din(new_net_3164),
		.dout(new_net_3165)
	);

	bfr new_net_3166_bfr_after (
		.din(new_net_3165),
		.dout(new_net_3166)
	);

	bfr new_net_3167_bfr_after (
		.din(new_net_3166),
		.dout(new_net_3167)
	);

	bfr new_net_3168_bfr_after (
		.din(new_net_3167),
		.dout(new_net_3168)
	);

	bfr new_net_3169_bfr_after (
		.din(new_net_3168),
		.dout(new_net_3169)
	);

	bfr new_net_3170_bfr_after (
		.din(new_net_3169),
		.dout(new_net_3170)
	);

	bfr new_net_3171_bfr_after (
		.din(new_net_3170),
		.dout(new_net_3171)
	);

	bfr new_net_3172_bfr_after (
		.din(new_net_3171),
		.dout(new_net_3172)
	);

	bfr new_net_3173_bfr_after (
		.din(new_net_3172),
		.dout(new_net_3173)
	);

	bfr new_net_3174_bfr_after (
		.din(new_net_3173),
		.dout(new_net_3174)
	);

	bfr new_net_3175_bfr_after (
		.din(new_net_3174),
		.dout(new_net_3175)
	);

	bfr new_net_3176_bfr_after (
		.din(new_net_3175),
		.dout(new_net_3176)
	);

	bfr new_net_3177_bfr_after (
		.din(new_net_3176),
		.dout(new_net_3177)
	);

	bfr new_net_3178_bfr_after (
		.din(new_net_3177),
		.dout(new_net_3178)
	);

	bfr new_net_3179_bfr_after (
		.din(new_net_3178),
		.dout(new_net_3179)
	);

	bfr new_net_3180_bfr_after (
		.din(new_net_3179),
		.dout(new_net_3180)
	);

	bfr new_net_3181_bfr_after (
		.din(new_net_3180),
		.dout(new_net_3181)
	);

	bfr new_net_3182_bfr_after (
		.din(new_net_3181),
		.dout(new_net_3182)
	);

	bfr new_net_3183_bfr_after (
		.din(new_net_3182),
		.dout(new_net_3183)
	);

	bfr new_net_3184_bfr_after (
		.din(new_net_3183),
		.dout(new_net_3184)
	);

	bfr new_net_3185_bfr_after (
		.din(new_net_3184),
		.dout(new_net_3185)
	);

	bfr new_net_3186_bfr_after (
		.din(new_net_3185),
		.dout(new_net_3186)
	);

	bfr new_net_3187_bfr_after (
		.din(new_net_3186),
		.dout(new_net_3187)
	);

	bfr new_net_3188_bfr_after (
		.din(new_net_3187),
		.dout(new_net_3188)
	);

	bfr new_net_3189_bfr_after (
		.din(new_net_3188),
		.dout(new_net_3189)
	);

	bfr new_net_3190_bfr_after (
		.din(new_net_3189),
		.dout(new_net_3190)
	);

	bfr new_net_3191_bfr_after (
		.din(new_net_3190),
		.dout(new_net_3191)
	);

	bfr new_net_3192_bfr_after (
		.din(new_net_3191),
		.dout(new_net_3192)
	);

	bfr new_net_3193_bfr_after (
		.din(new_net_3192),
		.dout(new_net_3193)
	);

	bfr new_net_3194_bfr_after (
		.din(new_net_3193),
		.dout(new_net_3194)
	);

	bfr new_net_3195_bfr_after (
		.din(new_net_3194),
		.dout(new_net_3195)
	);

	bfr G3520_bfr_after (
		.din(new_net_3195),
		.dout(G3520)
	);

	bfr new_net_1402_bfr_after (
		.din(_0589_),
		.dout(new_net_1402)
	);

	bfr new_net_1397_bfr_after (
		.din(_0580_),
		.dout(new_net_1397)
	);

	bfr new_net_1424_bfr_after (
		.din(_0666_),
		.dout(new_net_1424)
	);

	bfr new_net_3196_bfr_after (
		.din(_0721_),
		.dout(new_net_3196)
	);

	bfr new_net_3197_bfr_after (
		.din(new_net_3196),
		.dout(new_net_3197)
	);

	bfr new_net_1445_bfr_after (
		.din(new_net_3197),
		.dout(new_net_1445)
	);

	bfr new_net_3198_bfr_after (
		.din(_0335_),
		.dout(new_net_3198)
	);

	bfr new_net_3199_bfr_after (
		.din(new_net_3198),
		.dout(new_net_3199)
	);

	bfr new_net_3200_bfr_after (
		.din(new_net_3199),
		.dout(new_net_3200)
	);

	bfr new_net_3201_bfr_after (
		.din(new_net_3200),
		.dout(new_net_3201)
	);

	bfr new_net_1335_bfr_after (
		.din(new_net_3201),
		.dout(new_net_1335)
	);

	bfr new_net_3202_bfr_after (
		.din(_0654_),
		.dout(new_net_3202)
	);

	bfr new_net_3203_bfr_after (
		.din(new_net_3202),
		.dout(new_net_3203)
	);

	bfr new_net_3204_bfr_after (
		.din(new_net_3203),
		.dout(new_net_3204)
	);

	bfr new_net_3205_bfr_after (
		.din(new_net_3204),
		.dout(new_net_3205)
	);

	bfr new_net_1419_bfr_after (
		.din(new_net_3205),
		.dout(new_net_1419)
	);

	bfr new_net_3206_bfr_after (
		.din(_0297_),
		.dout(new_net_3206)
	);

	bfr new_net_3207_bfr_after (
		.din(new_net_3206),
		.dout(new_net_3207)
	);

	bfr new_net_3208_bfr_after (
		.din(new_net_3207),
		.dout(new_net_3208)
	);

	bfr new_net_3209_bfr_after (
		.din(new_net_3208),
		.dout(new_net_3209)
	);

	bfr new_net_3210_bfr_after (
		.din(new_net_3209),
		.dout(new_net_3210)
	);

	bfr new_net_3211_bfr_after (
		.din(new_net_3210),
		.dout(new_net_3211)
	);

	bfr new_net_3212_bfr_after (
		.din(new_net_3211),
		.dout(new_net_3212)
	);

	bfr new_net_1330_bfr_after (
		.din(new_net_3212),
		.dout(new_net_1330)
	);

	bfr new_net_1288_bfr_after (
		.din(_0144_),
		.dout(new_net_1288)
	);

	bfr new_net_1309_bfr_after (
		.din(_0219_),
		.dout(new_net_1309)
	);

	bfr new_net_1292_bfr_after (
		.din(_0159_),
		.dout(new_net_1292)
	);

	bfr new_net_1313_bfr_after (
		.din(_0232_),
		.dout(new_net_1313)
	);

	bfr new_net_1263_bfr_after (
		.din(_0029_),
		.dout(new_net_1263)
	);

	bfr new_net_1267_bfr_after (
		.din(_0067_),
		.dout(new_net_1267)
	);

	bfr new_net_1271_bfr_after (
		.din(_0073_),
		.dout(new_net_1271)
	);

	bfr new_net_1284_bfr_after (
		.din(_0127_),
		.dout(new_net_1284)
	);

	bfr new_net_1305_bfr_after (
		.din(_0208_),
		.dout(new_net_1305)
	);

	bfr new_net_3213_bfr_after (
		.din(_0449_),
		.dout(new_net_3213)
	);

	bfr new_net_3214_bfr_after (
		.din(new_net_3213),
		.dout(new_net_3214)
	);

	bfr new_net_3215_bfr_after (
		.din(new_net_3214),
		.dout(new_net_3215)
	);

	bfr new_net_3216_bfr_after (
		.din(new_net_3215),
		.dout(new_net_3216)
	);

	bfr new_net_3217_bfr_after (
		.din(new_net_3216),
		.dout(new_net_3217)
	);

	bfr new_net_3218_bfr_after (
		.din(new_net_3217),
		.dout(new_net_3218)
	);

	bfr new_net_3219_bfr_after (
		.din(new_net_3218),
		.dout(new_net_3219)
	);

	bfr new_net_3220_bfr_after (
		.din(new_net_3219),
		.dout(new_net_3220)
	);

	bfr new_net_3221_bfr_after (
		.din(new_net_3220),
		.dout(new_net_3221)
	);

	bfr new_net_3222_bfr_after (
		.din(new_net_3221),
		.dout(new_net_3222)
	);

	bfr new_net_3223_bfr_after (
		.din(new_net_3222),
		.dout(new_net_3223)
	);

	bfr new_net_3224_bfr_after (
		.din(new_net_3223),
		.dout(new_net_3224)
	);

	bfr new_net_3225_bfr_after (
		.din(new_net_3224),
		.dout(new_net_3225)
	);

	bfr new_net_3226_bfr_after (
		.din(new_net_3225),
		.dout(new_net_3226)
	);

	bfr new_net_3227_bfr_after (
		.din(new_net_3226),
		.dout(new_net_3227)
	);

	bfr new_net_3228_bfr_after (
		.din(new_net_3227),
		.dout(new_net_3228)
	);

	bfr new_net_3229_bfr_after (
		.din(new_net_3228),
		.dout(new_net_3229)
	);

	bfr new_net_3230_bfr_after (
		.din(new_net_3229),
		.dout(new_net_3230)
	);

	bfr new_net_1362_bfr_after (
		.din(new_net_3230),
		.dout(new_net_1362)
	);

	bfr new_net_1326_bfr_after (
		.din(_0293_),
		.dout(new_net_1326)
	);

	bfr new_net_3231_bfr_after (
		.din(_0615_),
		.dout(new_net_3231)
	);

	bfr new_net_3232_bfr_after (
		.din(new_net_3231),
		.dout(new_net_3232)
	);

	bfr new_net_3233_bfr_after (
		.din(new_net_3232),
		.dout(new_net_3233)
	);

	bfr new_net_3234_bfr_after (
		.din(new_net_3233),
		.dout(new_net_3234)
	);

	bfr new_net_3235_bfr_after (
		.din(new_net_3234),
		.dout(new_net_3235)
	);

	bfr new_net_3236_bfr_after (
		.din(new_net_3235),
		.dout(new_net_3236)
	);

	bfr new_net_3237_bfr_after (
		.din(new_net_3236),
		.dout(new_net_3237)
	);

	bfr new_net_3238_bfr_after (
		.din(new_net_3237),
		.dout(new_net_3238)
	);

	bfr new_net_3239_bfr_after (
		.din(new_net_3238),
		.dout(new_net_3239)
	);

	bfr new_net_1410_bfr_after (
		.din(new_net_3239),
		.dout(new_net_1410)
	);

	bfr new_net_1321_bfr_after (
		.din(_0261_),
		.dout(new_net_1321)
	);

	bfr new_net_3240_bfr_after (
		.din(_0522_),
		.dout(new_net_3240)
	);

	bfr new_net_1384_bfr_after (
		.din(new_net_3240),
		.dout(new_net_1384)
	);

	bfr new_net_3241_bfr_after (
		.din(_0046_),
		.dout(new_net_3241)
	);

	bfr new_net_1264_bfr_after (
		.din(new_net_3241),
		.dout(new_net_1264)
	);

	bfr new_net_1285_bfr_after (
		.din(_0134_),
		.dout(new_net_1285)
	);

	bfr new_net_3242_bfr_after (
		.din(_0418_),
		.dout(new_net_3242)
	);

	bfr new_net_3243_bfr_after (
		.din(new_net_3242),
		.dout(new_net_3243)
	);

	bfr new_net_1348_bfr_after (
		.din(new_net_3243),
		.dout(new_net_1348)
	);

	bfr new_net_3244_bfr_after (
		.din(_0604_),
		.dout(new_net_3244)
	);

	bfr new_net_3245_bfr_after (
		.din(new_net_3244),
		.dout(new_net_3245)
	);

	bfr new_net_1406_bfr_after (
		.din(new_net_3245),
		.dout(new_net_1406)
	);

	bfr new_net_1432_bfr_after (
		.din(_0685_),
		.dout(new_net_1432)
	);

	bfr new_net_1370_bfr_after (
		.din(_0483_),
		.dout(new_net_1370)
	);

	bfr new_net_1454_bfr_after (
		.din(_0743_),
		.dout(new_net_1454)
	);

	bfr new_net_1428_bfr_after (
		.din(G46),
		.dout(new_net_1428)
	);

	bfr new_net_3246_bfr_after (
		.din(_0731_),
		.dout(new_net_3246)
	);

	bfr new_net_1449_bfr_after (
		.din(new_net_3246),
		.dout(new_net_1449)
	);

	bfr new_net_1392_bfr_after (
		.din(_0560_),
		.dout(new_net_1392)
	);

	bfr new_net_1366_bfr_after (
		.din(_0476_),
		.dout(new_net_1366)
	);

	bfr new_net_3247_bfr_after (
		.din(_0637_),
		.dout(new_net_3247)
	);

	bfr new_net_3248_bfr_after (
		.din(new_net_3247),
		.dout(new_net_3248)
	);

	bfr new_net_3249_bfr_after (
		.din(new_net_3248),
		.dout(new_net_3249)
	);

	bfr new_net_3250_bfr_after (
		.din(new_net_3249),
		.dout(new_net_3250)
	);

	bfr new_net_3251_bfr_after (
		.din(new_net_3250),
		.dout(new_net_3251)
	);

	bfr new_net_1414_bfr_after (
		.din(new_net_3251),
		.dout(new_net_1414)
	);

	bfr new_net_3252_bfr_after (
		.din(_0537_),
		.dout(new_net_3252)
	);

	bfr new_net_3253_bfr_after (
		.din(new_net_3252),
		.dout(new_net_3253)
	);

	bfr new_net_1388_bfr_after (
		.din(new_net_3253),
		.dout(new_net_1388)
	);

	bfr new_net_3254_bfr_after (
		.din(_0283_),
		.dout(new_net_3254)
	);

	bfr new_net_3255_bfr_after (
		.din(new_net_3254),
		.dout(new_net_3255)
	);

	bfr new_net_1325_bfr_after (
		.din(new_net_3255),
		.dout(new_net_1325)
	);

	bfr new_net_1283_bfr_after (
		.din(_0131_),
		.dout(new_net_1283)
	);

	bfr new_net_1304_bfr_after (
		.din(_0204_),
		.dout(new_net_1304)
	);

	bfr new_net_1262_bfr_after (
		.din(_0026_),
		.dout(new_net_1262)
	);

	bfr new_net_1275_bfr_after (
		.din(_0092_),
		.dout(new_net_1275)
	);

	bfr new_net_1279_bfr_after (
		.din(_0108_),
		.dout(new_net_1279)
	);

	bfr new_net_3256_bfr_after (
		.din(_0177_),
		.dout(new_net_3256)
	);

	bfr new_net_1296_bfr_after (
		.din(new_net_3256),
		.dout(new_net_1296)
	);

	bfr new_net_1317_bfr_after (
		.din(_0249_),
		.dout(new_net_1317)
	);

	bfr new_net_3257_bfr_after (
		.din(G49),
		.dout(new_net_3257)
	);

	bfr new_net_3258_bfr_after (
		.din(new_net_3257),
		.dout(new_net_3258)
	);

	bfr new_net_1268_bfr_after (
		.din(new_net_3258),
		.dout(new_net_1268)
	);

	bfr new_net_3259_bfr_after (
		.din(_0193_),
		.dout(new_net_3259)
	);

	bfr new_net_1300_bfr_after (
		.din(new_net_3259),
		.dout(new_net_1300)
	);

	bfr new_net_3260_bfr_after (
		.din(_0426_),
		.dout(new_net_3260)
	);

	bfr new_net_3261_bfr_after (
		.din(new_net_3260),
		.dout(new_net_3261)
	);

	bfr new_net_1352_bfr_after (
		.din(new_net_3261),
		.dout(new_net_1352)
	);

	bfr new_net_3262_bfr_after (
		.din(_0444_),
		.dout(new_net_3262)
	);

	bfr new_net_1357_bfr_after (
		.din(new_net_3262),
		.dout(new_net_1357)
	);

	bfr new_net_3263_bfr_after (
		.din(_0693_),
		.dout(new_net_3263)
	);

	bfr new_net_1436_bfr_after (
		.din(new_net_3263),
		.dout(new_net_1436)
	);

	bfr new_net_1462_bfr_after (
		.din(_0781_),
		.dout(new_net_1462)
	);

	bfr new_net_3264_bfr_after (
		.din(new_net_1473),
		.dout(new_net_3264)
	);

	bfr new_net_3265_bfr_after (
		.din(new_net_3264),
		.dout(new_net_3265)
	);

	bfr new_net_3266_bfr_after (
		.din(new_net_3265),
		.dout(new_net_3266)
	);

	bfr G3538_bfr_after (
		.din(new_net_3266),
		.dout(G3538)
	);

	bfr new_net_3267_bfr_after (
		.din(_0511_),
		.dout(new_net_3267)
	);

	bfr new_net_3268_bfr_after (
		.din(new_net_3267),
		.dout(new_net_3268)
	);

	bfr new_net_3269_bfr_after (
		.din(new_net_3268),
		.dout(new_net_3269)
	);

	bfr new_net_3270_bfr_after (
		.din(new_net_3269),
		.dout(new_net_3270)
	);

	bfr new_net_3271_bfr_after (
		.din(new_net_3270),
		.dout(new_net_3271)
	);

	bfr new_net_1379_bfr_after (
		.din(new_net_3271),
		.dout(new_net_1379)
	);

	bfr new_net_3272_bfr_after (
		.din(_0498_),
		.dout(new_net_3272)
	);

	bfr new_net_3273_bfr_after (
		.din(new_net_3272),
		.dout(new_net_3273)
	);

	bfr new_net_3274_bfr_after (
		.din(new_net_3273),
		.dout(new_net_3274)
	);

	bfr new_net_3275_bfr_after (
		.din(new_net_3274),
		.dout(new_net_3275)
	);

	bfr new_net_3276_bfr_after (
		.din(new_net_3275),
		.dout(new_net_3276)
	);

	bfr new_net_3277_bfr_after (
		.din(new_net_3276),
		.dout(new_net_3277)
	);

	bfr new_net_3278_bfr_after (
		.din(new_net_3277),
		.dout(new_net_3278)
	);

	bfr new_net_3279_bfr_after (
		.din(new_net_3278),
		.dout(new_net_3279)
	);

	bfr new_net_3280_bfr_after (
		.din(new_net_3279),
		.dout(new_net_3280)
	);

	bfr new_net_3281_bfr_after (
		.din(new_net_3280),
		.dout(new_net_3281)
	);

	bfr new_net_3282_bfr_after (
		.din(new_net_3281),
		.dout(new_net_3282)
	);

	bfr new_net_3283_bfr_after (
		.din(new_net_3282),
		.dout(new_net_3283)
	);

	bfr new_net_3284_bfr_after (
		.din(new_net_3283),
		.dout(new_net_3284)
	);

	bfr new_net_3285_bfr_after (
		.din(new_net_3284),
		.dout(new_net_3285)
	);

	bfr new_net_3286_bfr_after (
		.din(new_net_3285),
		.dout(new_net_3286)
	);

	bfr new_net_3287_bfr_after (
		.din(new_net_3286),
		.dout(new_net_3287)
	);

	bfr new_net_3288_bfr_after (
		.din(new_net_3287),
		.dout(new_net_3288)
	);

	bfr new_net_3289_bfr_after (
		.din(new_net_3288),
		.dout(new_net_3289)
	);

	bfr new_net_3290_bfr_after (
		.din(new_net_3289),
		.dout(new_net_3290)
	);

	bfr new_net_3291_bfr_after (
		.din(new_net_3290),
		.dout(new_net_3291)
	);

	bfr new_net_3292_bfr_after (
		.din(new_net_3291),
		.dout(new_net_3292)
	);

	bfr new_net_3293_bfr_after (
		.din(new_net_3292),
		.dout(new_net_3293)
	);

	bfr new_net_3294_bfr_after (
		.din(new_net_3293),
		.dout(new_net_3294)
	);

	bfr new_net_3295_bfr_after (
		.din(new_net_3294),
		.dout(new_net_3295)
	);

	bfr new_net_1374_bfr_after (
		.din(new_net_3295),
		.dout(new_net_1374)
	);

	bfr new_net_3296_bfr_after (
		.din(_0771_),
		.dout(new_net_3296)
	);

	bfr new_net_3297_bfr_after (
		.din(new_net_3296),
		.dout(new_net_3297)
	);

	bfr new_net_3298_bfr_after (
		.din(new_net_3297),
		.dout(new_net_3298)
	);

	bfr new_net_3299_bfr_after (
		.din(new_net_3298),
		.dout(new_net_3299)
	);

	bfr new_net_3300_bfr_after (
		.din(new_net_3299),
		.dout(new_net_3300)
	);

	bfr new_net_3301_bfr_after (
		.din(new_net_3300),
		.dout(new_net_3301)
	);

	bfr new_net_3302_bfr_after (
		.din(new_net_3301),
		.dout(new_net_3302)
	);

	bfr new_net_3303_bfr_after (
		.din(new_net_3302),
		.dout(new_net_3303)
	);

	bfr new_net_3304_bfr_after (
		.din(new_net_3303),
		.dout(new_net_3304)
	);

	bfr new_net_3305_bfr_after (
		.din(new_net_3304),
		.dout(new_net_3305)
	);

	bfr new_net_3306_bfr_after (
		.din(new_net_3305),
		.dout(new_net_3306)
	);

	bfr new_net_3307_bfr_after (
		.din(new_net_3306),
		.dout(new_net_3307)
	);

	bfr new_net_3308_bfr_after (
		.din(new_net_3307),
		.dout(new_net_3308)
	);

	bfr new_net_3309_bfr_after (
		.din(new_net_3308),
		.dout(new_net_3309)
	);

	bfr new_net_3310_bfr_after (
		.din(new_net_3309),
		.dout(new_net_3310)
	);

	bfr new_net_3311_bfr_after (
		.din(new_net_3310),
		.dout(new_net_3311)
	);

	bfr new_net_3312_bfr_after (
		.din(new_net_3311),
		.dout(new_net_3312)
	);

	bfr new_net_3313_bfr_after (
		.din(new_net_3312),
		.dout(new_net_3313)
	);

	bfr new_net_3314_bfr_after (
		.din(new_net_3313),
		.dout(new_net_3314)
	);

	bfr new_net_3315_bfr_after (
		.din(new_net_3314),
		.dout(new_net_3315)
	);

	bfr new_net_3316_bfr_after (
		.din(new_net_3315),
		.dout(new_net_3316)
	);

	bfr new_net_3317_bfr_after (
		.din(new_net_3316),
		.dout(new_net_3317)
	);

	bfr new_net_3318_bfr_after (
		.din(new_net_3317),
		.dout(new_net_3318)
	);

	bfr new_net_3319_bfr_after (
		.din(new_net_3318),
		.dout(new_net_3319)
	);

	bfr new_net_3320_bfr_after (
		.din(new_net_3319),
		.dout(new_net_3320)
	);

	bfr new_net_3321_bfr_after (
		.din(new_net_3320),
		.dout(new_net_3321)
	);

	bfr new_net_3322_bfr_after (
		.din(new_net_3321),
		.dout(new_net_3322)
	);

	bfr new_net_3323_bfr_after (
		.din(new_net_3322),
		.dout(new_net_3323)
	);

	bfr new_net_1458_bfr_after (
		.din(new_net_3323),
		.dout(new_net_1458)
	);

	bfr new_net_3324_bfr_after (
		.din(_0373_),
		.dout(new_net_3324)
	);

	bfr new_net_1338_bfr_after (
		.din(new_net_3324),
		.dout(new_net_1338)
	);

	bfr new_net_3325_bfr_after (
		.din(_0590_),
		.dout(new_net_3325)
	);

	bfr new_net_3326_bfr_after (
		.din(new_net_3325),
		.dout(new_net_3326)
	);

	bfr new_net_3327_bfr_after (
		.din(new_net_3326),
		.dout(new_net_3327)
	);

	bfr new_net_3328_bfr_after (
		.din(new_net_3327),
		.dout(new_net_3328)
	);

	bfr new_net_3329_bfr_after (
		.din(new_net_3328),
		.dout(new_net_3329)
	);

	bfr new_net_3330_bfr_after (
		.din(new_net_3329),
		.dout(new_net_3330)
	);

	bfr new_net_3331_bfr_after (
		.din(new_net_3330),
		.dout(new_net_3331)
	);

	bfr new_net_1401_bfr_after (
		.din(new_net_3331),
		.dout(new_net_1401)
	);

	bfr new_net_3332_bfr_after (
		.din(_0579_),
		.dout(new_net_3332)
	);

	bfr new_net_3333_bfr_after (
		.din(new_net_3332),
		.dout(new_net_3333)
	);

	bfr new_net_3334_bfr_after (
		.din(new_net_3333),
		.dout(new_net_3334)
	);

	bfr new_net_3335_bfr_after (
		.din(new_net_3334),
		.dout(new_net_3335)
	);

	bfr new_net_3336_bfr_after (
		.din(new_net_3335),
		.dout(new_net_3336)
	);

	bfr new_net_1396_bfr_after (
		.din(new_net_3336),
		.dout(new_net_1396)
	);

	bfr new_net_3337_bfr_after (
		.din(new_net_1471),
		.dout(new_net_3337)
	);

	bfr new_net_3338_bfr_after (
		.din(new_net_3337),
		.dout(new_net_3338)
	);

	bfr new_net_3339_bfr_after (
		.din(new_net_3338),
		.dout(new_net_3339)
	);

	bfr new_net_3340_bfr_after (
		.din(new_net_3339),
		.dout(new_net_3340)
	);

	bfr new_net_3341_bfr_after (
		.din(new_net_3340),
		.dout(new_net_3341)
	);

	bfr new_net_3342_bfr_after (
		.din(new_net_3341),
		.dout(new_net_3342)
	);

	bfr new_net_3343_bfr_after (
		.din(new_net_3342),
		.dout(new_net_3343)
	);

	bfr new_net_3344_bfr_after (
		.din(new_net_3343),
		.dout(new_net_3344)
	);

	bfr new_net_3345_bfr_after (
		.din(new_net_3344),
		.dout(new_net_3345)
	);

	bfr new_net_3346_bfr_after (
		.din(new_net_3345),
		.dout(new_net_3346)
	);

	bfr new_net_3347_bfr_after (
		.din(new_net_3346),
		.dout(new_net_3347)
	);

	bfr new_net_3348_bfr_after (
		.din(new_net_3347),
		.dout(new_net_3348)
	);

	bfr new_net_3349_bfr_after (
		.din(new_net_3348),
		.dout(new_net_3349)
	);

	bfr new_net_3350_bfr_after (
		.din(new_net_3349),
		.dout(new_net_3350)
	);

	bfr new_net_3351_bfr_after (
		.din(new_net_3350),
		.dout(new_net_3351)
	);

	bfr new_net_3352_bfr_after (
		.din(new_net_3351),
		.dout(new_net_3352)
	);

	bfr new_net_3353_bfr_after (
		.din(new_net_3352),
		.dout(new_net_3353)
	);

	bfr new_net_3354_bfr_after (
		.din(new_net_3353),
		.dout(new_net_3354)
	);

	bfr new_net_3355_bfr_after (
		.din(new_net_3354),
		.dout(new_net_3355)
	);

	bfr new_net_3356_bfr_after (
		.din(new_net_3355),
		.dout(new_net_3356)
	);

	bfr new_net_3357_bfr_after (
		.din(new_net_3356),
		.dout(new_net_3357)
	);

	bfr new_net_3358_bfr_after (
		.din(new_net_3357),
		.dout(new_net_3358)
	);

	bfr new_net_3359_bfr_after (
		.din(new_net_3358),
		.dout(new_net_3359)
	);

	bfr new_net_3360_bfr_after (
		.din(new_net_3359),
		.dout(new_net_3360)
	);

	bfr new_net_3361_bfr_after (
		.din(new_net_3360),
		.dout(new_net_3361)
	);

	bfr new_net_3362_bfr_after (
		.din(new_net_3361),
		.dout(new_net_3362)
	);

	bfr new_net_3363_bfr_after (
		.din(new_net_3362),
		.dout(new_net_3363)
	);

	bfr new_net_3364_bfr_after (
		.din(new_net_3363),
		.dout(new_net_3364)
	);

	bfr new_net_3365_bfr_after (
		.din(new_net_3364),
		.dout(new_net_3365)
	);

	bfr G3524_bfr_after (
		.din(new_net_3365),
		.dout(G3524)
	);

	bfr new_net_3366_bfr_after (
		.din(new_net_1483),
		.dout(new_net_3366)
	);

	bfr new_net_3367_bfr_after (
		.din(new_net_3366),
		.dout(new_net_3367)
	);

	bfr new_net_3368_bfr_after (
		.din(new_net_3367),
		.dout(new_net_3368)
	);

	bfr new_net_3369_bfr_after (
		.din(new_net_3368),
		.dout(new_net_3369)
	);

	bfr new_net_3370_bfr_after (
		.din(new_net_3369),
		.dout(new_net_3370)
	);

	bfr new_net_3371_bfr_after (
		.din(new_net_3370),
		.dout(new_net_3371)
	);

	bfr new_net_3372_bfr_after (
		.din(new_net_3371),
		.dout(new_net_3372)
	);

	bfr new_net_3373_bfr_after (
		.din(new_net_3372),
		.dout(new_net_3373)
	);

	bfr new_net_3374_bfr_after (
		.din(new_net_3373),
		.dout(new_net_3374)
	);

	bfr new_net_3375_bfr_after (
		.din(new_net_3374),
		.dout(new_net_3375)
	);

	bfr new_net_3376_bfr_after (
		.din(new_net_3375),
		.dout(new_net_3376)
	);

	bfr new_net_3377_bfr_after (
		.din(new_net_3376),
		.dout(new_net_3377)
	);

	bfr new_net_3378_bfr_after (
		.din(new_net_3377),
		.dout(new_net_3378)
	);

	bfr new_net_3379_bfr_after (
		.din(new_net_3378),
		.dout(new_net_3379)
	);

	bfr new_net_3380_bfr_after (
		.din(new_net_3379),
		.dout(new_net_3380)
	);

	bfr new_net_3381_bfr_after (
		.din(new_net_3380),
		.dout(new_net_3381)
	);

	bfr new_net_3382_bfr_after (
		.din(new_net_3381),
		.dout(new_net_3382)
	);

	bfr new_net_3383_bfr_after (
		.din(new_net_3382),
		.dout(new_net_3383)
	);

	bfr new_net_3384_bfr_after (
		.din(new_net_3383),
		.dout(new_net_3384)
	);

	bfr new_net_3385_bfr_after (
		.din(new_net_3384),
		.dout(new_net_3385)
	);

	bfr new_net_3386_bfr_after (
		.din(new_net_3385),
		.dout(new_net_3386)
	);

	bfr new_net_3387_bfr_after (
		.din(new_net_3386),
		.dout(new_net_3387)
	);

	bfr new_net_3388_bfr_after (
		.din(new_net_3387),
		.dout(new_net_3388)
	);

	bfr new_net_3389_bfr_after (
		.din(new_net_3388),
		.dout(new_net_3389)
	);

	bfr G3527_bfr_after (
		.din(new_net_3389),
		.dout(G3527)
	);

	bfr new_net_3390_bfr_after (
		.din(_0661_),
		.dout(new_net_3390)
	);

	bfr new_net_3391_bfr_after (
		.din(new_net_3390),
		.dout(new_net_3391)
	);

	bfr new_net_3392_bfr_after (
		.din(new_net_3391),
		.dout(new_net_3392)
	);

	bfr new_net_3393_bfr_after (
		.din(new_net_3392),
		.dout(new_net_3393)
	);

	bfr new_net_3394_bfr_after (
		.din(new_net_3393),
		.dout(new_net_3394)
	);

	bfr new_net_3395_bfr_after (
		.din(new_net_3394),
		.dout(new_net_3395)
	);

	bfr new_net_3396_bfr_after (
		.din(new_net_3395),
		.dout(new_net_3396)
	);

	bfr new_net_3397_bfr_after (
		.din(new_net_3396),
		.dout(new_net_3397)
	);

	bfr new_net_3398_bfr_after (
		.din(new_net_3397),
		.dout(new_net_3398)
	);

	bfr new_net_3399_bfr_after (
		.din(new_net_3398),
		.dout(new_net_3399)
	);

	bfr new_net_3400_bfr_after (
		.din(new_net_3399),
		.dout(new_net_3400)
	);

	bfr new_net_3401_bfr_after (
		.din(new_net_3400),
		.dout(new_net_3401)
	);

	bfr new_net_3402_bfr_after (
		.din(new_net_3401),
		.dout(new_net_3402)
	);

	bfr new_net_1423_bfr_after (
		.din(new_net_3402),
		.dout(new_net_1423)
	);

	bfr new_net_1444_bfr_after (
		.din(_0723_),
		.dout(new_net_1444)
	);

	bfr new_net_3403_bfr_after (
		.din(_0330_),
		.dout(new_net_3403)
	);

	bfr new_net_3404_bfr_after (
		.din(new_net_3403),
		.dout(new_net_3404)
	);

	bfr new_net_3405_bfr_after (
		.din(new_net_3404),
		.dout(new_net_3405)
	);

	bfr new_net_3406_bfr_after (
		.din(new_net_3405),
		.dout(new_net_3406)
	);

	bfr new_net_1334_bfr_after (
		.din(new_net_3406),
		.dout(new_net_1334)
	);

	bfr new_net_1418_bfr_after (
		.din(_0649_),
		.dout(new_net_1418)
	);

	bfr new_net_3407_bfr_after (
		.din(_0462_),
		.dout(new_net_3407)
	);

	bfr new_net_3408_bfr_after (
		.din(new_net_3407),
		.dout(new_net_3408)
	);

	bfr new_net_3409_bfr_after (
		.din(new_net_3408),
		.dout(new_net_3409)
	);

	bfr new_net_3410_bfr_after (
		.din(new_net_3409),
		.dout(new_net_3410)
	);

	bfr new_net_3411_bfr_after (
		.din(new_net_3410),
		.dout(new_net_3411)
	);

	bfr new_net_3412_bfr_after (
		.din(new_net_3411),
		.dout(new_net_3412)
	);

	bfr new_net_1361_bfr_after (
		.din(new_net_3412),
		.dout(new_net_1361)
	);

	bfr new_net_1356_bfr_after (
		.din(_0440_),
		.dout(new_net_1356)
	);

	bfr new_net_1440_bfr_after (
		.din(_0707_),
		.dout(new_net_1440)
	);

	bfr new_net_1287_bfr_after (
		.din(_0141_),
		.dout(new_net_1287)
	);

	bfr new_net_1308_bfr_after (
		.din(_0218_),
		.dout(new_net_1308)
	);

	bfr new_net_3413_bfr_after (
		.din(_0301_),
		.dout(new_net_3413)
	);

	bfr new_net_3414_bfr_after (
		.din(new_net_3413),
		.dout(new_net_3414)
	);

	bfr new_net_1329_bfr_after (
		.din(new_net_3414),
		.dout(new_net_1329)
	);

	bfr new_net_1291_bfr_after (
		.din(_0152_),
		.dout(new_net_1291)
	);

	bfr new_net_1312_bfr_after (
		.din(_0227_),
		.dout(new_net_1312)
	);

	bfr new_net_3415_bfr_after (
		.din(_0056_),
		.dout(new_net_3415)
	);

	bfr new_net_3416_bfr_after (
		.din(new_net_3415),
		.dout(new_net_3416)
	);

	bfr new_net_1266_bfr_after (
		.din(new_net_3416),
		.dout(new_net_1266)
	);

	bfr new_net_3417_bfr_after (
		.din(_0077_),
		.dout(new_net_3417)
	);

	bfr new_net_1270_bfr_after (
		.din(new_net_3417),
		.dout(new_net_1270)
	);

	bfr new_net_1333_bfr_after (
		.din(_0329_),
		.dout(new_net_1333)
	);

	bfr new_net_3418_bfr_after (
		.din(_0422_),
		.dout(new_net_3418)
	);

	bfr new_net_3419_bfr_after (
		.din(new_net_3418),
		.dout(new_net_3419)
	);

	bfr new_net_3420_bfr_after (
		.din(new_net_3419),
		.dout(new_net_3420)
	);

	bfr new_net_3421_bfr_after (
		.din(new_net_3420),
		.dout(new_net_3421)
	);

	bfr new_net_3422_bfr_after (
		.din(new_net_3421),
		.dout(new_net_3422)
	);

	bfr new_net_3423_bfr_after (
		.din(new_net_3422),
		.dout(new_net_3423)
	);

	bfr new_net_3424_bfr_after (
		.din(new_net_3423),
		.dout(new_net_3424)
	);

	bfr new_net_1350_bfr_after (
		.din(new_net_3424),
		.dout(new_net_1350)
	);

	bfr new_net_3425_bfr_after (
		.din(_0417_),
		.dout(new_net_3425)
	);

	bfr new_net_3426_bfr_after (
		.din(new_net_3425),
		.dout(new_net_3426)
	);

	bfr new_net_3427_bfr_after (
		.din(new_net_3426),
		.dout(new_net_3427)
	);

	bfr new_net_3428_bfr_after (
		.din(new_net_3427),
		.dout(new_net_3428)
	);

	bfr new_net_3429_bfr_after (
		.din(new_net_3428),
		.dout(new_net_3429)
	);

	bfr new_net_1354_bfr_after (
		.din(new_net_3429),
		.dout(new_net_1354)
	);

	bfr new_net_3430_bfr_after (
		.din(_0523_),
		.dout(new_net_3430)
	);

	bfr new_net_1383_bfr_after (
		.din(new_net_3430),
		.dout(new_net_1383)
	);

	bfr new_net_1347_bfr_after (
		.din(_0353_),
		.dout(new_net_1347)
	);

	bfr new_net_3431_bfr_after (
		.din(_0668_),
		.dout(new_net_3431)
	);

	bfr new_net_1431_bfr_after (
		.din(new_net_3431),
		.dout(new_net_1431)
	);

	bfr new_net_1342_bfr_after (
		.din(_0389_),
		.dout(new_net_1342)
	);

	bfr new_net_3432_bfr_after (
		.din(_0596_),
		.dout(new_net_3432)
	);

	bfr new_net_1405_bfr_after (
		.din(new_net_3432),
		.dout(new_net_1405)
	);

	bfr new_net_1369_bfr_after (
		.din(_0485_),
		.dout(new_net_1369)
	);

	bfr new_net_3433_bfr_after (
		.din(G45),
		.dout(new_net_3433)
	);

	bfr new_net_1427_bfr_after (
		.din(new_net_3433),
		.dout(new_net_1427)
	);

endmodule