module apc32bits(in, out);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _apc16_1_adder1_lv1_a ;
  wire _apc16_1_adder1_lv1_b ;
  wire _apc16_1_adder1_lv1_cin ;
  wire _apc16_1_adder1_lv1_cout ;
  wire _apc16_1_adder1_lv1_d ;
  wire _apc16_1_adder1_lv1_m3_d ;
  wire _apc16_1_adder1_lv2_b ;
  wire _apc16_1_adder1_lv2_cin ;
  wire _apc16_1_adder1_lv2_cout ;
  wire _apc16_1_adder1_lv2_d ;
  wire _apc16_1_adder1_lv2_m3_d ;
  wire _apc16_1_adder2_lv1_a ;
  wire _apc16_1_adder2_lv1_b ;
  wire _apc16_1_adder2_lv1_cin ;
  wire _apc16_1_adder2_lv1_d ;
  wire _apc16_1_adder2_lv1_m3_d ;
  wire _apc16_1_adder2_lv2_cin ;
  wire _apc16_1_adder2_lv2_d ;
  wire _apc16_1_adder2_lv2_m3_d ;
  wire _apc16_1_half1_a ;
  wire _apc16_1_half1_cout ;
  wire _apc16_1_half1_s ;
  wire _apc16_1_half2_cout ;
  wire _apc16_1_half2_s ;
  wire _apc16_1_half3_cout ;
  wire _apc16_1_half3_s ;
  wire _apc16_2_adder1_lv1_a ;
  wire _apc16_2_adder1_lv1_b ;
  wire _apc16_2_adder1_lv1_cin ;
  wire _apc16_2_adder1_lv1_cout ;
  wire _apc16_2_adder1_lv1_d ;
  wire _apc16_2_adder1_lv1_m3_d ;
  wire _apc16_2_adder1_lv2_b ;
  wire _apc16_2_adder1_lv2_cin ;
  wire _apc16_2_adder1_lv2_cout ;
  wire _apc16_2_adder1_lv2_d ;
  wire _apc16_2_adder1_lv2_m3_d ;
  wire _apc16_2_adder2_lv1_a ;
  wire _apc16_2_adder2_lv1_b ;
  wire _apc16_2_adder2_lv1_cin ;
  wire _apc16_2_adder2_lv1_d ;
  wire _apc16_2_adder2_lv1_m3_d ;
  wire _apc16_2_adder2_lv2_cin ;
  wire _apc16_2_adder2_lv2_d ;
  wire _apc16_2_adder2_lv2_m3_d ;
  wire _apc16_2_half1_a ;
  wire _apc16_2_half1_cout ;
  wire _apc16_2_half1_s ;
  wire _apc16_2_half2_cout ;
  wire _apc16_2_half2_s ;
  wire _apc16_2_half3_cout ;
  wire _apc16_2_half3_s ;
  input in_0_;
  input in_1_;
  input in_2_;
  input in_3_;
  input in_4_;
  input in_5_;
  input in_6_;
  input in_7_;
  input in_8_;
  input in_9_;
  input in_10_;
  input in_11_;
  input in_12_;
  input in_13_;
  input in_14_;
  input in_15_;
  input in_16_;
  input in_17_;
  input in_18_;
  input in_19_;
  input in_20_;
  input in_21_;
  input in_22_;
  input in_23_;
  input in_24_;
  input in_25_;
  input in_26_;
  input in_27_;
  input in_28_;
  input in_29_;
  input in_30_;
  input in_31_;
  output out_0_;
  output out_1_;
  output out_2_;
  output out_3_;
  output out_4_;
  output out_5_;
  or_ii _031_ (
    .a(1'b0),
    .b(1'b0),
    .c(_000_)
  );
  and_ii _032_ (
    .a(1'b0),
    .b(1'b0),
    .c(_001_)
  );
  and_bi _033_ (
    .a(_000_),
    .b(_001_),
    .c(out_0_)
  );
  or_ii _034_ (
    .a(_apc16_2_half1_s ),
    .b(_apc16_1_half1_s ),
    .c(_002_)
  );
  and_ii _035_ (
    .a(_apc16_2_half1_s ),
    .b(_apc16_1_half1_s ),
    .c(_003_)
  );
  and_bi _036_ (
    .a(_002_),
    .b(_003_),
    .c(_004_)
  );
  or_bi _037_ (
    .a(_000_),
    .b(_004_),
    .c(_005_)
  );
  and_bi _038_ (
    .a(_000_),
    .b(_004_),
    .c(_006_)
  );
  and_bi _039_ (
    .a(_005_),
    .b(_006_),
    .c(out_1_)
  );
  maj_bii _040_ (
    .a(_000_),
    .b(_apc16_2_half1_s ),
    .c(_apc16_1_half1_s ),
    .d(_007_)
  );
  or_ii _041_ (
    .a(_apc16_2_half2_s ),
    .b(_apc16_1_half2_s ),
    .c(_008_)
  );
  and_ii _042_ (
    .a(_apc16_2_half2_s ),
    .b(_apc16_1_half2_s ),
    .c(_009_)
  );
  and_bi _043_ (
    .a(_008_),
    .b(_009_),
    .c(_010_)
  );
  or_bi _044_ (
    .a(_007_),
    .b(_010_),
    .c(_011_)
  );
  and_bi _045_ (
    .a(_007_),
    .b(_010_),
    .c(_012_)
  );
  and_bi _046_ (
    .a(_011_),
    .b(_012_),
    .c(out_2_)
  );
  maj_bii _047_ (
    .a(_007_),
    .b(_apc16_2_half2_s ),
    .c(_apc16_1_half2_s ),
    .d(_013_)
  );
  or_ii _048_ (
    .a(_apc16_2_half3_s ),
    .b(_apc16_1_half3_s ),
    .c(_014_)
  );
  and_ii _049_ (
    .a(_apc16_2_half3_s ),
    .b(_apc16_1_half3_s ),
    .c(_015_)
  );
  and_bi _050_ (
    .a(_014_),
    .b(_015_),
    .c(_016_)
  );
  or_bi _051_ (
    .a(_013_),
    .b(_016_),
    .c(_017_)
  );
  and_bi _052_ (
    .a(_013_),
    .b(_016_),
    .c(_018_)
  );
  and_bi _053_ (
    .a(_017_),
    .b(_018_),
    .c(out_3_)
  );
  maj_bii _054_ (
    .a(_013_),
    .b(_apc16_2_half3_s ),
    .c(_apc16_1_half3_s ),
    .d(_019_)
  );
  or_ii _055_ (
    .a(_apc16_2_half3_cout ),
    .b(_apc16_1_half3_cout ),
    .c(_020_)
  );
  and_ii _056_ (
    .a(_apc16_2_half3_cout ),
    .b(_apc16_1_half3_cout ),
    .c(_021_)
  );
  and_bi _057_ (
    .a(_020_),
    .b(_021_),
    .c(_022_)
  );
  or_bi _058_ (
    .a(_019_),
    .b(_022_),
    .c(_023_)
  );
  and_bi _059_ (
    .a(_019_),
    .b(_022_),
    .c(_024_)
  );
  and_bi _060_ (
    .a(_023_),
    .b(_024_),
    .c(out_4_)
  );
  maj_bbi _061_ (
    .a(_apc16_2_half3_cout ),
    .b(_apc16_1_half3_cout ),
    .c(_019_),
    .d(out_5_)
  );
  or_bb _062_ (
    .a(in_17_),
    .b(in_16_),
    .c(_apc16_1_adder1_lv1_a )
  );
  and_bb _063_ (
    .a(in_19_),
    .b(in_18_),
    .c(_apc16_1_adder1_lv1_b )
  );
  or_bb _064_ (
    .a(in_21_),
    .b(in_20_),
    .c(_apc16_1_adder1_lv1_cin )
  );
  and_bb _065_ (
    .a(in_23_),
    .b(in_22_),
    .c(_apc16_1_adder2_lv1_a )
  );
  or_bb _066_ (
    .a(in_25_),
    .b(in_24_),
    .c(_apc16_1_adder2_lv1_b )
  );
  and_bb _067_ (
    .a(in_27_),
    .b(in_26_),
    .c(_apc16_1_adder2_lv1_cin )
  );
  or_bb _068_ (
    .a(in_29_),
    .b(in_28_),
    .c(_apc16_1_adder2_lv2_cin )
  );
  and_bb _069_ (
    .a(in_31_),
    .b(in_30_),
    .c(_apc16_1_half1_a )
  );
  maj_bbb _070_ (
    .a(_apc16_1_adder1_lv1_cin ),
    .b(_apc16_1_adder1_lv1_b ),
    .c(_apc16_1_adder1_lv1_a ),
    .d(_apc16_1_adder1_lv1_cout )
  );
  maj_bbi _071_ (
    .a(_apc16_1_adder1_lv1_b ),
    .b(_apc16_1_adder1_lv1_a ),
    .c(_apc16_1_adder1_lv1_cin ),
    .d(_apc16_1_adder1_lv1_d )
  );
  maj_bbi _072_ (
    .a(_apc16_1_adder1_lv1_d ),
    .b(_apc16_1_adder1_lv1_cin ),
    .c(_apc16_1_adder1_lv1_cout ),
    .d(_apc16_1_adder1_lv1_m3_d )
  );
  maj_bbb _073_ (
    .a(_apc16_1_adder1_lv2_cin ),
    .b(_apc16_1_adder1_lv2_b ),
    .c(_apc16_1_adder1_lv1_cout ),
    .d(_apc16_1_adder1_lv2_cout )
  );
  maj_bbi _074_ (
    .a(_apc16_1_adder1_lv2_b ),
    .b(_apc16_1_adder1_lv1_cout ),
    .c(_apc16_1_adder1_lv2_cin ),
    .d(_apc16_1_adder1_lv2_d )
  );
  maj_bbi _075_ (
    .a(_apc16_1_adder1_lv2_d ),
    .b(_apc16_1_adder1_lv2_cin ),
    .c(_apc16_1_adder1_lv2_cout ),
    .d(_apc16_1_adder1_lv2_m3_d )
  );
  maj_bbb _076_ (
    .a(_apc16_1_adder2_lv1_cin ),
    .b(_apc16_1_adder2_lv1_b ),
    .c(_apc16_1_adder2_lv1_a ),
    .d(_apc16_1_adder1_lv2_b )
  );
  maj_bbi _077_ (
    .a(_apc16_1_adder2_lv1_b ),
    .b(_apc16_1_adder2_lv1_a ),
    .c(_apc16_1_adder2_lv1_cin ),
    .d(_apc16_1_adder2_lv1_d )
  );
  maj_bbi _078_ (
    .a(_apc16_1_adder2_lv1_d ),
    .b(_apc16_1_adder2_lv1_cin ),
    .c(_apc16_1_adder1_lv2_b ),
    .d(_apc16_1_adder2_lv1_m3_d )
  );
  maj_bbb _079_ (
    .a(_apc16_1_adder2_lv2_cin ),
    .b(_apc16_1_adder2_lv1_m3_d ),
    .c(_apc16_1_adder1_lv1_m3_d ),
    .d(_apc16_1_adder1_lv2_cin )
  );
  maj_bbi _080_ (
    .a(_apc16_1_adder2_lv1_m3_d ),
    .b(_apc16_1_adder1_lv1_m3_d ),
    .c(_apc16_1_adder2_lv2_cin ),
    .d(_apc16_1_adder2_lv2_d )
  );
  maj_bbi _081_ (
    .a(_apc16_1_adder2_lv2_d ),
    .b(_apc16_1_adder2_lv2_cin ),
    .c(_apc16_1_adder1_lv2_cin ),
    .d(_apc16_1_adder2_lv2_m3_d )
  );
  and_bb _082_ (
    .a(_apc16_1_adder2_lv2_m3_d ),
    .b(_apc16_1_half1_a ),
    .c(_apc16_1_half1_cout )
  );
  or_bb _083_ (
    .a(_apc16_1_adder2_lv2_m3_d ),
    .b(_apc16_1_half1_a ),
    .c(_025_)
  );
  and_bi _084_ (
    .a(_025_),
    .b(_apc16_1_half1_cout ),
    .c(_apc16_1_half1_s )
  );
  and_bb _085_ (
    .a(_apc16_1_half1_cout ),
    .b(_apc16_1_adder1_lv2_m3_d ),
    .c(_apc16_1_half2_cout )
  );
  or_bb _086_ (
    .a(_apc16_1_half1_cout ),
    .b(_apc16_1_adder1_lv2_m3_d ),
    .c(_026_)
  );
  and_bi _087_ (
    .a(_026_),
    .b(_apc16_1_half2_cout ),
    .c(_apc16_1_half2_s )
  );
  and_bb _088_ (
    .a(_apc16_1_half2_cout ),
    .b(_apc16_1_adder1_lv2_cout ),
    .c(_apc16_1_half3_cout )
  );
  or_bb _089_ (
    .a(_apc16_1_half2_cout ),
    .b(_apc16_1_adder1_lv2_cout ),
    .c(_027_)
  );
  and_bi _090_ (
    .a(_027_),
    .b(_apc16_1_half3_cout ),
    .c(_apc16_1_half3_s )
  );
  or_bb _091_ (
    .a(in_1_),
    .b(in_0_),
    .c(_apc16_2_adder1_lv1_a )
  );
  and_bb _092_ (
    .a(in_3_),
    .b(in_2_),
    .c(_apc16_2_adder1_lv1_b )
  );
  or_bb _093_ (
    .a(in_5_),
    .b(in_4_),
    .c(_apc16_2_adder1_lv1_cin )
  );
  and_bb _094_ (
    .a(in_7_),
    .b(in_6_),
    .c(_apc16_2_adder2_lv1_a )
  );
  or_bb _095_ (
    .a(in_9_),
    .b(in_8_),
    .c(_apc16_2_adder2_lv1_b )
  );
  and_bb _096_ (
    .a(in_11_),
    .b(in_10_),
    .c(_apc16_2_adder2_lv1_cin )
  );
  or_bb _097_ (
    .a(in_13_),
    .b(in_12_),
    .c(_apc16_2_adder2_lv2_cin )
  );
  and_bb _098_ (
    .a(in_15_),
    .b(in_14_),
    .c(_apc16_2_half1_a )
  );
  maj_bbb _099_ (
    .a(_apc16_2_adder1_lv1_cin ),
    .b(_apc16_2_adder1_lv1_b ),
    .c(_apc16_2_adder1_lv1_a ),
    .d(_apc16_2_adder1_lv1_cout )
  );
  maj_bbi _100_ (
    .a(_apc16_2_adder1_lv1_b ),
    .b(_apc16_2_adder1_lv1_a ),
    .c(_apc16_2_adder1_lv1_cin ),
    .d(_apc16_2_adder1_lv1_d )
  );
  maj_bbi _101_ (
    .a(_apc16_2_adder1_lv1_d ),
    .b(_apc16_2_adder1_lv1_cin ),
    .c(_apc16_2_adder1_lv1_cout ),
    .d(_apc16_2_adder1_lv1_m3_d )
  );
  maj_bbb _102_ (
    .a(_apc16_2_adder1_lv2_cin ),
    .b(_apc16_2_adder1_lv2_b ),
    .c(_apc16_2_adder1_lv1_cout ),
    .d(_apc16_2_adder1_lv2_cout )
  );
  maj_bbi _103_ (
    .a(_apc16_2_adder1_lv2_b ),
    .b(_apc16_2_adder1_lv1_cout ),
    .c(_apc16_2_adder1_lv2_cin ),
    .d(_apc16_2_adder1_lv2_d )
  );
  maj_bbi _104_ (
    .a(_apc16_2_adder1_lv2_d ),
    .b(_apc16_2_adder1_lv2_cin ),
    .c(_apc16_2_adder1_lv2_cout ),
    .d(_apc16_2_adder1_lv2_m3_d )
  );
  maj_bbb _105_ (
    .a(_apc16_2_adder2_lv1_cin ),
    .b(_apc16_2_adder2_lv1_b ),
    .c(_apc16_2_adder2_lv1_a ),
    .d(_apc16_2_adder1_lv2_b )
  );
  maj_bbi _106_ (
    .a(_apc16_2_adder2_lv1_b ),
    .b(_apc16_2_adder2_lv1_a ),
    .c(_apc16_2_adder2_lv1_cin ),
    .d(_apc16_2_adder2_lv1_d )
  );
  maj_bbi _107_ (
    .a(_apc16_2_adder2_lv1_d ),
    .b(_apc16_2_adder2_lv1_cin ),
    .c(_apc16_2_adder1_lv2_b ),
    .d(_apc16_2_adder2_lv1_m3_d )
  );
  maj_bbb _108_ (
    .a(_apc16_2_adder2_lv2_cin ),
    .b(_apc16_2_adder2_lv1_m3_d ),
    .c(_apc16_2_adder1_lv1_m3_d ),
    .d(_apc16_2_adder1_lv2_cin )
  );
  maj_bbi _109_ (
    .a(_apc16_2_adder2_lv1_m3_d ),
    .b(_apc16_2_adder1_lv1_m3_d ),
    .c(_apc16_2_adder2_lv2_cin ),
    .d(_apc16_2_adder2_lv2_d )
  );
  maj_bbi _110_ (
    .a(_apc16_2_adder2_lv2_d ),
    .b(_apc16_2_adder2_lv2_cin ),
    .c(_apc16_2_adder1_lv2_cin ),
    .d(_apc16_2_adder2_lv2_m3_d )
  );
  and_bb _111_ (
    .a(_apc16_2_adder2_lv2_m3_d ),
    .b(_apc16_2_half1_a ),
    .c(_apc16_2_half1_cout )
  );
  or_bb _112_ (
    .a(_apc16_2_adder2_lv2_m3_d ),
    .b(_apc16_2_half1_a ),
    .c(_028_)
  );
  and_bi _113_ (
    .a(_028_),
    .b(_apc16_2_half1_cout ),
    .c(_apc16_2_half1_s )
  );
  and_bb _114_ (
    .a(_apc16_2_half1_cout ),
    .b(_apc16_2_adder1_lv2_m3_d ),
    .c(_apc16_2_half2_cout )
  );
  or_bb _115_ (
    .a(_apc16_2_half1_cout ),
    .b(_apc16_2_adder1_lv2_m3_d ),
    .c(_029_)
  );
  and_bi _116_ (
    .a(_029_),
    .b(_apc16_2_half2_cout ),
    .c(_apc16_2_half2_s )
  );
  and_bb _117_ (
    .a(_apc16_2_half2_cout ),
    .b(_apc16_2_adder1_lv2_cout ),
    .c(_apc16_2_half3_cout )
  );
  or_bb _118_ (
    .a(_apc16_2_half2_cout ),
    .b(_apc16_2_adder1_lv2_cout ),
    .c(_030_)
  );
  and_bi _119_ (
    .a(_030_),
    .b(_apc16_2_half3_cout ),
    .c(_apc16_2_half3_s )
  );
endmodule
