module ALU32(clock, reset, io_fn, io_in1, io_in2, io_out, io_adder_out, io_test_adder_Cout);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  wire _0913_;
  wire _0914_;
  wire _0915_;
  wire _0916_;
  wire _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  wire _0971_;
  wire _0972_;
  wire _0973_;
  wire _0974_;
  wire _0975_;
  wire _0976_;
  wire _0977_;
  wire _0978_;
  wire _0979_;
  wire _0980_;
  wire _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  wire _0985_;
  wire _0986_;
  wire _0987_;
  wire _0988_;
  wire _0989_;
  wire _0990_;
  wire _0991_;
  wire _0992_;
  wire _0993_;
  wire _0994_;
  wire _0995_;
  wire _0996_;
  wire _0997_;
  wire _0998_;
  wire _0999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire _1031_;
  wire _1032_;
  wire _1033_;
  wire _1034_;
  wire _1035_;
  wire _1036_;
  wire _1037_;
  wire _1038_;
  wire _1039_;
  wire _1040_;
  wire _1041_;
  wire _1042_;
  wire _1043_;
  wire _1044_;
  wire _1045_;
  wire _1046_;
  wire _1047_;
  wire _1048_;
  wire _1049_;
  wire _1050_;
  wire _1051_;
  wire _1052_;
  wire _1053_;
  wire _1054_;
  wire _1055_;
  wire _1056_;
  wire _1057_;
  wire _1058_;
  wire _1059_;
  wire _1060_;
  wire _1061_;
  wire _1062_;
  wire _1063_;
  wire _1064_;
  wire _1065_;
  wire _1066_;
  wire _1067_;
  wire _1068_;
  wire _1069_;
  wire _1070_;
  wire _1071_;
  wire _1072_;
  wire _1073_;
  wire _1074_;
  wire _1075_;
  wire _1076_;
  wire _1077_;
  wire _1078_;
  wire _1079_;
  wire _1080_;
  wire _1081_;
  wire _1082_;
  wire _1083_;
  wire _1084_;
  wire _1085_;
  wire _1086_;
  wire _1087_;
  wire _1088_;
  wire _1089_;
  wire _1090_;
  wire _1091_;
  wire _1092_;
  wire _1093_;
  wire _1094_;
  wire _1095_;
  wire _1096_;
  wire _1097_;
  wire _1098_;
  wire _1099_;
  wire _1100_;
  wire _1101_;
  wire _1102_;
  wire _1103_;
  wire _1104_;
  wire _1105_;
  wire _1106_;
  wire _1107_;
  wire _1108_;
  wire _1109_;
  wire _1110_;
  wire _1111_;
  wire _1112_;
  wire _1113_;
  wire _1114_;
  wire _1115_;
  wire _1116_;
  wire _1117_;
  wire _1118_;
  wire _1119_;
  wire _1120_;
  wire _1121_;
  wire _1122_;
  wire _1123_;
  wire _1124_;
  wire _1125_;
  wire _1126_;
  wire _1127_;
  wire _1128_;
  wire _1129_;
  wire _1130_;
  wire _1131_;
  wire _1132_;
  wire _1133_;
  wire _1134_;
  wire _1135_;
  wire _1136_;
  wire _1137_;
  wire _1138_;
  wire _1139_;
  wire _1140_;
  wire _1141_;
  wire _1142_;
  wire _1143_;
  wire _1144_;
  wire _1145_;
  wire _1146_;
  wire _1147_;
  wire _1148_;
  wire _1149_;
  wire _1150_;
  wire _1151_;
  wire _1152_;
  wire _1153_;
  wire _1154_;
  wire _1155_;
  wire _1156_;
  wire _1157_;
  wire _1158_;
  wire _1159_;
  wire _1160_;
  wire _1161_;
  wire _1162_;
  wire _1163_;
  wire _1164_;
  wire _1165_;
  wire _1166_;
  wire _1167_;
  wire _1168_;
  wire _1169_;
  wire _1170_;
  wire _1171_;
  wire _1172_;
  wire _1173_;
  wire _1174_;
  wire _1175_;
  wire _1176_;
  wire _1177_;
  wire _1178_;
  wire _1179_;
  wire _1180_;
  wire _1181_;
  wire _1182_;
  wire _1183_;
  wire _1184_;
  wire _1185_;
  wire _1186_;
  wire _1187_;
  wire _1188_;
  wire _1189_;
  wire _1190_;
  wire _1191_;
  wire _1192_;
  wire _1193_;
  wire _1194_;
  wire _1195_;
  wire _1196_;
  wire _1197_;
  wire _1198_;
  wire _1199_;
  wire _1200_;
  wire _1201_;
  wire _1202_;
  wire _1203_;
  wire _1204_;
  wire _1205_;
  wire _1206_;
  wire _1207_;
  wire _1208_;
  wire _1209_;
  wire _1210_;
  wire _1211_;
  wire _1212_;
  wire _1213_;
  wire _1214_;
  wire _1215_;
  wire _1216_;
  wire _1217_;
  wire _1218_;
  wire _1219_;
  wire _1220_;
  wire _1221_;
  wire _1222_;
  wire _1223_;
  wire _1224_;
  wire _1225_;
  wire _1226_;
  wire _1227_;
  wire _1228_;
  wire _1229_;
  wire _1230_;
  wire _1231_;
  wire _1232_;
  wire _1233_;
  wire _1234_;
  wire _1235_;
  wire _1236_;
  wire _1237_;
  wire _1238_;
  wire _1239_;
  wire _1240_;
  wire _1241_;
  wire _1242_;
  wire _1243_;
  wire _1244_;
  wire _1245_;
  wire _1246_;
  wire _1247_;
  wire _1248_;
  wire _1249_;
  wire _1250_;
  wire _1251_;
  wire _1252_;
  wire _1253_;
  wire _1254_;
  wire _1255_;
  wire _1256_;
  wire _1257_;
  wire _1258_;
  wire _1259_;
  wire _1260_;
  wire _1261_;
  wire _1262_;
  wire _1263_;
  wire _1264_;
  wire _1265_;
  wire _1266_;
  wire _1267_;
  wire _1268_;
  wire _1269_;
  wire _1270_;
  wire _1271_;
  wire _1272_;
  wire _1273_;
  wire _1274_;
  wire _1275_;
  wire _1276_;
  wire _1277_;
  wire _1278_;
  wire _1279_;
  wire _1280_;
  wire _1281_;
  wire _1282_;
  wire _1283_;
  wire _1284_;
  wire _1285_;
  wire _1286_;
  wire _1287_;
  wire _1288_;
  wire _1289_;
  wire _1290_;
  wire _1291_;
  wire _1292_;
  wire _1293_;
  wire _1294_;
  wire _1295_;
  wire _1296_;
  wire _1297_;
  wire _1298_;
  wire _1299_;
  wire _1300_;
  wire _1301_;
  wire _1302_;
  wire _1303_;
  wire _1304_;
  wire _1305_;
  wire _1306_;
  wire _1307_;
  wire _1308_;
  wire _1309_;
  wire _1310_;
  wire _1311_;
  wire _1312_;
  wire _1313_;
  wire _1314_;
  wire _1315_;
  wire _1316_;
  wire _1317_;
  wire _1318_;
  wire _1319_;
  wire _1320_;
  wire _1321_;
  wire _1322_;
  wire _1323_;
  wire _1324_;
  wire _1325_;
  wire _1326_;
  wire _1327_;
  wire _1328_;
  wire _1329_;
  wire _1330_;
  wire _1331_;
  wire _1332_;
  wire _1333_;
  wire _1334_;
  wire _1335_;
  wire _1336_;
  wire _1337_;
  wire _1338_;
  wire _1339_;
  wire _1340_;
  wire _1341_;
  wire _1342_;
  wire _1343_;
  wire _1344_;
  wire _1345_;
  wire _1346_;
  wire _1347_;
  wire _1348_;
  wire _1349_;
  wire _1350_;
  wire _1351_;
  wire _1352_;
  wire _1353_;
  wire _1354_;
  wire _1355_;
  wire _1356_;
  wire _1357_;
  wire _1358_;
  wire _1359_;
  wire _1360_;
  wire _1361_;
  wire _1362_;
  wire _1363_;
  wire _1364_;
  wire _1365_;
  wire _1366_;
  wire _1367_;
  wire _1368_;
  wire _1369_;
  wire _1370_;
  wire _1371_;
  wire _1372_;
  wire _1373_;
  wire _1374_;
  wire _1375_;
  wire _1376_;
  wire _1377_;
  wire _1378_;
  wire _1379_;
  wire _1380_;
  wire _1381_;
  wire _1382_;
  wire _1383_;
  wire _1384_;
  wire _1385_;
  wire _1386_;
  wire _1387_;
  wire _1388_;
  wire _1389_;
  wire _1390_;
  wire _1391_;
  wire _1392_;
  wire _1393_;
  wire _1394_;
  wire _1395_;
  wire _1396_;
  wire _1397_;
  wire _1398_;
  wire _1399_;
  wire _1400_;
  wire _1401_;
  wire _1402_;
  wire _1403_;
  wire _1404_;
  wire _1405_;
  wire _1406_;
  wire _1407_;
  wire _1408_;
  wire _1409_;
  wire _1410_;
  wire _1411_;
  wire _1412_;
  wire _1413_;
  wire _1414_;
  wire _1415_;
  wire _1416_;
  wire _1417_;
  wire _1418_;
  wire _1419_;
  wire _1420_;
  wire _1421_;
  wire _1422_;
  wire _1423_;
  wire _1424_;
  wire _1425_;
  wire _1426_;
  wire _1427_;
  wire _1428_;
  wire _1429_;
  wire _1430_;
  wire _1431_;
  wire _1432_;
  wire _1433_;
  wire _1434_;
  wire _1435_;
  wire _1436_;
  wire _1437_;
  wire _1438_;
  wire _1439_;
  wire _1440_;
  wire _1441_;
  wire _1442_;
  wire _1443_;
  wire _1444_;
  wire _1445_;
  wire _1446_;
  wire _1447_;
  wire _1448_;
  wire _1449_;
  wire _1450_;
  wire _1451_;
  wire _1452_;
  wire _1453_;
  wire _1454_;
  wire _1455_;
  wire _1456_;
  wire _1457_;
  wire _1458_;
  wire _1459_;
  wire _1460_;
  wire _1461_;
  wire _1462_;
  wire _1463_;
  wire _1464_;
  wire _1465_;
  wire _1466_;
  wire _1467_;
  wire _1468_;
  wire _1469_;
  wire _1470_;
  wire _1471_;
  wire _1472_;
  wire _1473_;
  wire _1474_;
  wire _1475_;
  wire _1476_;
  wire _1477_;
  wire _1478_;
  wire _1479_;
  wire _1480_;
  wire _1481_;
  wire _1482_;
  wire _1483_;
  wire _1484_;
  wire _1485_;
  wire _1486_;
  wire _1487_;
  wire _1488_;
  wire _1489_;
  wire _1490_;
  wire _1491_;
  wire _1492_;
  wire _1493_;
  wire _1494_;
  wire _1495_;
  wire _1496_;
  wire _1497_;
  wire _1498_;
  wire _1499_;
  wire _1500_;
  wire _1501_;
  wire _1502_;
  wire _1503_;
  wire _1504_;
  wire _1505_;
  wire _1506_;
  wire _1507_;
  wire _1508_;
  wire _1509_;
  wire _1510_;
  wire _1511_;
  wire _1512_;
  wire _1513_;
  wire _1514_;
  wire _1515_;
  wire _1516_;
  wire _1517_;
  output io_adder_out_0_;
  output io_adder_out_1_;
  output io_adder_out_2_;
  output io_adder_out_3_;
  output io_adder_out_4_;
  output io_adder_out_5_;
  output io_adder_out_6_;
  output io_adder_out_7_;
  output io_adder_out_8_;
  output io_adder_out_9_;
  output io_adder_out_10_;
  output io_adder_out_11_;
  output io_adder_out_12_;
  output io_adder_out_13_;
  output io_adder_out_14_;
  output io_adder_out_15_;
  output io_adder_out_16_;
  output io_adder_out_17_;
  output io_adder_out_18_;
  output io_adder_out_19_;
  output io_adder_out_20_;
  output io_adder_out_21_;
  output io_adder_out_22_;
  output io_adder_out_23_;
  output io_adder_out_24_;
  output io_adder_out_25_;
  output io_adder_out_26_;
  output io_adder_out_27_;
  output io_adder_out_28_;
  output io_adder_out_29_;
  output io_adder_out_30_;
  output io_adder_out_31_;
  input io_fn_0_;
  input io_fn_1_;
  input io_fn_2_;
  input io_fn_3_;
  input io_in1_0_;
  input io_in1_1_;
  input io_in1_2_;
  input io_in1_3_;
  input io_in1_4_;
  input io_in1_5_;
  input io_in1_6_;
  input io_in1_7_;
  input io_in1_8_;
  input io_in1_9_;
  input io_in1_10_;
  input io_in1_11_;
  input io_in1_12_;
  input io_in1_13_;
  input io_in1_14_;
  input io_in1_15_;
  input io_in1_16_;
  input io_in1_17_;
  input io_in1_18_;
  input io_in1_19_;
  input io_in1_20_;
  input io_in1_21_;
  input io_in1_22_;
  input io_in1_23_;
  input io_in1_24_;
  input io_in1_25_;
  input io_in1_26_;
  input io_in1_27_;
  input io_in1_28_;
  input io_in1_29_;
  input io_in1_30_;
  input io_in1_31_;
  input io_in2_0_;
  input io_in2_1_;
  input io_in2_2_;
  input io_in2_3_;
  input io_in2_4_;
  input io_in2_5_;
  input io_in2_6_;
  input io_in2_7_;
  input io_in2_8_;
  input io_in2_9_;
  input io_in2_10_;
  input io_in2_11_;
  input io_in2_12_;
  input io_in2_13_;
  input io_in2_14_;
  input io_in2_15_;
  input io_in2_16_;
  input io_in2_17_;
  input io_in2_18_;
  input io_in2_19_;
  input io_in2_20_;
  input io_in2_21_;
  input io_in2_22_;
  input io_in2_23_;
  input io_in2_24_;
  input io_in2_25_;
  input io_in2_26_;
  input io_in2_27_;
  input io_in2_28_;
  input io_in2_29_;
  input io_in2_30_;
  input io_in2_31_;
  output io_out_0_;
  output io_out_1_;
  output io_out_2_;
  output io_out_3_;
  output io_out_4_;
  output io_out_5_;
  output io_out_6_;
  output io_out_7_;
  output io_out_8_;
  output io_out_9_;
  output io_out_10_;
  output io_out_11_;
  output io_out_12_;
  output io_out_13_;
  output io_out_14_;
  output io_out_15_;
  output io_out_16_;
  output io_out_17_;
  output io_out_18_;
  output io_out_19_;
  output io_out_20_;
  output io_out_21_;
  output io_out_22_;
  output io_out_23_;
  output io_out_24_;
  output io_out_25_;
  output io_out_26_;
  output io_out_27_;
  output io_out_28_;
  output io_out_29_;
  output io_out_30_;
  output io_out_31_;
  output io_test_adder_Cout;

  inv _1518_ (
    .din(io_in1_31_),
    .dout(_0340_)
  );
  inv _1519_ (
    .din(io_in2_31_),
    .dout(_0341_)
  );
  inv _1520_ (
    .din(io_fn_3_),
    .dout(_0352_)
  );
  inv _1521_ (
    .din(io_in2_29_),
    .dout(_0363_)
  );
  inv _1522_ (
    .din(io_in2_2_),
    .dout(_0383_)
  );
  or_bb _1523_ (
    .a(io_in2_1_),
    .b(io_in2_0_),
    .c(_0384_)
  );
  and_bi _1524_ (
    .a(_0383_),
    .b(_0384_),
    .c(_0394_)
  );
  and_bi _1525_ (
    .a(_0394_),
    .b(io_in2_3_),
    .c(_0405_)
  );
  and_bi _1526_ (
    .a(_0405_),
    .b(io_in2_4_),
    .c(_0415_)
  );
  and_bi _1527_ (
    .a(_0415_),
    .b(io_in2_5_),
    .c(_0436_)
  );
  and_bi _1528_ (
    .a(_0436_),
    .b(io_in2_6_),
    .c(_0437_)
  );
  and_bi _1529_ (
    .a(_0437_),
    .b(io_in2_7_),
    .c(_0447_)
  );
  and_bi _1530_ (
    .a(_0447_),
    .b(io_in2_8_),
    .c(_0458_)
  );
  and_bi _1531_ (
    .a(_0458_),
    .b(io_in2_9_),
    .c(_0477_)
  );
  and_bi _1532_ (
    .a(_0477_),
    .b(io_in2_10_),
    .c(_0478_)
  );
  and_bi _1533_ (
    .a(_0478_),
    .b(io_in2_11_),
    .c(_0489_)
  );
  and_bi _1534_ (
    .a(_0489_),
    .b(io_in2_12_),
    .c(_0499_)
  );
  and_bi _1535_ (
    .a(_0499_),
    .b(io_in2_13_),
    .c(_0510_)
  );
  and_bi _1536_ (
    .a(_0510_),
    .b(io_in2_14_),
    .c(_0530_)
  );
  and_bi _1537_ (
    .a(_0530_),
    .b(io_in2_15_),
    .c(_0531_)
  );
  and_bi _1538_ (
    .a(_0531_),
    .b(io_in2_16_),
    .c(_0541_)
  );
  and_bi _1539_ (
    .a(_0541_),
    .b(io_in2_17_),
    .c(_0551_)
  );
  and_bi _1540_ (
    .a(_0551_),
    .b(io_in2_18_),
    .c(_0571_)
  );
  and_bi _1541_ (
    .a(_0571_),
    .b(io_in2_19_),
    .c(_0572_)
  );
  and_bi _1542_ (
    .a(_0572_),
    .b(io_in2_20_),
    .c(_0583_)
  );
  and_bi _1543_ (
    .a(_0583_),
    .b(io_in2_21_),
    .c(_0593_)
  );
  and_bi _1544_ (
    .a(_0593_),
    .b(io_in2_22_),
    .c(_0603_)
  );
  and_bi _1545_ (
    .a(_0603_),
    .b(io_in2_23_),
    .c(_0623_)
  );
  and_bi _1546_ (
    .a(_0623_),
    .b(io_in2_24_),
    .c(_0624_)
  );
  and_bi _1547_ (
    .a(_0624_),
    .b(io_in2_25_),
    .c(_0635_)
  );
  and_bi _1548_ (
    .a(_0635_),
    .b(io_in2_26_),
    .c(_0645_)
  );
  and_bi _1549_ (
    .a(_0645_),
    .b(io_in2_27_),
    .c(_0665_)
  );
  or_bb _1550_ (
    .a(_0665_),
    .b(_0352_),
    .c(_0666_)
  );
  and_bi _1551_ (
    .a(_0666_),
    .b(io_in2_28_),
    .c(_0676_)
  );
  and_bi _1552_ (
    .a(io_fn_3_),
    .b(_0676_),
    .c(_0687_)
  );
  and_bi _1553_ (
    .a(_0363_),
    .b(_0687_),
    .c(_0697_)
  );
  or_bb _1554_ (
    .a(_0697_),
    .b(_0352_),
    .c(_0717_)
  );
  and_bb _1555_ (
    .a(io_in2_30_),
    .b(io_fn_3_),
    .c(_0718_)
  );
  and_bi _1556_ (
    .a(_0717_),
    .b(_0718_),
    .c(_0725_)
  );
  and_bi _1557_ (
    .a(_0341_),
    .b(_0725_),
    .c(_0726_)
  );
  and_bi _1558_ (
    .a(_0725_),
    .b(_0341_),
    .c(_0727_)
  );
  or_bb _1559_ (
    .a(_0727_),
    .b(_0726_),
    .c(_0728_)
  );
  and_bi _1560_ (
    .a(_0728_),
    .b(_0340_),
    .c(_0729_)
  );
  inv _1561_ (
    .din(_0729_),
    .dout(_0730_)
  );
  and_bi _1562_ (
    .a(_0340_),
    .b(_0728_),
    .c(_0731_)
  );
  and_bi _1563_ (
    .a(_0730_),
    .b(_0731_),
    .c(_0732_)
  );
  inv _1564_ (
    .din(io_in1_30_),
    .dout(_0733_)
  );
  inv _1565_ (
    .din(io_in1_27_),
    .dout(_0734_)
  );
  inv _1566_ (
    .din(io_in1_26_),
    .dout(_0735_)
  );
  inv _1567_ (
    .din(io_in1_25_),
    .dout(_0736_)
  );
  inv _1568_ (
    .din(io_in1_23_),
    .dout(_0737_)
  );
  inv _1569_ (
    .din(io_in1_17_),
    .dout(_0738_)
  );
  inv _1570_ (
    .din(io_in1_13_),
    .dout(_0739_)
  );
  inv _1571_ (
    .din(io_in1_11_),
    .dout(_0740_)
  );
  inv _1572_ (
    .din(io_in1_7_),
    .dout(_0741_)
  );
  inv _1573_ (
    .din(io_in1_1_),
    .dout(_0742_)
  );
  and_bb _1574_ (
    .a(io_in2_0_),
    .b(io_in1_0_),
    .c(_0743_)
  );
  and_bi _1575_ (
    .a(_0742_),
    .b(_0743_),
    .c(_0744_)
  );
  or_ii _1576_ (
    .a(_0743_),
    .b(io_in1_1_),
    .c(_0745_)
  );
  and_bi _1577_ (
    .a(io_in2_1_),
    .b(io_fn_3_),
    .c(_0746_)
  );
  or_ii _1578_ (
    .a(io_in2_1_),
    .b(io_in2_0_),
    .c(_0747_)
  );
  or_ii _1579_ (
    .a(_0384_),
    .b(io_fn_3_),
    .c(_0748_)
  );
  and_bi _1580_ (
    .a(_0747_),
    .b(_0748_),
    .c(_0749_)
  );
  or_bb _1581_ (
    .a(_0749_),
    .b(_0746_),
    .c(_0750_)
  );
  and_bi _1582_ (
    .a(_0745_),
    .b(_0750_),
    .c(_0751_)
  );
  or_bb _1583_ (
    .a(_0751_),
    .b(_0744_),
    .c(_0752_)
  );
  and_bi _1584_ (
    .a(_0752_),
    .b(io_in1_2_),
    .c(_0753_)
  );
  inv _1585_ (
    .din(io_in1_2_),
    .dout(_0754_)
  );
  or_bb _1586_ (
    .a(_0752_),
    .b(_0754_),
    .c(_0755_)
  );
  and_bi _1587_ (
    .a(_0383_),
    .b(_0748_),
    .c(_0756_)
  );
  and_bi _1588_ (
    .a(_0748_),
    .b(_0383_),
    .c(_0757_)
  );
  or_bb _1589_ (
    .a(_0757_),
    .b(_0756_),
    .c(_0758_)
  );
  and_bi _1590_ (
    .a(_0755_),
    .b(_0758_),
    .c(_0759_)
  );
  or_bb _1591_ (
    .a(_0759_),
    .b(_0753_),
    .c(_0760_)
  );
  and_bi _1592_ (
    .a(_0760_),
    .b(io_in1_3_),
    .c(_0761_)
  );
  inv _1593_ (
    .din(io_in1_3_),
    .dout(_0762_)
  );
  or_bb _1594_ (
    .a(_0760_),
    .b(_0762_),
    .c(_0763_)
  );
  inv _1595_ (
    .din(io_in2_3_),
    .dout(_0764_)
  );
  and_bi _1596_ (
    .a(io_fn_3_),
    .b(_0394_),
    .c(_0765_)
  );
  and_bi _1597_ (
    .a(_0765_),
    .b(_0764_),
    .c(_0766_)
  );
  and_bi _1598_ (
    .a(_0764_),
    .b(_0765_),
    .c(_0767_)
  );
  or_bb _1599_ (
    .a(_0767_),
    .b(_0766_),
    .c(_0768_)
  );
  inv _1600_ (
    .din(_0768_),
    .dout(_0769_)
  );
  and_bi _1601_ (
    .a(_0763_),
    .b(_0769_),
    .c(_0770_)
  );
  or_bb _1602_ (
    .a(_0770_),
    .b(_0761_),
    .c(_0771_)
  );
  and_bi _1603_ (
    .a(_0771_),
    .b(io_in1_4_),
    .c(_0772_)
  );
  inv _1604_ (
    .din(io_in1_4_),
    .dout(_0773_)
  );
  or_bb _1605_ (
    .a(_0771_),
    .b(_0773_),
    .c(_0774_)
  );
  and_bi _1606_ (
    .a(io_fn_3_),
    .b(_0405_),
    .c(_0775_)
  );
  and_bi _1607_ (
    .a(_0775_),
    .b(io_in2_4_),
    .c(_0776_)
  );
  and_bi _1608_ (
    .a(io_in2_4_),
    .b(_0775_),
    .c(_0777_)
  );
  or_bb _1609_ (
    .a(_0777_),
    .b(_0776_),
    .c(_0778_)
  );
  and_bi _1610_ (
    .a(_0774_),
    .b(_0778_),
    .c(_0779_)
  );
  or_bb _1611_ (
    .a(_0779_),
    .b(_0772_),
    .c(_0780_)
  );
  and_bi _1612_ (
    .a(_0780_),
    .b(io_in1_5_),
    .c(_0781_)
  );
  inv _1613_ (
    .din(io_in1_5_),
    .dout(_0782_)
  );
  or_bb _1614_ (
    .a(_0780_),
    .b(_0782_),
    .c(_0783_)
  );
  inv _1615_ (
    .din(io_in2_5_),
    .dout(_0784_)
  );
  and_bi _1616_ (
    .a(io_fn_3_),
    .b(_0415_),
    .c(_0785_)
  );
  and_bi _1617_ (
    .a(_0785_),
    .b(_0784_),
    .c(_0786_)
  );
  and_bi _1618_ (
    .a(_0784_),
    .b(_0785_),
    .c(_0787_)
  );
  or_bb _1619_ (
    .a(_0787_),
    .b(_0786_),
    .c(_0788_)
  );
  inv _1620_ (
    .din(_0788_),
    .dout(_0789_)
  );
  and_bi _1621_ (
    .a(_0783_),
    .b(_0789_),
    .c(_0790_)
  );
  or_bb _1622_ (
    .a(_0790_),
    .b(_0781_),
    .c(_0791_)
  );
  and_bi _1623_ (
    .a(io_in1_6_),
    .b(_0791_),
    .c(_0792_)
  );
  inv _1624_ (
    .din(io_in1_6_),
    .dout(_0793_)
  );
  or_ii _1625_ (
    .a(_0791_),
    .b(_0793_),
    .c(_0794_)
  );
  and_bi _1626_ (
    .a(io_fn_3_),
    .b(_0436_),
    .c(_0795_)
  );
  and_bi _1627_ (
    .a(_0795_),
    .b(io_in2_6_),
    .c(_0796_)
  );
  and_bi _1628_ (
    .a(io_in2_6_),
    .b(_0795_),
    .c(_0797_)
  );
  or_bb _1629_ (
    .a(_0797_),
    .b(_0796_),
    .c(_0798_)
  );
  and_bb _1630_ (
    .a(_0798_),
    .b(_0794_),
    .c(_0799_)
  );
  or_bb _1631_ (
    .a(_0799_),
    .b(_0792_),
    .c(_0800_)
  );
  and_bi _1632_ (
    .a(_0741_),
    .b(_0800_),
    .c(_0801_)
  );
  or_ii _1633_ (
    .a(_0800_),
    .b(io_in1_7_),
    .c(_0802_)
  );
  inv _1634_ (
    .din(io_in2_7_),
    .dout(_0803_)
  );
  and_bi _1635_ (
    .a(io_fn_3_),
    .b(_0437_),
    .c(_0804_)
  );
  and_bi _1636_ (
    .a(_0804_),
    .b(_0803_),
    .c(_0805_)
  );
  and_bi _1637_ (
    .a(_0803_),
    .b(_0804_),
    .c(_0806_)
  );
  or_bb _1638_ (
    .a(_0806_),
    .b(_0805_),
    .c(_0807_)
  );
  inv _1639_ (
    .din(_0807_),
    .dout(_0808_)
  );
  and_bi _1640_ (
    .a(_0802_),
    .b(_0808_),
    .c(_0809_)
  );
  or_bb _1641_ (
    .a(_0809_),
    .b(_0801_),
    .c(_0810_)
  );
  and_bi _1642_ (
    .a(_0810_),
    .b(io_in1_8_),
    .c(_0811_)
  );
  inv _1643_ (
    .din(io_in1_8_),
    .dout(_0812_)
  );
  or_bb _1644_ (
    .a(_0810_),
    .b(_0812_),
    .c(_0813_)
  );
  and_bi _1645_ (
    .a(io_fn_3_),
    .b(_0447_),
    .c(_0814_)
  );
  and_bi _1646_ (
    .a(_0814_),
    .b(io_in2_8_),
    .c(_0815_)
  );
  and_bi _1647_ (
    .a(io_in2_8_),
    .b(_0814_),
    .c(_0816_)
  );
  or_bb _1648_ (
    .a(_0816_),
    .b(_0815_),
    .c(_0817_)
  );
  and_bi _1649_ (
    .a(_0813_),
    .b(_0817_),
    .c(_0818_)
  );
  or_bb _1650_ (
    .a(_0818_),
    .b(_0811_),
    .c(_0819_)
  );
  and_bi _1651_ (
    .a(_0819_),
    .b(io_in1_9_),
    .c(_0820_)
  );
  inv _1652_ (
    .din(io_in1_9_),
    .dout(_0821_)
  );
  or_bb _1653_ (
    .a(_0819_),
    .b(_0821_),
    .c(_0822_)
  );
  inv _1654_ (
    .din(io_in2_9_),
    .dout(_0823_)
  );
  and_bi _1655_ (
    .a(io_fn_3_),
    .b(_0458_),
    .c(_0824_)
  );
  and_bi _1656_ (
    .a(_0824_),
    .b(_0823_),
    .c(_0825_)
  );
  and_bi _1657_ (
    .a(_0823_),
    .b(_0824_),
    .c(_0826_)
  );
  or_bb _1658_ (
    .a(_0826_),
    .b(_0825_),
    .c(_0827_)
  );
  inv _1659_ (
    .din(_0827_),
    .dout(_0828_)
  );
  and_bi _1660_ (
    .a(_0822_),
    .b(_0828_),
    .c(_0829_)
  );
  or_bb _1661_ (
    .a(_0829_),
    .b(_0820_),
    .c(_0830_)
  );
  and_bi _1662_ (
    .a(_0830_),
    .b(io_in1_10_),
    .c(_0831_)
  );
  inv _1663_ (
    .din(io_in1_10_),
    .dout(_0832_)
  );
  or_bb _1664_ (
    .a(_0830_),
    .b(_0832_),
    .c(_0833_)
  );
  and_bi _1665_ (
    .a(io_fn_3_),
    .b(_0477_),
    .c(_0834_)
  );
  and_bi _1666_ (
    .a(_0834_),
    .b(io_in2_10_),
    .c(_0835_)
  );
  and_bi _1667_ (
    .a(io_in2_10_),
    .b(_0834_),
    .c(_0836_)
  );
  or_bb _1668_ (
    .a(_0836_),
    .b(_0835_),
    .c(_0837_)
  );
  and_bi _1669_ (
    .a(_0833_),
    .b(_0837_),
    .c(_0838_)
  );
  or_bb _1670_ (
    .a(_0838_),
    .b(_0831_),
    .c(_0839_)
  );
  or_ii _1671_ (
    .a(_0839_),
    .b(_0740_),
    .c(_0840_)
  );
  or_bb _1672_ (
    .a(_0839_),
    .b(_0740_),
    .c(_0841_)
  );
  and_bi _1673_ (
    .a(io_fn_3_),
    .b(_0478_),
    .c(_0842_)
  );
  or_ii _1674_ (
    .a(_0842_),
    .b(io_in2_11_),
    .c(_0843_)
  );
  inv _1675_ (
    .din(io_in2_11_),
    .dout(_0844_)
  );
  and_bi _1676_ (
    .a(_0844_),
    .b(_0842_),
    .c(_0845_)
  );
  and_bi _1677_ (
    .a(_0843_),
    .b(_0845_),
    .c(_0846_)
  );
  and_bi _1678_ (
    .a(_0841_),
    .b(_0846_),
    .c(_0847_)
  );
  or_bi _1679_ (
    .a(_0847_),
    .b(_0840_),
    .c(_0848_)
  );
  and_bi _1680_ (
    .a(_0848_),
    .b(io_in1_12_),
    .c(_0849_)
  );
  inv _1681_ (
    .din(io_in1_12_),
    .dout(_0850_)
  );
  or_bb _1682_ (
    .a(_0848_),
    .b(_0850_),
    .c(_0851_)
  );
  and_bi _1683_ (
    .a(io_fn_3_),
    .b(_0489_),
    .c(_0852_)
  );
  and_bi _1684_ (
    .a(_0852_),
    .b(io_in2_12_),
    .c(_0853_)
  );
  and_bi _1685_ (
    .a(io_in2_12_),
    .b(_0852_),
    .c(_0854_)
  );
  or_bb _1686_ (
    .a(_0854_),
    .b(_0853_),
    .c(_0855_)
  );
  and_bi _1687_ (
    .a(_0851_),
    .b(_0855_),
    .c(_0856_)
  );
  or_bb _1688_ (
    .a(_0856_),
    .b(_0849_),
    .c(_0857_)
  );
  or_ii _1689_ (
    .a(_0857_),
    .b(_0739_),
    .c(_0858_)
  );
  or_bb _1690_ (
    .a(_0857_),
    .b(_0739_),
    .c(_0859_)
  );
  and_bi _1691_ (
    .a(io_fn_3_),
    .b(_0499_),
    .c(_0860_)
  );
  or_ii _1692_ (
    .a(_0860_),
    .b(io_in2_13_),
    .c(_0861_)
  );
  inv _1693_ (
    .din(io_in2_13_),
    .dout(_0862_)
  );
  and_bi _1694_ (
    .a(_0862_),
    .b(_0860_),
    .c(_0863_)
  );
  and_bi _1695_ (
    .a(_0861_),
    .b(_0863_),
    .c(_0864_)
  );
  and_bi _1696_ (
    .a(_0859_),
    .b(_0864_),
    .c(_0865_)
  );
  or_bi _1697_ (
    .a(_0865_),
    .b(_0858_),
    .c(_0866_)
  );
  and_bi _1698_ (
    .a(_0866_),
    .b(io_in1_14_),
    .c(_0867_)
  );
  inv _1699_ (
    .din(io_in1_14_),
    .dout(_0868_)
  );
  or_bb _1700_ (
    .a(_0866_),
    .b(_0868_),
    .c(_0869_)
  );
  and_bi _1701_ (
    .a(io_fn_3_),
    .b(_0510_),
    .c(_0870_)
  );
  and_bi _1702_ (
    .a(_0870_),
    .b(io_in2_14_),
    .c(_0871_)
  );
  and_bi _1703_ (
    .a(io_in2_14_),
    .b(_0870_),
    .c(_0872_)
  );
  or_bb _1704_ (
    .a(_0872_),
    .b(_0871_),
    .c(_0873_)
  );
  and_bi _1705_ (
    .a(_0869_),
    .b(_0873_),
    .c(_0874_)
  );
  or_bb _1706_ (
    .a(_0874_),
    .b(_0867_),
    .c(_0875_)
  );
  and_bi _1707_ (
    .a(_0875_),
    .b(io_in1_15_),
    .c(_0876_)
  );
  inv _1708_ (
    .din(io_in1_15_),
    .dout(_0877_)
  );
  or_bb _1709_ (
    .a(_0875_),
    .b(_0877_),
    .c(_0878_)
  );
  inv _1710_ (
    .din(io_in2_15_),
    .dout(_0879_)
  );
  and_bi _1711_ (
    .a(io_fn_3_),
    .b(_0530_),
    .c(_0880_)
  );
  and_bi _1712_ (
    .a(_0880_),
    .b(_0879_),
    .c(_0881_)
  );
  and_bi _1713_ (
    .a(_0879_),
    .b(_0880_),
    .c(_0882_)
  );
  or_bb _1714_ (
    .a(_0882_),
    .b(_0881_),
    .c(_0883_)
  );
  inv _1715_ (
    .din(_0883_),
    .dout(_0884_)
  );
  and_bi _1716_ (
    .a(_0878_),
    .b(_0884_),
    .c(_0885_)
  );
  or_bb _1717_ (
    .a(_0885_),
    .b(_0876_),
    .c(_0886_)
  );
  and_bi _1718_ (
    .a(io_in1_16_),
    .b(_0886_),
    .c(_0887_)
  );
  inv _1719_ (
    .din(io_in1_16_),
    .dout(_0888_)
  );
  or_ii _1720_ (
    .a(_0886_),
    .b(_0888_),
    .c(_0889_)
  );
  and_bi _1721_ (
    .a(io_fn_3_),
    .b(_0531_),
    .c(_0890_)
  );
  and_bi _1722_ (
    .a(_0890_),
    .b(io_in2_16_),
    .c(_0891_)
  );
  and_bi _1723_ (
    .a(io_in2_16_),
    .b(_0890_),
    .c(_0892_)
  );
  or_bb _1724_ (
    .a(_0892_),
    .b(_0891_),
    .c(_0893_)
  );
  and_bb _1725_ (
    .a(_0893_),
    .b(_0889_),
    .c(_0894_)
  );
  or_bb _1726_ (
    .a(_0894_),
    .b(_0887_),
    .c(_0895_)
  );
  and_bi _1727_ (
    .a(_0895_),
    .b(_0738_),
    .c(_0896_)
  );
  or_bb _1728_ (
    .a(_0895_),
    .b(io_in1_17_),
    .c(_0897_)
  );
  inv _1729_ (
    .din(io_in2_17_),
    .dout(_0898_)
  );
  and_bi _1730_ (
    .a(io_fn_3_),
    .b(_0541_),
    .c(_0899_)
  );
  and_bi _1731_ (
    .a(_0899_),
    .b(_0898_),
    .c(_0900_)
  );
  and_bi _1732_ (
    .a(_0898_),
    .b(_0899_),
    .c(_0901_)
  );
  or_bb _1733_ (
    .a(_0901_),
    .b(_0900_),
    .c(_0902_)
  );
  and_bi _1734_ (
    .a(_0897_),
    .b(_0902_),
    .c(_0903_)
  );
  or_bb _1735_ (
    .a(_0903_),
    .b(_0896_),
    .c(_0904_)
  );
  or_ii _1736_ (
    .a(_0904_),
    .b(io_in1_18_),
    .c(_0905_)
  );
  or_bb _1737_ (
    .a(_0904_),
    .b(io_in1_18_),
    .c(_0906_)
  );
  and_bi _1738_ (
    .a(io_fn_3_),
    .b(_0551_),
    .c(_0907_)
  );
  and_bi _1739_ (
    .a(_0907_),
    .b(io_in2_18_),
    .c(_0908_)
  );
  and_bi _1740_ (
    .a(io_in2_18_),
    .b(_0907_),
    .c(_0909_)
  );
  or_bb _1741_ (
    .a(_0909_),
    .b(_0908_),
    .c(_0910_)
  );
  and_bb _1742_ (
    .a(_0910_),
    .b(_0906_),
    .c(_0911_)
  );
  and_bi _1743_ (
    .a(_0905_),
    .b(_0911_),
    .c(_0912_)
  );
  and_bi _1744_ (
    .a(_0912_),
    .b(io_in1_19_),
    .c(_0913_)
  );
  inv _1745_ (
    .din(io_in1_19_),
    .dout(_0914_)
  );
  or_bb _1746_ (
    .a(_0912_),
    .b(_0914_),
    .c(_0915_)
  );
  inv _1747_ (
    .din(io_in2_19_),
    .dout(_0916_)
  );
  and_bi _1748_ (
    .a(io_fn_3_),
    .b(_0571_),
    .c(_0917_)
  );
  and_bi _1749_ (
    .a(_0917_),
    .b(_0916_),
    .c(_0918_)
  );
  and_bi _1750_ (
    .a(_0916_),
    .b(_0917_),
    .c(_0919_)
  );
  or_bb _1751_ (
    .a(_0919_),
    .b(_0918_),
    .c(_0920_)
  );
  inv _1752_ (
    .din(_0920_),
    .dout(_0921_)
  );
  and_bi _1753_ (
    .a(_0915_),
    .b(_0921_),
    .c(_0922_)
  );
  or_bb _1754_ (
    .a(_0922_),
    .b(_0913_),
    .c(_0923_)
  );
  and_bi _1755_ (
    .a(_0923_),
    .b(io_in1_20_),
    .c(_0924_)
  );
  inv _1756_ (
    .din(io_in1_20_),
    .dout(_0925_)
  );
  or_bb _1757_ (
    .a(_0923_),
    .b(_0925_),
    .c(_0926_)
  );
  and_bi _1758_ (
    .a(io_fn_3_),
    .b(_0572_),
    .c(_0927_)
  );
  and_bi _1759_ (
    .a(_0927_),
    .b(io_in2_20_),
    .c(_0928_)
  );
  and_bi _1760_ (
    .a(io_in2_20_),
    .b(_0927_),
    .c(_0929_)
  );
  or_bb _1761_ (
    .a(_0929_),
    .b(_0928_),
    .c(_0930_)
  );
  and_bi _1762_ (
    .a(_0926_),
    .b(_0930_),
    .c(_0931_)
  );
  or_bb _1763_ (
    .a(_0931_),
    .b(_0924_),
    .c(_0932_)
  );
  and_bi _1764_ (
    .a(_0932_),
    .b(io_in1_21_),
    .c(_0933_)
  );
  inv _1765_ (
    .din(io_in1_21_),
    .dout(_0934_)
  );
  or_bb _1766_ (
    .a(_0932_),
    .b(_0934_),
    .c(_0935_)
  );
  inv _1767_ (
    .din(io_in2_21_),
    .dout(_0936_)
  );
  and_bi _1768_ (
    .a(io_fn_3_),
    .b(_0583_),
    .c(_0937_)
  );
  and_bi _1769_ (
    .a(_0937_),
    .b(_0936_),
    .c(_0938_)
  );
  and_bi _1770_ (
    .a(_0936_),
    .b(_0937_),
    .c(_0939_)
  );
  or_bb _1771_ (
    .a(_0939_),
    .b(_0938_),
    .c(_0940_)
  );
  inv _1772_ (
    .din(_0940_),
    .dout(_0941_)
  );
  and_bi _1773_ (
    .a(_0935_),
    .b(_0941_),
    .c(_0942_)
  );
  or_bb _1774_ (
    .a(_0942_),
    .b(_0933_),
    .c(_0943_)
  );
  and_bi _1775_ (
    .a(io_in1_22_),
    .b(_0943_),
    .c(_0944_)
  );
  inv _1776_ (
    .din(io_in1_22_),
    .dout(_0945_)
  );
  or_ii _1777_ (
    .a(_0943_),
    .b(_0945_),
    .c(_0946_)
  );
  and_bi _1778_ (
    .a(io_fn_3_),
    .b(_0593_),
    .c(_0947_)
  );
  and_bi _1779_ (
    .a(_0947_),
    .b(io_in2_22_),
    .c(_0948_)
  );
  and_bi _1780_ (
    .a(io_in2_22_),
    .b(_0947_),
    .c(_0949_)
  );
  or_bb _1781_ (
    .a(_0949_),
    .b(_0948_),
    .c(_0950_)
  );
  and_bb _1782_ (
    .a(_0950_),
    .b(_0946_),
    .c(_0951_)
  );
  or_bb _1783_ (
    .a(_0951_),
    .b(_0944_),
    .c(_0952_)
  );
  and_bi _1784_ (
    .a(_0737_),
    .b(_0952_),
    .c(_0953_)
  );
  or_ii _1785_ (
    .a(_0952_),
    .b(io_in1_23_),
    .c(_0954_)
  );
  inv _1786_ (
    .din(io_in2_23_),
    .dout(_0955_)
  );
  and_bi _1787_ (
    .a(io_fn_3_),
    .b(_0603_),
    .c(_0956_)
  );
  and_bi _1788_ (
    .a(_0956_),
    .b(_0955_),
    .c(_0957_)
  );
  and_bi _1789_ (
    .a(_0955_),
    .b(_0956_),
    .c(_0958_)
  );
  or_bb _1790_ (
    .a(_0958_),
    .b(_0957_),
    .c(_0959_)
  );
  inv _1791_ (
    .din(_0959_),
    .dout(_0960_)
  );
  and_bi _1792_ (
    .a(_0954_),
    .b(_0960_),
    .c(_0961_)
  );
  or_bb _1793_ (
    .a(_0961_),
    .b(_0953_),
    .c(_0962_)
  );
  and_bi _1794_ (
    .a(io_in1_24_),
    .b(_0962_),
    .c(_0963_)
  );
  inv _1795_ (
    .din(io_in1_24_),
    .dout(_0964_)
  );
  or_ii _1796_ (
    .a(_0962_),
    .b(_0964_),
    .c(_0965_)
  );
  and_bi _1797_ (
    .a(io_fn_3_),
    .b(_0623_),
    .c(_0966_)
  );
  and_bi _1798_ (
    .a(_0966_),
    .b(io_in2_24_),
    .c(_0967_)
  );
  and_bi _1799_ (
    .a(io_in2_24_),
    .b(_0966_),
    .c(_0968_)
  );
  or_bb _1800_ (
    .a(_0968_),
    .b(_0967_),
    .c(_0969_)
  );
  and_bb _1801_ (
    .a(_0969_),
    .b(_0965_),
    .c(_0970_)
  );
  or_bb _1802_ (
    .a(_0970_),
    .b(_0963_),
    .c(_0971_)
  );
  and_bi _1803_ (
    .a(_0971_),
    .b(_0736_),
    .c(_0972_)
  );
  inv _1804_ (
    .din(_0972_),
    .dout(_0973_)
  );
  or_bb _1805_ (
    .a(_0971_),
    .b(io_in1_25_),
    .c(_0974_)
  );
  and_bi _1806_ (
    .a(io_fn_3_),
    .b(_0624_),
    .c(_0975_)
  );
  and_bi _1807_ (
    .a(io_in2_25_),
    .b(_0975_),
    .c(_0976_)
  );
  and_bi _1808_ (
    .a(_0975_),
    .b(io_in2_25_),
    .c(_0977_)
  );
  or_bb _1809_ (
    .a(_0977_),
    .b(_0976_),
    .c(_0978_)
  );
  and_bb _1810_ (
    .a(_0978_),
    .b(_0974_),
    .c(_0979_)
  );
  and_bi _1811_ (
    .a(_0973_),
    .b(_0979_),
    .c(_0980_)
  );
  or_bb _1812_ (
    .a(_0980_),
    .b(_0735_),
    .c(_0981_)
  );
  or_ii _1813_ (
    .a(_0980_),
    .b(_0735_),
    .c(_0982_)
  );
  or_bb _1814_ (
    .a(_0635_),
    .b(_0352_),
    .c(_0983_)
  );
  and_bi _1815_ (
    .a(io_in2_26_),
    .b(_0983_),
    .c(_0984_)
  );
  and_bi _1816_ (
    .a(_0983_),
    .b(io_in2_26_),
    .c(_0985_)
  );
  or_bb _1817_ (
    .a(_0985_),
    .b(_0984_),
    .c(_0986_)
  );
  and_bi _1818_ (
    .a(_0982_),
    .b(_0986_),
    .c(_0987_)
  );
  and_bi _1819_ (
    .a(_0981_),
    .b(_0987_),
    .c(_0988_)
  );
  or_ii _1820_ (
    .a(_0988_),
    .b(_0734_),
    .c(_0989_)
  );
  or_bb _1821_ (
    .a(_0988_),
    .b(_0734_),
    .c(_0990_)
  );
  or_bb _1822_ (
    .a(_0645_),
    .b(_0352_),
    .c(_0991_)
  );
  or_bb _1823_ (
    .a(_0991_),
    .b(io_in2_27_),
    .c(_0992_)
  );
  or_ii _1824_ (
    .a(_0991_),
    .b(io_in2_27_),
    .c(_0993_)
  );
  or_ii _1825_ (
    .a(_0993_),
    .b(_0992_),
    .c(_0994_)
  );
  and_bi _1826_ (
    .a(_0990_),
    .b(_0994_),
    .c(_0995_)
  );
  and_bi _1827_ (
    .a(_0989_),
    .b(_0995_),
    .c(_0996_)
  );
  or_ii _1828_ (
    .a(_0996_),
    .b(io_in1_28_),
    .c(_0997_)
  );
  or_bb _1829_ (
    .a(_0996_),
    .b(io_in1_28_),
    .c(_0998_)
  );
  and_bi _1830_ (
    .a(io_in2_28_),
    .b(_0666_),
    .c(_0999_)
  );
  or_bb _1831_ (
    .a(_0999_),
    .b(_0676_),
    .c(_1000_)
  );
  and_bi _1832_ (
    .a(_0998_),
    .b(_1000_),
    .c(_1001_)
  );
  and_bi _1833_ (
    .a(_0997_),
    .b(_1001_),
    .c(_1002_)
  );
  and_bi _1834_ (
    .a(_1002_),
    .b(io_in1_29_),
    .c(_1003_)
  );
  inv _1835_ (
    .din(io_in1_29_),
    .dout(_1004_)
  );
  or_bb _1836_ (
    .a(_1002_),
    .b(_1004_),
    .c(_1005_)
  );
  and_bi _1837_ (
    .a(_0687_),
    .b(_0363_),
    .c(_1006_)
  );
  or_bb _1838_ (
    .a(_1006_),
    .b(_0697_),
    .c(_1007_)
  );
  inv _1839_ (
    .din(_1007_),
    .dout(_1008_)
  );
  and_bi _1840_ (
    .a(_1005_),
    .b(_1008_),
    .c(_1009_)
  );
  or_bb _1841_ (
    .a(_1009_),
    .b(_1003_),
    .c(_1010_)
  );
  or_bb _1842_ (
    .a(_1010_),
    .b(_0733_),
    .c(_1011_)
  );
  and_bi _1843_ (
    .a(_1010_),
    .b(io_in1_30_),
    .c(_1012_)
  );
  and_bi _1844_ (
    .a(io_in2_30_),
    .b(_0717_),
    .c(_1013_)
  );
  and_bi _1845_ (
    .a(_0717_),
    .b(io_in2_30_),
    .c(_1014_)
  );
  or_bb _1846_ (
    .a(_1014_),
    .b(_1013_),
    .c(_1015_)
  );
  inv _1847_ (
    .din(_1015_),
    .dout(_1016_)
  );
  and_bi _1848_ (
    .a(_1016_),
    .b(_1012_),
    .c(_1017_)
  );
  or_bi _1849_ (
    .a(_1017_),
    .b(_1011_),
    .c(_1018_)
  );
  and_bi _1850_ (
    .a(_1018_),
    .b(_0732_),
    .c(_1019_)
  );
  and_bi _1851_ (
    .a(_0732_),
    .b(_1018_),
    .c(_1020_)
  );
  or_bb _1852_ (
    .a(_1020_),
    .b(_1019_),
    .c(io_adder_out_31_)
  );
  and_bi _1853_ (
    .a(_1011_),
    .b(_1012_),
    .c(_1021_)
  );
  or_bb _1854_ (
    .a(_1021_),
    .b(_1016_),
    .c(_1022_)
  );
  and_bb _1855_ (
    .a(_1017_),
    .b(_1011_),
    .c(_1023_)
  );
  and_bi _1856_ (
    .a(_1022_),
    .b(_1023_),
    .c(io_adder_out_30_)
  );
  and_bi _1857_ (
    .a(_1005_),
    .b(_1003_),
    .c(_1024_)
  );
  and_bi _1858_ (
    .a(_1008_),
    .b(_1024_),
    .c(_1025_)
  );
  and_bi _1859_ (
    .a(_1024_),
    .b(_1008_),
    .c(_1026_)
  );
  or_bb _1860_ (
    .a(_1026_),
    .b(_1025_),
    .c(io_adder_out_29_)
  );
  and_bb _1861_ (
    .a(_0998_),
    .b(_0997_),
    .c(_1027_)
  );
  and_bi _1862_ (
    .a(_1000_),
    .b(_1027_),
    .c(_1028_)
  );
  or_ii _1863_ (
    .a(_1001_),
    .b(_0997_),
    .c(_1029_)
  );
  and_bi _1864_ (
    .a(_1029_),
    .b(_1028_),
    .c(io_adder_out_28_)
  );
  and_bb _1865_ (
    .a(_0990_),
    .b(_0989_),
    .c(_1030_)
  );
  and_bi _1866_ (
    .a(_0994_),
    .b(_1030_),
    .c(_1031_)
  );
  and_bb _1867_ (
    .a(_0995_),
    .b(_0989_),
    .c(_1032_)
  );
  or_bb _1868_ (
    .a(_1032_),
    .b(_1031_),
    .c(io_adder_out_27_)
  );
  and_bb _1869_ (
    .a(_0982_),
    .b(_0981_),
    .c(_1033_)
  );
  or_ii _1870_ (
    .a(_1033_),
    .b(_0986_),
    .c(_1034_)
  );
  or_bb _1871_ (
    .a(_1033_),
    .b(_0986_),
    .c(_1035_)
  );
  or_ii _1872_ (
    .a(_1035_),
    .b(_1034_),
    .c(io_adder_out_26_)
  );
  and_bi _1873_ (
    .a(_0974_),
    .b(_0972_),
    .c(_1036_)
  );
  or_bb _1874_ (
    .a(_1036_),
    .b(_0978_),
    .c(_1037_)
  );
  and_bb _1875_ (
    .a(_1036_),
    .b(_0978_),
    .c(_1038_)
  );
  and_bi _1876_ (
    .a(_1037_),
    .b(_1038_),
    .c(io_adder_out_25_)
  );
  and_bi _1877_ (
    .a(_0965_),
    .b(_0963_),
    .c(_1039_)
  );
  or_bb _1878_ (
    .a(_1039_),
    .b(_0969_),
    .c(_1040_)
  );
  and_bb _1879_ (
    .a(_1039_),
    .b(_0969_),
    .c(_1041_)
  );
  and_bi _1880_ (
    .a(_1040_),
    .b(_1041_),
    .c(io_adder_out_24_)
  );
  and_bi _1881_ (
    .a(_0954_),
    .b(_0953_),
    .c(_1042_)
  );
  and_bi _1882_ (
    .a(_1042_),
    .b(_0960_),
    .c(_1043_)
  );
  and_bi _1883_ (
    .a(_0960_),
    .b(_1042_),
    .c(_1044_)
  );
  or_bb _1884_ (
    .a(_1044_),
    .b(_1043_),
    .c(io_adder_out_23_)
  );
  and_bi _1885_ (
    .a(_0946_),
    .b(_0944_),
    .c(_1045_)
  );
  or_bb _1886_ (
    .a(_1045_),
    .b(_0950_),
    .c(_1046_)
  );
  and_bb _1887_ (
    .a(_1045_),
    .b(_0950_),
    .c(_1047_)
  );
  and_bi _1888_ (
    .a(_1046_),
    .b(_1047_),
    .c(io_adder_out_22_)
  );
  and_bi _1889_ (
    .a(_0935_),
    .b(_0933_),
    .c(_1048_)
  );
  and_bi _1890_ (
    .a(_0941_),
    .b(_1048_),
    .c(_1049_)
  );
  and_bi _1891_ (
    .a(_1048_),
    .b(_0941_),
    .c(_1050_)
  );
  or_bb _1892_ (
    .a(_1050_),
    .b(_1049_),
    .c(io_adder_out_21_)
  );
  and_bi _1893_ (
    .a(_0926_),
    .b(_0924_),
    .c(_1051_)
  );
  or_bb _1894_ (
    .a(_1051_),
    .b(_0930_),
    .c(_1052_)
  );
  and_bb _1895_ (
    .a(_1051_),
    .b(_0930_),
    .c(_1053_)
  );
  and_bi _1896_ (
    .a(_1052_),
    .b(_1053_),
    .c(io_adder_out_20_)
  );
  and_bi _1897_ (
    .a(_0915_),
    .b(_0913_),
    .c(_1054_)
  );
  and_bi _1898_ (
    .a(_1054_),
    .b(_0921_),
    .c(_1055_)
  );
  and_bi _1899_ (
    .a(_0921_),
    .b(_1054_),
    .c(_1056_)
  );
  or_bb _1900_ (
    .a(_1056_),
    .b(_1055_),
    .c(io_adder_out_19_)
  );
  and_bb _1901_ (
    .a(_0906_),
    .b(_0905_),
    .c(_1057_)
  );
  and_bi _1902_ (
    .a(_1057_),
    .b(_0910_),
    .c(_1058_)
  );
  and_bi _1903_ (
    .a(_0910_),
    .b(_1057_),
    .c(_1059_)
  );
  or_bb _1904_ (
    .a(_1059_),
    .b(_1058_),
    .c(io_adder_out_18_)
  );
  and_bi _1905_ (
    .a(_0897_),
    .b(_0896_),
    .c(_1060_)
  );
  or_ii _1906_ (
    .a(_1060_),
    .b(_0902_),
    .c(_1061_)
  );
  or_bb _1907_ (
    .a(_1060_),
    .b(_0902_),
    .c(_1062_)
  );
  or_ii _1908_ (
    .a(_1062_),
    .b(_1061_),
    .c(io_adder_out_17_)
  );
  and_bi _1909_ (
    .a(_0889_),
    .b(_0887_),
    .c(_1063_)
  );
  or_bb _1910_ (
    .a(_1063_),
    .b(_0893_),
    .c(_1064_)
  );
  and_bb _1911_ (
    .a(_1063_),
    .b(_0893_),
    .c(_1065_)
  );
  and_bi _1912_ (
    .a(_1064_),
    .b(_1065_),
    .c(io_adder_out_16_)
  );
  and_bi _1913_ (
    .a(_0878_),
    .b(_0876_),
    .c(_1066_)
  );
  and_bi _1914_ (
    .a(_0884_),
    .b(_1066_),
    .c(_1067_)
  );
  and_bi _1915_ (
    .a(_1066_),
    .b(_0884_),
    .c(_1068_)
  );
  or_bb _1916_ (
    .a(_1068_),
    .b(_1067_),
    .c(io_adder_out_15_)
  );
  and_bi _1917_ (
    .a(_0869_),
    .b(_0867_),
    .c(_1069_)
  );
  or_ii _1918_ (
    .a(_1069_),
    .b(_0873_),
    .c(_1070_)
  );
  or_bb _1919_ (
    .a(_1069_),
    .b(_0873_),
    .c(_1071_)
  );
  and_bb _1920_ (
    .a(_1071_),
    .b(_1070_),
    .c(io_adder_out_14_)
  );
  and_bb _1921_ (
    .a(_0865_),
    .b(_0858_),
    .c(_1072_)
  );
  and_bb _1922_ (
    .a(_0859_),
    .b(_0858_),
    .c(_1073_)
  );
  and_bi _1923_ (
    .a(_0864_),
    .b(_1073_),
    .c(_1074_)
  );
  or_bb _1924_ (
    .a(_1074_),
    .b(_1072_),
    .c(io_adder_out_13_)
  );
  and_bi _1925_ (
    .a(_0851_),
    .b(_0849_),
    .c(_1075_)
  );
  or_ii _1926_ (
    .a(_1075_),
    .b(_0855_),
    .c(_1076_)
  );
  or_bb _1927_ (
    .a(_1075_),
    .b(_0855_),
    .c(_1077_)
  );
  and_bb _1928_ (
    .a(_1077_),
    .b(_1076_),
    .c(io_adder_out_12_)
  );
  and_bb _1929_ (
    .a(_0847_),
    .b(_0840_),
    .c(_1078_)
  );
  and_bb _1930_ (
    .a(_0841_),
    .b(_0840_),
    .c(_1079_)
  );
  and_bi _1931_ (
    .a(_0846_),
    .b(_1079_),
    .c(_1080_)
  );
  or_bb _1932_ (
    .a(_1080_),
    .b(_1078_),
    .c(io_adder_out_11_)
  );
  and_bi _1933_ (
    .a(_0833_),
    .b(_0831_),
    .c(_1081_)
  );
  or_bb _1934_ (
    .a(_1081_),
    .b(_0837_),
    .c(_1082_)
  );
  and_bb _1935_ (
    .a(_1081_),
    .b(_0837_),
    .c(_1083_)
  );
  and_bi _1936_ (
    .a(_1082_),
    .b(_1083_),
    .c(io_adder_out_10_)
  );
  and_bi _1937_ (
    .a(_0822_),
    .b(_0820_),
    .c(_1084_)
  );
  and_bi _1938_ (
    .a(_0828_),
    .b(_1084_),
    .c(_1085_)
  );
  and_bi _1939_ (
    .a(_1084_),
    .b(_0828_),
    .c(_1086_)
  );
  or_bb _1940_ (
    .a(_1086_),
    .b(_1085_),
    .c(io_adder_out_9_)
  );
  and_bi _1941_ (
    .a(_0813_),
    .b(_0811_),
    .c(_1087_)
  );
  or_bb _1942_ (
    .a(_1087_),
    .b(_0817_),
    .c(_1088_)
  );
  and_bb _1943_ (
    .a(_1087_),
    .b(_0817_),
    .c(_1089_)
  );
  and_bi _1944_ (
    .a(_1088_),
    .b(_1089_),
    .c(io_adder_out_8_)
  );
  and_bi _1945_ (
    .a(_0802_),
    .b(_0801_),
    .c(_1090_)
  );
  and_bi _1946_ (
    .a(_1090_),
    .b(_0808_),
    .c(_1091_)
  );
  and_bi _1947_ (
    .a(_0808_),
    .b(_1090_),
    .c(_1092_)
  );
  or_bb _1948_ (
    .a(_1092_),
    .b(_1091_),
    .c(io_adder_out_7_)
  );
  and_bi _1949_ (
    .a(_0794_),
    .b(_0792_),
    .c(_1093_)
  );
  or_bb _1950_ (
    .a(_1093_),
    .b(_0798_),
    .c(_1094_)
  );
  and_bb _1951_ (
    .a(_1093_),
    .b(_0798_),
    .c(_1095_)
  );
  and_bi _1952_ (
    .a(_1094_),
    .b(_1095_),
    .c(io_adder_out_6_)
  );
  and_bi _1953_ (
    .a(_0783_),
    .b(_0781_),
    .c(_1096_)
  );
  and_bi _1954_ (
    .a(_0789_),
    .b(_1096_),
    .c(_1097_)
  );
  and_bi _1955_ (
    .a(_1096_),
    .b(_0789_),
    .c(_1098_)
  );
  or_bb _1956_ (
    .a(_1098_),
    .b(_1097_),
    .c(io_adder_out_5_)
  );
  and_bi _1957_ (
    .a(_0774_),
    .b(_0772_),
    .c(_1099_)
  );
  or_bb _1958_ (
    .a(_1099_),
    .b(_0778_),
    .c(_1100_)
  );
  and_bb _1959_ (
    .a(_1099_),
    .b(_0778_),
    .c(_1101_)
  );
  and_bi _1960_ (
    .a(_1100_),
    .b(_1101_),
    .c(io_adder_out_4_)
  );
  and_bi _1961_ (
    .a(_0763_),
    .b(_0761_),
    .c(_1102_)
  );
  and_bi _1962_ (
    .a(_0769_),
    .b(_1102_),
    .c(_1103_)
  );
  and_bi _1963_ (
    .a(_1102_),
    .b(_0769_),
    .c(_1104_)
  );
  or_bb _1964_ (
    .a(_1104_),
    .b(_1103_),
    .c(io_adder_out_3_)
  );
  and_bi _1965_ (
    .a(_0755_),
    .b(_0753_),
    .c(_1105_)
  );
  and_bi _1966_ (
    .a(_0758_),
    .b(_1105_),
    .c(_1106_)
  );
  and_bi _1967_ (
    .a(_1105_),
    .b(_0758_),
    .c(_1107_)
  );
  or_bb _1968_ (
    .a(_1107_),
    .b(_1106_),
    .c(io_adder_out_2_)
  );
  and_bi _1969_ (
    .a(_0745_),
    .b(_0744_),
    .c(_1108_)
  );
  or_bb _1970_ (
    .a(_1108_),
    .b(_0750_),
    .c(_1109_)
  );
  and_bb _1971_ (
    .a(_1108_),
    .b(_0750_),
    .c(_1110_)
  );
  and_bi _1972_ (
    .a(_1109_),
    .b(_1110_),
    .c(io_adder_out_1_)
  );
  inv _1973_ (
    .din(_0743_),
    .dout(_1111_)
  );
  inv _1974_ (
    .din(io_in1_0_),
    .dout(_1112_)
  );
  and_bi _1975_ (
    .a(_1112_),
    .b(io_in2_0_),
    .c(_1113_)
  );
  and_bi _1976_ (
    .a(_1111_),
    .b(_1113_),
    .c(io_adder_out_0_)
  );
  or_bb _1977_ (
    .a(_1018_),
    .b(_0729_),
    .c(_1114_)
  );
  and_bi _1978_ (
    .a(_1114_),
    .b(_0731_),
    .c(io_test_adder_Cout)
  );
  or_bi _1979_ (
    .a(io_fn_0_),
    .b(io_fn_3_),
    .c(_1115_)
  );
  or_bi _1980_ (
    .a(io_fn_2_),
    .b(io_fn_1_),
    .c(_1116_)
  );
  or_bb _1981_ (
    .a(_1116_),
    .b(_1115_),
    .c(_1117_)
  );
  or_bb _1982_ (
    .a(io_fn_2_),
    .b(io_fn_3_),
    .c(_1118_)
  );
  or_bb _1983_ (
    .a(io_fn_1_),
    .b(io_fn_0_),
    .c(_1119_)
  );
  or_bb _1984_ (
    .a(_1119_),
    .b(_1118_),
    .c(_1120_)
  );
  and_bb _1985_ (
    .a(_1120_),
    .b(_1117_),
    .c(_1121_)
  );
  or_bb _1986_ (
    .a(_1121_),
    .b(io_adder_out_0_),
    .c(_1122_)
  );
  and_bi _1987_ (
    .a(io_fn_2_),
    .b(_1115_),
    .c(_1123_)
  );
  and_bi _1988_ (
    .a(io_in1_31_),
    .b(io_in2_31_),
    .c(_1124_)
  );
  and_bi _1989_ (
    .a(io_in2_31_),
    .b(io_in1_31_),
    .c(_1125_)
  );
  or_bb _1990_ (
    .a(_1125_),
    .b(_1124_),
    .c(_1126_)
  );
  or_bi _1991_ (
    .a(_1126_),
    .b(io_adder_out_31_),
    .c(_1127_)
  );
  or_ii _1992_ (
    .a(_1123_),
    .b(io_fn_1_),
    .c(_1128_)
  );
  or_bb _1993_ (
    .a(_1128_),
    .b(_1125_),
    .c(_1129_)
  );
  and_bi _1994_ (
    .a(_1128_),
    .b(_1124_),
    .c(_1130_)
  );
  and_bi _1995_ (
    .a(_1129_),
    .b(_1130_),
    .c(_1131_)
  );
  and_bi _1996_ (
    .a(_1127_),
    .b(_1131_),
    .c(_1132_)
  );
  or_bi _1997_ (
    .a(_1132_),
    .b(_1123_),
    .c(_1133_)
  );
  and_bi _1998_ (
    .a(io_fn_0_),
    .b(io_fn_1_),
    .c(_1134_)
  );
  and_bi _1999_ (
    .a(io_fn_2_),
    .b(io_fn_3_),
    .c(_1135_)
  );
  and_bb _2000_ (
    .a(_1135_),
    .b(_1134_),
    .c(_1136_)
  );
  and_bi _2001_ (
    .a(io_fn_3_),
    .b(io_fn_2_),
    .c(_1137_)
  );
  or_ii _2002_ (
    .a(io_fn_1_),
    .b(io_fn_0_),
    .c(_1138_)
  );
  and_bi _2003_ (
    .a(_1137_),
    .b(_1138_),
    .c(_1139_)
  );
  or_bb _2004_ (
    .a(_1139_),
    .b(_1136_),
    .c(_1140_)
  );
  inv _2005_ (
    .din(io_in2_4_),
    .dout(_1141_)
  );
  or_bb _2006_ (
    .a(_1140_),
    .b(_0737_),
    .c(_1142_)
  );
  and_bi _2007_ (
    .a(_1140_),
    .b(_0812_),
    .c(_1143_)
  );
  and_bi _2008_ (
    .a(_1142_),
    .b(_1143_),
    .c(_1144_)
  );
  or_bb _2009_ (
    .a(_1144_),
    .b(io_in2_0_),
    .c(_1145_)
  );
  or_bb _2010_ (
    .a(_1140_),
    .b(_0945_),
    .c(_1146_)
  );
  and_bi _2011_ (
    .a(_1140_),
    .b(_0821_),
    .c(_1147_)
  );
  and_bi _2012_ (
    .a(_1146_),
    .b(_1147_),
    .c(_1148_)
  );
  and_bi _2013_ (
    .a(io_in2_0_),
    .b(_1148_),
    .c(_1149_)
  );
  and_bi _2014_ (
    .a(_1145_),
    .b(_1149_),
    .c(_1150_)
  );
  or_bb _2015_ (
    .a(_1150_),
    .b(io_in2_1_),
    .c(_1151_)
  );
  or_bb _2016_ (
    .a(_1140_),
    .b(_0934_),
    .c(_1152_)
  );
  and_bi _2017_ (
    .a(_1140_),
    .b(_0832_),
    .c(_1153_)
  );
  and_bi _2018_ (
    .a(_1152_),
    .b(_1153_),
    .c(_1154_)
  );
  or_bb _2019_ (
    .a(_1154_),
    .b(io_in2_0_),
    .c(_1155_)
  );
  or_bb _2020_ (
    .a(_1140_),
    .b(_0925_),
    .c(_1156_)
  );
  and_bi _2021_ (
    .a(_1140_),
    .b(_0740_),
    .c(_1157_)
  );
  and_bi _2022_ (
    .a(_1156_),
    .b(_1157_),
    .c(_1158_)
  );
  and_bi _2023_ (
    .a(io_in2_0_),
    .b(_1158_),
    .c(_1159_)
  );
  and_bi _2024_ (
    .a(_1155_),
    .b(_1159_),
    .c(_1160_)
  );
  and_bi _2025_ (
    .a(io_in2_1_),
    .b(_1160_),
    .c(_1161_)
  );
  and_bi _2026_ (
    .a(_1151_),
    .b(_1161_),
    .c(_1162_)
  );
  and_bi _2027_ (
    .a(_0383_),
    .b(_1162_),
    .c(_1163_)
  );
  or_bb _2028_ (
    .a(_1140_),
    .b(_0914_),
    .c(_1164_)
  );
  and_bi _2029_ (
    .a(_1140_),
    .b(_0850_),
    .c(_1165_)
  );
  and_bi _2030_ (
    .a(_1164_),
    .b(_1165_),
    .c(_1166_)
  );
  or_bb _2031_ (
    .a(_1166_),
    .b(io_in2_0_),
    .c(_1167_)
  );
  inv _2032_ (
    .din(io_in1_18_),
    .dout(_1168_)
  );
  or_bb _2033_ (
    .a(_1140_),
    .b(_1168_),
    .c(_1169_)
  );
  and_bi _2034_ (
    .a(_1140_),
    .b(_0739_),
    .c(_1170_)
  );
  and_bi _2035_ (
    .a(_1169_),
    .b(_1170_),
    .c(_1171_)
  );
  and_bi _2036_ (
    .a(io_in2_0_),
    .b(_1171_),
    .c(_1172_)
  );
  and_bi _2037_ (
    .a(_1167_),
    .b(_1172_),
    .c(_1173_)
  );
  or_bb _2038_ (
    .a(_1173_),
    .b(io_in2_1_),
    .c(_1174_)
  );
  or_bb _2039_ (
    .a(_1140_),
    .b(_0738_),
    .c(_1175_)
  );
  and_bi _2040_ (
    .a(_1140_),
    .b(_0868_),
    .c(_1176_)
  );
  and_bi _2041_ (
    .a(_1175_),
    .b(_1176_),
    .c(_1177_)
  );
  or_bb _2042_ (
    .a(_1177_),
    .b(io_in2_0_),
    .c(_1178_)
  );
  inv _2043_ (
    .din(io_in2_0_),
    .dout(_1179_)
  );
  and_bi _2044_ (
    .a(io_in1_16_),
    .b(_1140_),
    .c(_1180_)
  );
  and_bi _2045_ (
    .a(_1140_),
    .b(_0877_),
    .c(_1181_)
  );
  or_bb _2046_ (
    .a(_1181_),
    .b(_1180_),
    .c(_1182_)
  );
  and_bi _2047_ (
    .a(_1182_),
    .b(_1179_),
    .c(_1183_)
  );
  and_bi _2048_ (
    .a(_1178_),
    .b(_1183_),
    .c(_1184_)
  );
  and_bi _2049_ (
    .a(io_in2_1_),
    .b(_1184_),
    .c(_1185_)
  );
  and_bi _2050_ (
    .a(_1174_),
    .b(_1185_),
    .c(_1186_)
  );
  and_bi _2051_ (
    .a(io_in2_2_),
    .b(_1186_),
    .c(_1187_)
  );
  or_bb _2052_ (
    .a(_1187_),
    .b(_1163_),
    .c(_1188_)
  );
  or_ii _2053_ (
    .a(_1188_),
    .b(io_in2_3_),
    .c(_1189_)
  );
  inv _2054_ (
    .din(io_in2_1_),
    .dout(_1190_)
  );
  or_bb _2055_ (
    .a(_1140_),
    .b(_0734_),
    .c(_1191_)
  );
  and_bi _2056_ (
    .a(_1140_),
    .b(_0773_),
    .c(_1192_)
  );
  and_bi _2057_ (
    .a(_1191_),
    .b(_1192_),
    .c(_1193_)
  );
  or_bb _2058_ (
    .a(_1193_),
    .b(io_in2_0_),
    .c(_1194_)
  );
  or_bb _2059_ (
    .a(_1140_),
    .b(_0735_),
    .c(_1195_)
  );
  and_bi _2060_ (
    .a(_1140_),
    .b(_0782_),
    .c(_1196_)
  );
  and_bi _2061_ (
    .a(_1195_),
    .b(_1196_),
    .c(_1197_)
  );
  and_bi _2062_ (
    .a(io_in2_0_),
    .b(_1197_),
    .c(_1198_)
  );
  and_bi _2063_ (
    .a(_1194_),
    .b(_1198_),
    .c(_1199_)
  );
  and_bi _2064_ (
    .a(_1190_),
    .b(_1199_),
    .c(_1200_)
  );
  or_bb _2065_ (
    .a(_1140_),
    .b(_0736_),
    .c(_1201_)
  );
  and_bi _2066_ (
    .a(_1140_),
    .b(_0793_),
    .c(_1202_)
  );
  and_bi _2067_ (
    .a(_1201_),
    .b(_1202_),
    .c(_1203_)
  );
  or_bb _2068_ (
    .a(_1203_),
    .b(io_in2_0_),
    .c(_1204_)
  );
  or_bb _2069_ (
    .a(_1140_),
    .b(_0964_),
    .c(_1205_)
  );
  and_bi _2070_ (
    .a(_1140_),
    .b(_0741_),
    .c(_1206_)
  );
  and_bi _2071_ (
    .a(_1205_),
    .b(_1206_),
    .c(_1207_)
  );
  and_bi _2072_ (
    .a(io_in2_0_),
    .b(_1207_),
    .c(_1208_)
  );
  and_bi _2073_ (
    .a(_1204_),
    .b(_1208_),
    .c(_1209_)
  );
  and_bi _2074_ (
    .a(io_in2_1_),
    .b(_1209_),
    .c(_1210_)
  );
  or_bb _2075_ (
    .a(_1210_),
    .b(_1200_),
    .c(_1211_)
  );
  and_bi _2076_ (
    .a(io_in2_2_),
    .b(_1211_),
    .c(_1212_)
  );
  and_bi _2077_ (
    .a(io_in1_29_),
    .b(_1140_),
    .c(_1213_)
  );
  and_bi _2078_ (
    .a(_1140_),
    .b(_0754_),
    .c(_1214_)
  );
  or_bb _2079_ (
    .a(_1214_),
    .b(_1213_),
    .c(_1215_)
  );
  or_ii _2080_ (
    .a(_1215_),
    .b(_1179_),
    .c(_1216_)
  );
  inv _2081_ (
    .din(io_in1_28_),
    .dout(_1217_)
  );
  or_bb _2082_ (
    .a(_1140_),
    .b(_1217_),
    .c(_1218_)
  );
  and_bi _2083_ (
    .a(_1140_),
    .b(_0762_),
    .c(_1219_)
  );
  and_bi _2084_ (
    .a(_1218_),
    .b(_1219_),
    .c(_1220_)
  );
  and_bi _2085_ (
    .a(io_in2_0_),
    .b(_1220_),
    .c(_1221_)
  );
  and_bi _2086_ (
    .a(_1216_),
    .b(_1221_),
    .c(_1222_)
  );
  or_bb _2087_ (
    .a(_1222_),
    .b(_1190_),
    .c(_1223_)
  );
  and_bi _2088_ (
    .a(io_in2_0_),
    .b(io_in2_1_),
    .c(_1224_)
  );
  or_bb _2089_ (
    .a(_1140_),
    .b(_0733_),
    .c(_1225_)
  );
  and_bi _2090_ (
    .a(_1140_),
    .b(_0742_),
    .c(_1226_)
  );
  and_bi _2091_ (
    .a(_1225_),
    .b(_1226_),
    .c(_1227_)
  );
  and_bi _2092_ (
    .a(_1224_),
    .b(_1227_),
    .c(_1228_)
  );
  and_bi _2093_ (
    .a(_1223_),
    .b(_1228_),
    .c(_1229_)
  );
  or_ii _2094_ (
    .a(_1140_),
    .b(_1112_),
    .c(_1230_)
  );
  and_bi _2095_ (
    .a(_0340_),
    .b(_1140_),
    .c(_1231_)
  );
  or_bb _2096_ (
    .a(_1231_),
    .b(_0384_),
    .c(_1232_)
  );
  and_bi _2097_ (
    .a(_1230_),
    .b(_1232_),
    .c(_1233_)
  );
  or_bb _2098_ (
    .a(_1233_),
    .b(io_in2_2_),
    .c(_1234_)
  );
  and_bi _2099_ (
    .a(_1229_),
    .b(_1234_),
    .c(_1235_)
  );
  or_bb _2100_ (
    .a(_1235_),
    .b(_1212_),
    .c(_1236_)
  );
  and_bi _2101_ (
    .a(_0764_),
    .b(_1236_),
    .c(_1237_)
  );
  and_bi _2102_ (
    .a(_1189_),
    .b(_1237_),
    .c(_1238_)
  );
  and_bi _2103_ (
    .a(_1141_),
    .b(_1238_),
    .c(_1239_)
  );
  and_bi _2104_ (
    .a(io_in1_15_),
    .b(_1140_),
    .c(_1240_)
  );
  and_bi _2105_ (
    .a(_1140_),
    .b(_0888_),
    .c(_1241_)
  );
  or_bb _2106_ (
    .a(_1241_),
    .b(_1240_),
    .c(_1242_)
  );
  or_ii _2107_ (
    .a(_1242_),
    .b(_1179_),
    .c(_1243_)
  );
  or_bb _2108_ (
    .a(_1140_),
    .b(_0868_),
    .c(_1244_)
  );
  and_bi _2109_ (
    .a(_1140_),
    .b(_0738_),
    .c(_1245_)
  );
  and_bi _2110_ (
    .a(_1244_),
    .b(_1245_),
    .c(_1246_)
  );
  and_bi _2111_ (
    .a(io_in2_0_),
    .b(_1246_),
    .c(_1247_)
  );
  and_bi _2112_ (
    .a(_1243_),
    .b(_1247_),
    .c(_1248_)
  );
  or_bb _2113_ (
    .a(_1248_),
    .b(io_in2_1_),
    .c(_1249_)
  );
  or_bb _2114_ (
    .a(_1140_),
    .b(_0739_),
    .c(_1250_)
  );
  and_bi _2115_ (
    .a(_1140_),
    .b(_1168_),
    .c(_1251_)
  );
  and_bi _2116_ (
    .a(_1250_),
    .b(_1251_),
    .c(_1252_)
  );
  or_bb _2117_ (
    .a(_1252_),
    .b(io_in2_0_),
    .c(_1253_)
  );
  or_bb _2118_ (
    .a(_1140_),
    .b(_0850_),
    .c(_1254_)
  );
  and_bi _2119_ (
    .a(_1140_),
    .b(_0914_),
    .c(_1255_)
  );
  and_bi _2120_ (
    .a(_1254_),
    .b(_1255_),
    .c(_1256_)
  );
  and_bi _2121_ (
    .a(io_in2_0_),
    .b(_1256_),
    .c(_1257_)
  );
  and_bi _2122_ (
    .a(_1253_),
    .b(_1257_),
    .c(_1258_)
  );
  and_bi _2123_ (
    .a(io_in2_1_),
    .b(_1258_),
    .c(_1259_)
  );
  and_bi _2124_ (
    .a(_1249_),
    .b(_1259_),
    .c(_1260_)
  );
  and_bi _2125_ (
    .a(_0383_),
    .b(_1260_),
    .c(_1261_)
  );
  or_bb _2126_ (
    .a(_1140_),
    .b(_0740_),
    .c(_1262_)
  );
  and_bi _2127_ (
    .a(_1140_),
    .b(_0925_),
    .c(_1263_)
  );
  and_bi _2128_ (
    .a(_1262_),
    .b(_1263_),
    .c(_1264_)
  );
  or_bb _2129_ (
    .a(_1264_),
    .b(io_in2_0_),
    .c(_1265_)
  );
  or_bb _2130_ (
    .a(_1140_),
    .b(_0832_),
    .c(_1266_)
  );
  and_bi _2131_ (
    .a(_1140_),
    .b(_0934_),
    .c(_1267_)
  );
  and_bi _2132_ (
    .a(_1266_),
    .b(_1267_),
    .c(_1268_)
  );
  and_bi _2133_ (
    .a(io_in2_0_),
    .b(_1268_),
    .c(_1269_)
  );
  and_bi _2134_ (
    .a(_1265_),
    .b(_1269_),
    .c(_1270_)
  );
  or_bb _2135_ (
    .a(_1270_),
    .b(io_in2_1_),
    .c(_1271_)
  );
  or_bb _2136_ (
    .a(_1140_),
    .b(_0821_),
    .c(_1272_)
  );
  and_bi _2137_ (
    .a(_1140_),
    .b(_0945_),
    .c(_1273_)
  );
  and_bi _2138_ (
    .a(_1272_),
    .b(_1273_),
    .c(_1274_)
  );
  or_bb _2139_ (
    .a(_1274_),
    .b(io_in2_0_),
    .c(_1275_)
  );
  or_bb _2140_ (
    .a(_1140_),
    .b(_0812_),
    .c(_1276_)
  );
  and_bi _2141_ (
    .a(_1140_),
    .b(_0737_),
    .c(_1277_)
  );
  and_bi _2142_ (
    .a(_1276_),
    .b(_1277_),
    .c(_1278_)
  );
  and_bi _2143_ (
    .a(io_in2_0_),
    .b(_1278_),
    .c(_1279_)
  );
  and_bi _2144_ (
    .a(_1275_),
    .b(_1279_),
    .c(_1280_)
  );
  and_bi _2145_ (
    .a(io_in2_1_),
    .b(_1280_),
    .c(_1281_)
  );
  and_bi _2146_ (
    .a(_1271_),
    .b(_1281_),
    .c(_1282_)
  );
  and_bi _2147_ (
    .a(io_in2_2_),
    .b(_1282_),
    .c(_1283_)
  );
  or_bb _2148_ (
    .a(_1283_),
    .b(_1261_),
    .c(_1284_)
  );
  or_ii _2149_ (
    .a(_1284_),
    .b(_0764_),
    .c(_1285_)
  );
  or_bb _2150_ (
    .a(_1140_),
    .b(_0741_),
    .c(_1286_)
  );
  and_bi _2151_ (
    .a(_1140_),
    .b(_0964_),
    .c(_1287_)
  );
  and_bi _2152_ (
    .a(_1286_),
    .b(_1287_),
    .c(_1288_)
  );
  or_bb _2153_ (
    .a(_1288_),
    .b(io_in2_0_),
    .c(_1289_)
  );
  or_bb _2154_ (
    .a(_1140_),
    .b(_0793_),
    .c(_1290_)
  );
  and_bi _2155_ (
    .a(_1140_),
    .b(_0736_),
    .c(_1291_)
  );
  and_bi _2156_ (
    .a(_1290_),
    .b(_1291_),
    .c(_1292_)
  );
  and_bi _2157_ (
    .a(io_in2_0_),
    .b(_1292_),
    .c(_1293_)
  );
  and_bi _2158_ (
    .a(_1289_),
    .b(_1293_),
    .c(_1294_)
  );
  or_bb _2159_ (
    .a(_1294_),
    .b(io_in2_1_),
    .c(_1295_)
  );
  or_bb _2160_ (
    .a(_1140_),
    .b(_0782_),
    .c(_1296_)
  );
  and_bi _2161_ (
    .a(_1140_),
    .b(_0735_),
    .c(_1297_)
  );
  and_bi _2162_ (
    .a(_1296_),
    .b(_1297_),
    .c(_1298_)
  );
  or_bb _2163_ (
    .a(_1298_),
    .b(io_in2_0_),
    .c(_1299_)
  );
  or_bb _2164_ (
    .a(_1140_),
    .b(_0773_),
    .c(_1300_)
  );
  and_bi _2165_ (
    .a(_1140_),
    .b(_0734_),
    .c(_1301_)
  );
  and_bi _2166_ (
    .a(_1300_),
    .b(_1301_),
    .c(_1302_)
  );
  and_bi _2167_ (
    .a(io_in2_0_),
    .b(_1302_),
    .c(_1303_)
  );
  and_bi _2168_ (
    .a(_1299_),
    .b(_1303_),
    .c(_1304_)
  );
  and_bi _2169_ (
    .a(io_in2_1_),
    .b(_1304_),
    .c(_1305_)
  );
  and_bi _2170_ (
    .a(_1295_),
    .b(_1305_),
    .c(_1306_)
  );
  or_bb _2171_ (
    .a(_1306_),
    .b(io_in2_2_),
    .c(_1307_)
  );
  or_bb _2172_ (
    .a(_1140_),
    .b(_0762_),
    .c(_1308_)
  );
  and_bi _2173_ (
    .a(_1140_),
    .b(_1217_),
    .c(_1309_)
  );
  and_bi _2174_ (
    .a(_1308_),
    .b(_1309_),
    .c(_1310_)
  );
  or_bb _2175_ (
    .a(_1310_),
    .b(io_in2_0_),
    .c(_1311_)
  );
  or_bb _2176_ (
    .a(_1140_),
    .b(_0754_),
    .c(_1312_)
  );
  and_bi _2177_ (
    .a(_1140_),
    .b(_1004_),
    .c(_1313_)
  );
  and_bi _2178_ (
    .a(_1312_),
    .b(_1313_),
    .c(_1314_)
  );
  and_bi _2179_ (
    .a(io_in2_0_),
    .b(_1314_),
    .c(_1315_)
  );
  and_bi _2180_ (
    .a(_1311_),
    .b(_1315_),
    .c(_1316_)
  );
  or_bb _2181_ (
    .a(_1316_),
    .b(io_in2_1_),
    .c(_1317_)
  );
  or_bb _2182_ (
    .a(_1140_),
    .b(_0742_),
    .c(_1318_)
  );
  and_bi _2183_ (
    .a(_1140_),
    .b(_0733_),
    .c(_1319_)
  );
  and_bi _2184_ (
    .a(_1318_),
    .b(_1319_),
    .c(_1320_)
  );
  and_bi _2185_ (
    .a(_1179_),
    .b(_1320_),
    .c(_1321_)
  );
  and_bi _2186_ (
    .a(io_in1_0_),
    .b(_1140_),
    .c(_1322_)
  );
  and_bi _2187_ (
    .a(_1140_),
    .b(_0340_),
    .c(_1323_)
  );
  or_bb _2188_ (
    .a(_1323_),
    .b(_1322_),
    .c(_1324_)
  );
  and_bi _2189_ (
    .a(_1324_),
    .b(_1179_),
    .c(_1325_)
  );
  or_bb _2190_ (
    .a(_1325_),
    .b(_1321_),
    .c(_1326_)
  );
  and_bi _2191_ (
    .a(_1326_),
    .b(_1190_),
    .c(_1327_)
  );
  and_bi _2192_ (
    .a(_1317_),
    .b(_1327_),
    .c(_1328_)
  );
  and_bi _2193_ (
    .a(io_in2_2_),
    .b(_1328_),
    .c(_1329_)
  );
  and_bi _2194_ (
    .a(_1307_),
    .b(_1329_),
    .c(_1330_)
  );
  and_bi _2195_ (
    .a(io_in2_3_),
    .b(_1330_),
    .c(_1331_)
  );
  and_bi _2196_ (
    .a(_1285_),
    .b(_1331_),
    .c(_1332_)
  );
  and_bi _2197_ (
    .a(io_in2_4_),
    .b(_1332_),
    .c(_1333_)
  );
  or_bb _2198_ (
    .a(_1333_),
    .b(_1239_),
    .c(_1334_)
  );
  or_bi _2199_ (
    .a(_1334_),
    .b(_1140_),
    .c(_1335_)
  );
  and_bi _2200_ (
    .a(_1134_),
    .b(_1118_),
    .c(_1336_)
  );
  inv _2201_ (
    .din(_1336_),
    .dout(_1337_)
  );
  and_bi _2202_ (
    .a(_0352_),
    .b(_0415_),
    .c(_1338_)
  );
  or_bi _2203_ (
    .a(_1338_),
    .b(_1324_),
    .c(_1339_)
  );
  or_bb _2204_ (
    .a(_1339_),
    .b(_1337_),
    .c(_1340_)
  );
  and_bi _2205_ (
    .a(_1135_),
    .b(_1119_),
    .c(_1341_)
  );
  and_bb _2206_ (
    .a(_1341_),
    .b(_0743_),
    .c(_1342_)
  );
  and_bi _2207_ (
    .a(_1135_),
    .b(io_fn_0_),
    .c(_1343_)
  );
  and_bi _2208_ (
    .a(_1112_),
    .b(_1343_),
    .c(_1344_)
  );
  and_bi _2209_ (
    .a(_1135_),
    .b(_1138_),
    .c(_1345_)
  );
  or_bb _2210_ (
    .a(_1345_),
    .b(_1113_),
    .c(_1346_)
  );
  or_bb _2211_ (
    .a(_1346_),
    .b(_1344_),
    .c(_1347_)
  );
  or_bb _2212_ (
    .a(_1347_),
    .b(_1342_),
    .c(_1348_)
  );
  and_bi _2213_ (
    .a(_1345_),
    .b(_1111_),
    .c(_1349_)
  );
  and_bi _2214_ (
    .a(_1348_),
    .b(_1349_),
    .c(_1350_)
  );
  and_bi _2215_ (
    .a(_1337_),
    .b(_1350_),
    .c(_1351_)
  );
  or_bb _2216_ (
    .a(_1351_),
    .b(_1140_),
    .c(_1352_)
  );
  and_bi _2217_ (
    .a(_1340_),
    .b(_1352_),
    .c(_1353_)
  );
  or_bb _2218_ (
    .a(_1353_),
    .b(_1123_),
    .c(_1354_)
  );
  and_bi _2219_ (
    .a(_1335_),
    .b(_1354_),
    .c(_1355_)
  );
  or_bi _2220_ (
    .a(_1355_),
    .b(_1121_),
    .c(_1356_)
  );
  and_bi _2221_ (
    .a(_1133_),
    .b(_1356_),
    .c(_1357_)
  );
  and_bi _2222_ (
    .a(_1122_),
    .b(_1357_),
    .c(io_out_0_)
  );
  and_bi _2223_ (
    .a(io_adder_out_1_),
    .b(_1121_),
    .c(_1358_)
  );
  or_ii _2224_ (
    .a(_1324_),
    .b(io_fn_3_),
    .c(_1359_)
  );
  and_bi _2225_ (
    .a(io_in2_4_),
    .b(_1359_),
    .c(_1360_)
  );
  inv _2226_ (
    .din(_1360_),
    .dout(_1361_)
  );
  or_bb _2227_ (
    .a(_1359_),
    .b(_0764_),
    .c(_1362_)
  );
  and_bi _2228_ (
    .a(io_in2_2_),
    .b(_1359_),
    .c(_1363_)
  );
  inv _2229_ (
    .din(_1363_),
    .dout(_1364_)
  );
  and_bi _2230_ (
    .a(_1359_),
    .b(_1190_),
    .c(_1365_)
  );
  and_bi _2231_ (
    .a(_1190_),
    .b(_1326_),
    .c(_1366_)
  );
  or_bb _2232_ (
    .a(_1366_),
    .b(_1365_),
    .c(_1367_)
  );
  and_bi _2233_ (
    .a(_0383_),
    .b(_1367_),
    .c(_1368_)
  );
  and_bi _2234_ (
    .a(_1364_),
    .b(_1368_),
    .c(_1369_)
  );
  and_bi _2235_ (
    .a(_0764_),
    .b(_1369_),
    .c(_1370_)
  );
  and_bi _2236_ (
    .a(_1362_),
    .b(_1370_),
    .c(_1371_)
  );
  and_bi _2237_ (
    .a(_1141_),
    .b(_1371_),
    .c(_1372_)
  );
  and_bi _2238_ (
    .a(_1361_),
    .b(_1372_),
    .c(_1373_)
  );
  and_bi _2239_ (
    .a(_1336_),
    .b(_1373_),
    .c(_1374_)
  );
  and_bi _2240_ (
    .a(_1343_),
    .b(_1190_),
    .c(_1375_)
  );
  or_bb _2241_ (
    .a(_1375_),
    .b(io_in1_1_),
    .c(_1376_)
  );
  and_bb _2242_ (
    .a(io_in2_1_),
    .b(io_in1_1_),
    .c(_1377_)
  );
  and_bb _2243_ (
    .a(_1377_),
    .b(_1341_),
    .c(_1378_)
  );
  and_bi _2244_ (
    .a(_1376_),
    .b(_1378_),
    .c(_1379_)
  );
  or_bb _2245_ (
    .a(_1379_),
    .b(_1345_),
    .c(_1380_)
  );
  and_bi _2246_ (
    .a(_1345_),
    .b(_1377_),
    .c(_1381_)
  );
  or_bb _2247_ (
    .a(_1381_),
    .b(_1336_),
    .c(_1382_)
  );
  and_bi _2248_ (
    .a(_1380_),
    .b(_1382_),
    .c(_1383_)
  );
  or_bb _2249_ (
    .a(_1383_),
    .b(_1140_),
    .c(_1384_)
  );
  or_bb _2250_ (
    .a(_1384_),
    .b(_1374_),
    .c(_1385_)
  );
  or_bb _2251_ (
    .a(_1148_),
    .b(io_in2_0_),
    .c(_1386_)
  );
  and_bi _2252_ (
    .a(io_in2_0_),
    .b(_1154_),
    .c(_1387_)
  );
  and_bi _2253_ (
    .a(_1386_),
    .b(_1387_),
    .c(_1388_)
  );
  and_bi _2254_ (
    .a(_1190_),
    .b(_1388_),
    .c(_1389_)
  );
  or_bb _2255_ (
    .a(_1158_),
    .b(io_in2_0_),
    .c(_1390_)
  );
  and_bi _2256_ (
    .a(io_in2_0_),
    .b(_1166_),
    .c(_1391_)
  );
  and_bi _2257_ (
    .a(_1390_),
    .b(_1391_),
    .c(_1392_)
  );
  and_bi _2258_ (
    .a(io_in2_1_),
    .b(_1392_),
    .c(_1393_)
  );
  or_bb _2259_ (
    .a(_1393_),
    .b(_1389_),
    .c(_1394_)
  );
  or_ii _2260_ (
    .a(_1394_),
    .b(_0383_),
    .c(_1395_)
  );
  or_bb _2261_ (
    .a(_1171_),
    .b(io_in2_0_),
    .c(_1396_)
  );
  and_bi _2262_ (
    .a(io_in2_0_),
    .b(_1177_),
    .c(_1397_)
  );
  and_bi _2263_ (
    .a(_1396_),
    .b(_1397_),
    .c(_1398_)
  );
  or_bb _2264_ (
    .a(_1398_),
    .b(io_in2_1_),
    .c(_1399_)
  );
  and_bi _2265_ (
    .a(io_in2_0_),
    .b(_1242_),
    .c(_1400_)
  );
  and_bi _2266_ (
    .a(_1179_),
    .b(_1182_),
    .c(_1401_)
  );
  or_bb _2267_ (
    .a(_1401_),
    .b(_1400_),
    .c(_1402_)
  );
  and_bi _2268_ (
    .a(io_in2_1_),
    .b(_1402_),
    .c(_1403_)
  );
  and_bi _2269_ (
    .a(_1399_),
    .b(_1403_),
    .c(_1404_)
  );
  and_bi _2270_ (
    .a(io_in2_2_),
    .b(_1404_),
    .c(_1405_)
  );
  and_bi _2271_ (
    .a(_1395_),
    .b(_1405_),
    .c(_1406_)
  );
  or_bb _2272_ (
    .a(_1406_),
    .b(_0764_),
    .c(_1407_)
  );
  or_bb _2273_ (
    .a(_1220_),
    .b(io_in2_0_),
    .c(_1408_)
  );
  and_bi _2274_ (
    .a(io_in2_0_),
    .b(_1193_),
    .c(_1409_)
  );
  and_bi _2275_ (
    .a(_1408_),
    .b(_1409_),
    .c(_1410_)
  );
  or_bb _2276_ (
    .a(_1410_),
    .b(_1190_),
    .c(_1411_)
  );
  and_bb _2277_ (
    .a(_1224_),
    .b(_1215_),
    .c(_1412_)
  );
  or_bb _2278_ (
    .a(_1227_),
    .b(_0384_),
    .c(_1413_)
  );
  or_ii _2279_ (
    .a(_1413_),
    .b(_0383_),
    .c(_1414_)
  );
  or_bb _2280_ (
    .a(_1414_),
    .b(_1412_),
    .c(_1415_)
  );
  and_bi _2281_ (
    .a(_1411_),
    .b(_1415_),
    .c(_1416_)
  );
  or_bb _2282_ (
    .a(_1197_),
    .b(io_in2_0_),
    .c(_1417_)
  );
  and_bi _2283_ (
    .a(io_in2_0_),
    .b(_1203_),
    .c(_1418_)
  );
  and_bi _2284_ (
    .a(_1417_),
    .b(_1418_),
    .c(_1419_)
  );
  and_bi _2285_ (
    .a(_1190_),
    .b(_1419_),
    .c(_1420_)
  );
  or_bb _2286_ (
    .a(_1207_),
    .b(io_in2_0_),
    .c(_1421_)
  );
  and_bi _2287_ (
    .a(io_in2_0_),
    .b(_1144_),
    .c(_1422_)
  );
  and_bi _2288_ (
    .a(_1421_),
    .b(_1422_),
    .c(_1423_)
  );
  and_bi _2289_ (
    .a(io_in2_1_),
    .b(_1423_),
    .c(_1424_)
  );
  or_bb _2290_ (
    .a(_1424_),
    .b(_1420_),
    .c(_1425_)
  );
  and_bi _2291_ (
    .a(io_in2_2_),
    .b(_1425_),
    .c(_1426_)
  );
  or_bb _2292_ (
    .a(_1426_),
    .b(_1416_),
    .c(_1427_)
  );
  and_bi _2293_ (
    .a(_0764_),
    .b(_1427_),
    .c(_1428_)
  );
  and_bi _2294_ (
    .a(_1407_),
    .b(_1428_),
    .c(_1429_)
  );
  and_bi _2295_ (
    .a(_1141_),
    .b(_1429_),
    .c(_1430_)
  );
  or_bb _2296_ (
    .a(_1246_),
    .b(io_in2_0_),
    .c(_1431_)
  );
  and_bi _2297_ (
    .a(io_in2_0_),
    .b(_1252_),
    .c(_1432_)
  );
  and_bi _2298_ (
    .a(_1431_),
    .b(_1432_),
    .c(_1433_)
  );
  or_bb _2299_ (
    .a(_1433_),
    .b(io_in2_1_),
    .c(_1434_)
  );
  or_bb _2300_ (
    .a(_1256_),
    .b(io_in2_0_),
    .c(_1435_)
  );
  and_bi _2301_ (
    .a(io_in2_0_),
    .b(_1264_),
    .c(_1436_)
  );
  and_bi _2302_ (
    .a(_1435_),
    .b(_1436_),
    .c(_1437_)
  );
  and_bi _2303_ (
    .a(io_in2_1_),
    .b(_1437_),
    .c(_1438_)
  );
  and_bi _2304_ (
    .a(_1434_),
    .b(_1438_),
    .c(_1439_)
  );
  or_bb _2305_ (
    .a(_1439_),
    .b(io_in2_2_),
    .c(_1440_)
  );
  or_bb _2306_ (
    .a(_1268_),
    .b(io_in2_0_),
    .c(_1441_)
  );
  and_bi _2307_ (
    .a(io_in2_0_),
    .b(_1274_),
    .c(_1442_)
  );
  and_bi _2308_ (
    .a(_1441_),
    .b(_1442_),
    .c(_1443_)
  );
  or_bb _2309_ (
    .a(_1443_),
    .b(io_in2_1_),
    .c(_1444_)
  );
  or_bb _2310_ (
    .a(_1278_),
    .b(io_in2_0_),
    .c(_1445_)
  );
  and_bi _2311_ (
    .a(io_in2_0_),
    .b(_1288_),
    .c(_1446_)
  );
  and_bi _2312_ (
    .a(_1445_),
    .b(_1446_),
    .c(_1447_)
  );
  and_bi _2313_ (
    .a(io_in2_1_),
    .b(_1447_),
    .c(_1448_)
  );
  and_bi _2314_ (
    .a(_1444_),
    .b(_1448_),
    .c(_1449_)
  );
  and_bi _2315_ (
    .a(io_in2_2_),
    .b(_1449_),
    .c(_1450_)
  );
  and_bi _2316_ (
    .a(_1440_),
    .b(_1450_),
    .c(_1451_)
  );
  or_bb _2317_ (
    .a(_1451_),
    .b(io_in2_3_),
    .c(_1452_)
  );
  or_bb _2318_ (
    .a(_1292_),
    .b(io_in2_0_),
    .c(_1453_)
  );
  and_bi _2319_ (
    .a(io_in2_0_),
    .b(_1298_),
    .c(_1454_)
  );
  and_bi _2320_ (
    .a(_1453_),
    .b(_1454_),
    .c(_1455_)
  );
  or_bb _2321_ (
    .a(_1455_),
    .b(io_in2_1_),
    .c(_1456_)
  );
  or_bb _2322_ (
    .a(_1302_),
    .b(io_in2_0_),
    .c(_1457_)
  );
  and_bi _2323_ (
    .a(io_in2_0_),
    .b(_1310_),
    .c(_1458_)
  );
  and_bi _2324_ (
    .a(_1457_),
    .b(_1458_),
    .c(_1459_)
  );
  and_bi _2325_ (
    .a(io_in2_1_),
    .b(_1459_),
    .c(_1460_)
  );
  and_bi _2326_ (
    .a(_1456_),
    .b(_1460_),
    .c(_1461_)
  );
  or_bb _2327_ (
    .a(_1461_),
    .b(io_in2_2_),
    .c(_1462_)
  );
  and_bi _2328_ (
    .a(_1324_),
    .b(io_in2_0_),
    .c(_1463_)
  );
  and_bi _2329_ (
    .a(_1365_),
    .b(_1463_),
    .c(_1464_)
  );
  and_bi _2330_ (
    .a(_1179_),
    .b(_1314_),
    .c(_1465_)
  );
  and_bi _2331_ (
    .a(io_in2_0_),
    .b(_1320_),
    .c(_1466_)
  );
  or_bb _2332_ (
    .a(_1466_),
    .b(_1465_),
    .c(_1467_)
  );
  and_bi _2333_ (
    .a(_1190_),
    .b(_1467_),
    .c(_1468_)
  );
  or_bb _2334_ (
    .a(_1468_),
    .b(_1464_),
    .c(_1469_)
  );
  and_bi _2335_ (
    .a(io_in2_2_),
    .b(_1469_),
    .c(_1470_)
  );
  and_bi _2336_ (
    .a(_1462_),
    .b(_1470_),
    .c(_1471_)
  );
  and_bi _2337_ (
    .a(io_in2_3_),
    .b(_1471_),
    .c(_1472_)
  );
  and_bi _2338_ (
    .a(_1452_),
    .b(_1472_),
    .c(_1473_)
  );
  and_bi _2339_ (
    .a(io_in2_4_),
    .b(_1473_),
    .c(_1474_)
  );
  or_bb _2340_ (
    .a(_1474_),
    .b(_1430_),
    .c(_1475_)
  );
  and_bi _2341_ (
    .a(_1140_),
    .b(_1475_),
    .c(_1476_)
  );
  or_bi _2342_ (
    .a(_1123_),
    .b(_1121_),
    .c(_1477_)
  );
  or_bb _2343_ (
    .a(_1477_),
    .b(_1476_),
    .c(_1478_)
  );
  and_bi _2344_ (
    .a(_1385_),
    .b(_1478_),
    .c(_1479_)
  );
  or_bb _2345_ (
    .a(_1479_),
    .b(_1358_),
    .c(io_out_1_)
  );
  and_bi _2346_ (
    .a(io_adder_out_2_),
    .b(_1121_),
    .c(_1480_)
  );
  and_bi _2347_ (
    .a(_0383_),
    .b(_1469_),
    .c(_1481_)
  );
  and_bi _2348_ (
    .a(_1364_),
    .b(_1481_),
    .c(_1482_)
  );
  and_bi _2349_ (
    .a(_0764_),
    .b(_1482_),
    .c(_1483_)
  );
  and_bi _2350_ (
    .a(_1362_),
    .b(_1483_),
    .c(_1484_)
  );
  and_bi _2351_ (
    .a(_1141_),
    .b(_1484_),
    .c(_1485_)
  );
  and_bi _2352_ (
    .a(_1361_),
    .b(_1485_),
    .c(_1486_)
  );
  and_bi _2353_ (
    .a(_1336_),
    .b(_1486_),
    .c(_1487_)
  );
  and_bi _2354_ (
    .a(_1343_),
    .b(_0383_),
    .c(_1488_)
  );
  or_bb _2355_ (
    .a(_1488_),
    .b(io_in1_2_),
    .c(_1489_)
  );
  and_bb _2356_ (
    .a(io_in2_2_),
    .b(io_in1_2_),
    .c(_1490_)
  );
  and_bb _2357_ (
    .a(_1490_),
    .b(_1341_),
    .c(_1491_)
  );
  and_bi _2358_ (
    .a(_1489_),
    .b(_1491_),
    .c(_1492_)
  );
  or_bb _2359_ (
    .a(_1492_),
    .b(_1345_),
    .c(_1493_)
  );
  and_bi _2360_ (
    .a(_1345_),
    .b(_1490_),
    .c(_1494_)
  );
  or_bb _2361_ (
    .a(_1494_),
    .b(_1336_),
    .c(_1495_)
  );
  and_bi _2362_ (
    .a(_1493_),
    .b(_1495_),
    .c(_1496_)
  );
  or_bb _2363_ (
    .a(_1496_),
    .b(_1140_),
    .c(_1497_)
  );
  or_bb _2364_ (
    .a(_1497_),
    .b(_1487_),
    .c(_1498_)
  );
  or_bb _2365_ (
    .a(_1222_),
    .b(io_in2_1_),
    .c(_1499_)
  );
  and_bi _2366_ (
    .a(io_in2_1_),
    .b(_1199_),
    .c(_1500_)
  );
  or_bb _2367_ (
    .a(_1500_),
    .b(io_in2_2_),
    .c(_1501_)
  );
  and_bi _2368_ (
    .a(_1499_),
    .b(_1501_),
    .c(_1502_)
  );
  and_bi _2369_ (
    .a(_1190_),
    .b(_1209_),
    .c(_1503_)
  );
  and_bi _2370_ (
    .a(io_in2_1_),
    .b(_1150_),
    .c(_1504_)
  );
  or_bb _2371_ (
    .a(_1504_),
    .b(_1503_),
    .c(_1505_)
  );
  and_bi _2372_ (
    .a(io_in2_2_),
    .b(_1505_),
    .c(_1506_)
  );
  or_bb _2373_ (
    .a(_1506_),
    .b(_1502_),
    .c(_1507_)
  );
  and_bi _2374_ (
    .a(_0764_),
    .b(_1507_),
    .c(_1508_)
  );
  and_bi _2375_ (
    .a(_1190_),
    .b(_1160_),
    .c(_1509_)
  );
  and_bi _2376_ (
    .a(io_in2_1_),
    .b(_1173_),
    .c(_1510_)
  );
  or_bb _2377_ (
    .a(_1510_),
    .b(_1509_),
    .c(_1511_)
  );
  or_ii _2378_ (
    .a(_1511_),
    .b(_0383_),
    .c(_1512_)
  );
  or_bb _2379_ (
    .a(_1184_),
    .b(io_in2_1_),
    .c(_1513_)
  );
  and_bi _2380_ (
    .a(io_in2_1_),
    .b(_1248_),
    .c(_1514_)
  );
  and_bi _2381_ (
    .a(_1513_),
    .b(_1514_),
    .c(_1515_)
  );
  and_bi _2382_ (
    .a(io_in2_2_),
    .b(_1515_),
    .c(_1516_)
  );
  and_bi _2383_ (
    .a(_1512_),
    .b(_1516_),
    .c(_1517_)
  );
  and_bi _2384_ (
    .a(io_in2_3_),
    .b(_1517_),
    .c(_0000_)
  );
  or_bb _2385_ (
    .a(_0000_),
    .b(io_in2_4_),
    .c(_0001_)
  );
  or_bb _2386_ (
    .a(_0001_),
    .b(_1508_),
    .c(_0002_)
  );
  or_bb _2387_ (
    .a(_1258_),
    .b(io_in2_1_),
    .c(_0003_)
  );
  and_bi _2388_ (
    .a(io_in2_1_),
    .b(_1270_),
    .c(_0004_)
  );
  and_bi _2389_ (
    .a(_0003_),
    .b(_0004_),
    .c(_0005_)
  );
  or_bb _2390_ (
    .a(_0005_),
    .b(io_in2_2_),
    .c(_0006_)
  );
  or_bb _2391_ (
    .a(_1280_),
    .b(io_in2_1_),
    .c(_0007_)
  );
  and_bi _2392_ (
    .a(io_in2_1_),
    .b(_1294_),
    .c(_0008_)
  );
  and_bi _2393_ (
    .a(_0007_),
    .b(_0008_),
    .c(_0009_)
  );
  and_bi _2394_ (
    .a(io_in2_2_),
    .b(_0009_),
    .c(_0010_)
  );
  and_bi _2395_ (
    .a(_0006_),
    .b(_0010_),
    .c(_0011_)
  );
  and_bi _2396_ (
    .a(_0764_),
    .b(_0011_),
    .c(_0012_)
  );
  and_bi _2397_ (
    .a(_1367_),
    .b(_0383_),
    .c(_0013_)
  );
  and_bi _2398_ (
    .a(_1190_),
    .b(_1304_),
    .c(_0014_)
  );
  and_bi _2399_ (
    .a(io_in2_1_),
    .b(_1316_),
    .c(_0015_)
  );
  or_bb _2400_ (
    .a(_0015_),
    .b(_0014_),
    .c(_0016_)
  );
  and_bi _2401_ (
    .a(_0383_),
    .b(_0016_),
    .c(_0017_)
  );
  or_bb _2402_ (
    .a(_0017_),
    .b(_0013_),
    .c(_0018_)
  );
  and_bi _2403_ (
    .a(io_in2_3_),
    .b(_0018_),
    .c(_0019_)
  );
  or_bb _2404_ (
    .a(_0019_),
    .b(_0012_),
    .c(_0020_)
  );
  and_bi _2405_ (
    .a(io_in2_4_),
    .b(_0020_),
    .c(_0021_)
  );
  or_bi _2406_ (
    .a(_0021_),
    .b(_0002_),
    .c(_0022_)
  );
  and_bb _2407_ (
    .a(_0022_),
    .b(_1140_),
    .c(_0023_)
  );
  or_bb _2408_ (
    .a(_0023_),
    .b(_1477_),
    .c(_0024_)
  );
  and_bi _2409_ (
    .a(_1498_),
    .b(_0024_),
    .c(_0025_)
  );
  or_bb _2410_ (
    .a(_0025_),
    .b(_1480_),
    .c(io_out_2_)
  );
  and_bi _2411_ (
    .a(io_adder_out_3_),
    .b(_1121_),
    .c(_0026_)
  );
  and_bi _2412_ (
    .a(_0383_),
    .b(_1328_),
    .c(_0027_)
  );
  or_bb _2413_ (
    .a(_0027_),
    .b(_1363_),
    .c(_0028_)
  );
  and_bi _2414_ (
    .a(_0028_),
    .b(io_in2_3_),
    .c(_0029_)
  );
  and_bi _2415_ (
    .a(_1362_),
    .b(_0029_),
    .c(_0030_)
  );
  and_bi _2416_ (
    .a(_1141_),
    .b(_0030_),
    .c(_0031_)
  );
  and_bi _2417_ (
    .a(_1361_),
    .b(_0031_),
    .c(_0032_)
  );
  and_bi _2418_ (
    .a(_1336_),
    .b(_0032_),
    .c(_0033_)
  );
  or_ii _2419_ (
    .a(io_in2_3_),
    .b(io_in1_3_),
    .c(_0034_)
  );
  or_bi _2420_ (
    .a(_0034_),
    .b(_1345_),
    .c(_0035_)
  );
  and_bi _2421_ (
    .a(_1343_),
    .b(_0764_),
    .c(_0036_)
  );
  or_bb _2422_ (
    .a(_0036_),
    .b(io_in1_3_),
    .c(_0037_)
  );
  and_bi _2423_ (
    .a(_1341_),
    .b(_0034_),
    .c(_0038_)
  );
  or_bb _2424_ (
    .a(_0038_),
    .b(_1345_),
    .c(_0039_)
  );
  and_bi _2425_ (
    .a(_0037_),
    .b(_0039_),
    .c(_0040_)
  );
  and_bi _2426_ (
    .a(_0035_),
    .b(_0040_),
    .c(_0041_)
  );
  and_bi _2427_ (
    .a(_1337_),
    .b(_0041_),
    .c(_0042_)
  );
  or_bb _2428_ (
    .a(_0042_),
    .b(_1140_),
    .c(_0043_)
  );
  or_bb _2429_ (
    .a(_0043_),
    .b(_0033_),
    .c(_0044_)
  );
  or_bb _2430_ (
    .a(_1419_),
    .b(_1190_),
    .c(_0045_)
  );
  and_bi _2431_ (
    .a(_1190_),
    .b(_1410_),
    .c(_0046_)
  );
  and_bi _2432_ (
    .a(_0045_),
    .b(_0046_),
    .c(_0047_)
  );
  or_bb _2433_ (
    .a(_0047_),
    .b(io_in2_2_),
    .c(_0048_)
  );
  or_bb _2434_ (
    .a(_1423_),
    .b(io_in2_1_),
    .c(_0049_)
  );
  and_bi _2435_ (
    .a(io_in2_1_),
    .b(_1388_),
    .c(_0050_)
  );
  and_bi _2436_ (
    .a(_0049_),
    .b(_0050_),
    .c(_0051_)
  );
  and_bi _2437_ (
    .a(io_in2_2_),
    .b(_0051_),
    .c(_0052_)
  );
  and_bi _2438_ (
    .a(_0048_),
    .b(_0052_),
    .c(_0053_)
  );
  or_bb _2439_ (
    .a(_0053_),
    .b(io_in2_3_),
    .c(_0054_)
  );
  or_bb _2440_ (
    .a(_1392_),
    .b(io_in2_1_),
    .c(_0055_)
  );
  and_bi _2441_ (
    .a(io_in2_1_),
    .b(_1398_),
    .c(_0056_)
  );
  and_bi _2442_ (
    .a(_0055_),
    .b(_0056_),
    .c(_0057_)
  );
  or_bb _2443_ (
    .a(_0057_),
    .b(io_in2_2_),
    .c(_0058_)
  );
  or_bb _2444_ (
    .a(_1402_),
    .b(io_in2_1_),
    .c(_0059_)
  );
  and_bi _2445_ (
    .a(io_in2_1_),
    .b(_1433_),
    .c(_0060_)
  );
  and_bi _2446_ (
    .a(_0059_),
    .b(_0060_),
    .c(_0061_)
  );
  and_bi _2447_ (
    .a(io_in2_2_),
    .b(_0061_),
    .c(_0062_)
  );
  and_bi _2448_ (
    .a(_0058_),
    .b(_0062_),
    .c(_0063_)
  );
  and_bi _2449_ (
    .a(io_in2_3_),
    .b(_0063_),
    .c(_0064_)
  );
  and_bi _2450_ (
    .a(_0054_),
    .b(_0064_),
    .c(_0065_)
  );
  and_bi _2451_ (
    .a(_1141_),
    .b(_0065_),
    .c(_0066_)
  );
  or_bb _2452_ (
    .a(_1437_),
    .b(io_in2_1_),
    .c(_0067_)
  );
  and_bi _2453_ (
    .a(io_in2_1_),
    .b(_1443_),
    .c(_0068_)
  );
  and_bi _2454_ (
    .a(_0067_),
    .b(_0068_),
    .c(_0069_)
  );
  or_bb _2455_ (
    .a(_0069_),
    .b(io_in2_2_),
    .c(_0070_)
  );
  or_bb _2456_ (
    .a(_1447_),
    .b(io_in2_1_),
    .c(_0071_)
  );
  and_bi _2457_ (
    .a(io_in2_1_),
    .b(_1455_),
    .c(_0072_)
  );
  and_bi _2458_ (
    .a(_0071_),
    .b(_0072_),
    .c(_0073_)
  );
  and_bi _2459_ (
    .a(io_in2_2_),
    .b(_0073_),
    .c(_0074_)
  );
  and_bi _2460_ (
    .a(_0070_),
    .b(_0074_),
    .c(_0075_)
  );
  or_bb _2461_ (
    .a(_0075_),
    .b(io_in2_3_),
    .c(_0076_)
  );
  and_bi _2462_ (
    .a(_0384_),
    .b(io_fn_3_),
    .c(_0077_)
  );
  and_bi _2463_ (
    .a(_1324_),
    .b(_0077_),
    .c(_0078_)
  );
  and_bi _2464_ (
    .a(io_in2_2_),
    .b(_0078_),
    .c(_0079_)
  );
  and_bi _2465_ (
    .a(_1190_),
    .b(_1459_),
    .c(_0080_)
  );
  and_bi _2466_ (
    .a(_1467_),
    .b(_1190_),
    .c(_0081_)
  );
  or_bb _2467_ (
    .a(_0081_),
    .b(_0080_),
    .c(_0082_)
  );
  and_bi _2468_ (
    .a(_0383_),
    .b(_0082_),
    .c(_0083_)
  );
  or_bb _2469_ (
    .a(_0083_),
    .b(_0079_),
    .c(_0084_)
  );
  and_bi _2470_ (
    .a(io_in2_3_),
    .b(_0084_),
    .c(_0085_)
  );
  and_bi _2471_ (
    .a(_0076_),
    .b(_0085_),
    .c(_0086_)
  );
  and_bi _2472_ (
    .a(io_in2_4_),
    .b(_0086_),
    .c(_0087_)
  );
  or_bb _2473_ (
    .a(_0087_),
    .b(_0066_),
    .c(_0088_)
  );
  and_bi _2474_ (
    .a(_1140_),
    .b(_0088_),
    .c(_0089_)
  );
  or_bb _2475_ (
    .a(_0089_),
    .b(_1477_),
    .c(_0090_)
  );
  and_bi _2476_ (
    .a(_0044_),
    .b(_0090_),
    .c(_0091_)
  );
  or_bb _2477_ (
    .a(_0091_),
    .b(_0026_),
    .c(io_out_3_)
  );
  and_bi _2478_ (
    .a(io_adder_out_4_),
    .b(_1121_),
    .c(_0092_)
  );
  and_bi _2479_ (
    .a(_0764_),
    .b(_0084_),
    .c(_0093_)
  );
  and_bi _2480_ (
    .a(_1362_),
    .b(_0093_),
    .c(_0094_)
  );
  and_bi _2481_ (
    .a(_1141_),
    .b(_0094_),
    .c(_0095_)
  );
  and_bi _2482_ (
    .a(_1361_),
    .b(_0095_),
    .c(_0096_)
  );
  and_bi _2483_ (
    .a(_1336_),
    .b(_0096_),
    .c(_0097_)
  );
  and_bi _2484_ (
    .a(_1343_),
    .b(_1141_),
    .c(_0098_)
  );
  or_bb _2485_ (
    .a(_0098_),
    .b(io_in1_4_),
    .c(_0099_)
  );
  and_bb _2486_ (
    .a(io_in2_4_),
    .b(io_in1_4_),
    .c(_0100_)
  );
  and_bb _2487_ (
    .a(_0100_),
    .b(_1341_),
    .c(_0101_)
  );
  and_bi _2488_ (
    .a(_0099_),
    .b(_0101_),
    .c(_0102_)
  );
  or_bb _2489_ (
    .a(_0102_),
    .b(_1345_),
    .c(_0103_)
  );
  and_bi _2490_ (
    .a(_1345_),
    .b(_0100_),
    .c(_0104_)
  );
  or_bb _2491_ (
    .a(_0104_),
    .b(_1336_),
    .c(_0105_)
  );
  and_bi _2492_ (
    .a(_0103_),
    .b(_0105_),
    .c(_0106_)
  );
  or_bb _2493_ (
    .a(_0106_),
    .b(_1140_),
    .c(_0107_)
  );
  or_bb _2494_ (
    .a(_0107_),
    .b(_0097_),
    .c(_0108_)
  );
  or_bb _2495_ (
    .a(_0028_),
    .b(_0764_),
    .c(_0109_)
  );
  and_bi _2496_ (
    .a(_0383_),
    .b(_1282_),
    .c(_0110_)
  );
  and_bi _2497_ (
    .a(io_in2_2_),
    .b(_1306_),
    .c(_0111_)
  );
  or_bb _2498_ (
    .a(_0111_),
    .b(_0110_),
    .c(_0112_)
  );
  and_bi _2499_ (
    .a(_0764_),
    .b(_0112_),
    .c(_0113_)
  );
  and_bi _2500_ (
    .a(_0109_),
    .b(_0113_),
    .c(_0114_)
  );
  and_bi _2501_ (
    .a(io_in2_4_),
    .b(_0114_),
    .c(_0115_)
  );
  or_ii _2502_ (
    .a(_1211_),
    .b(_0383_),
    .c(_0116_)
  );
  and_bi _2503_ (
    .a(io_in2_2_),
    .b(_1162_),
    .c(_0117_)
  );
  and_bi _2504_ (
    .a(_0116_),
    .b(_0117_),
    .c(_0118_)
  );
  and_bi _2505_ (
    .a(_0764_),
    .b(_0118_),
    .c(_0119_)
  );
  and_bi _2506_ (
    .a(_0383_),
    .b(_1186_),
    .c(_0120_)
  );
  and_bi _2507_ (
    .a(io_in2_2_),
    .b(_1260_),
    .c(_0121_)
  );
  or_bb _2508_ (
    .a(_0121_),
    .b(_0120_),
    .c(_0122_)
  );
  and_bi _2509_ (
    .a(_0122_),
    .b(_0764_),
    .c(_0123_)
  );
  or_bb _2510_ (
    .a(_0123_),
    .b(_0119_),
    .c(_0124_)
  );
  and_bi _2511_ (
    .a(_1141_),
    .b(_0124_),
    .c(_0125_)
  );
  or_bb _2512_ (
    .a(_0125_),
    .b(_0115_),
    .c(_0126_)
  );
  and_bb _2513_ (
    .a(_0126_),
    .b(_1140_),
    .c(_0127_)
  );
  or_bb _2514_ (
    .a(_0127_),
    .b(_1477_),
    .c(_0128_)
  );
  and_bi _2515_ (
    .a(_0108_),
    .b(_0128_),
    .c(_0129_)
  );
  or_bb _2516_ (
    .a(_0129_),
    .b(_0092_),
    .c(io_out_4_)
  );
  and_bi _2517_ (
    .a(io_adder_out_5_),
    .b(_1121_),
    .c(_0130_)
  );
  and_bi _2518_ (
    .a(_0764_),
    .b(_0018_),
    .c(_0131_)
  );
  and_bi _2519_ (
    .a(_1362_),
    .b(_0131_),
    .c(_0132_)
  );
  and_bi _2520_ (
    .a(_1141_),
    .b(_0132_),
    .c(_0133_)
  );
  and_bi _2521_ (
    .a(_1361_),
    .b(_0133_),
    .c(_0134_)
  );
  and_bi _2522_ (
    .a(_1336_),
    .b(_0134_),
    .c(_0135_)
  );
  and_bi _2523_ (
    .a(io_in1_5_),
    .b(_1345_),
    .c(_0136_)
  );
  and_bi _2524_ (
    .a(_1341_),
    .b(_0784_),
    .c(_0137_)
  );
  and_bi _2525_ (
    .a(_0136_),
    .b(_0137_),
    .c(_0138_)
  );
  and_bi _2526_ (
    .a(io_in2_5_),
    .b(_0136_),
    .c(_0139_)
  );
  or_bb _2527_ (
    .a(_0139_),
    .b(_0138_),
    .c(_0140_)
  );
  and_bi _2528_ (
    .a(_0782_),
    .b(_1343_),
    .c(_0141_)
  );
  or_bb _2529_ (
    .a(_0141_),
    .b(_1336_),
    .c(_0142_)
  );
  and_bi _2530_ (
    .a(_0140_),
    .b(_0142_),
    .c(_0143_)
  );
  or_bb _2531_ (
    .a(_0143_),
    .b(_1140_),
    .c(_0144_)
  );
  or_bb _2532_ (
    .a(_0144_),
    .b(_0135_),
    .c(_0145_)
  );
  or_bb _2533_ (
    .a(_1425_),
    .b(io_in2_2_),
    .c(_0146_)
  );
  and_bi _2534_ (
    .a(io_in2_2_),
    .b(_1394_),
    .c(_0147_)
  );
  and_bi _2535_ (
    .a(_0146_),
    .b(_0147_),
    .c(_0148_)
  );
  and_bi _2536_ (
    .a(_0764_),
    .b(_0148_),
    .c(_0149_)
  );
  and_bi _2537_ (
    .a(_0383_),
    .b(_1404_),
    .c(_0150_)
  );
  and_bi _2538_ (
    .a(io_in2_2_),
    .b(_1439_),
    .c(_0151_)
  );
  or_bb _2539_ (
    .a(_0151_),
    .b(_0150_),
    .c(_0152_)
  );
  and_bi _2540_ (
    .a(io_in2_3_),
    .b(_0152_),
    .c(_0153_)
  );
  or_bb _2541_ (
    .a(_0153_),
    .b(_0149_),
    .c(_0154_)
  );
  and_bi _2542_ (
    .a(_1141_),
    .b(_0154_),
    .c(_0155_)
  );
  and_bi _2543_ (
    .a(_1482_),
    .b(_0764_),
    .c(_0156_)
  );
  and_bi _2544_ (
    .a(_0383_),
    .b(_1449_),
    .c(_0157_)
  );
  and_bi _2545_ (
    .a(io_in2_2_),
    .b(_1461_),
    .c(_0158_)
  );
  or_bb _2546_ (
    .a(_0158_),
    .b(_0157_),
    .c(_0159_)
  );
  and_bi _2547_ (
    .a(_0764_),
    .b(_0159_),
    .c(_0160_)
  );
  or_bb _2548_ (
    .a(_0160_),
    .b(_0156_),
    .c(_0161_)
  );
  and_bi _2549_ (
    .a(io_in2_4_),
    .b(_0161_),
    .c(_0162_)
  );
  or_bb _2550_ (
    .a(_0162_),
    .b(_0155_),
    .c(_0163_)
  );
  and_bi _2551_ (
    .a(_1140_),
    .b(_0163_),
    .c(_0164_)
  );
  or_bb _2552_ (
    .a(_0164_),
    .b(_1477_),
    .c(_0165_)
  );
  and_bi _2553_ (
    .a(_0145_),
    .b(_0165_),
    .c(_0166_)
  );
  or_bb _2554_ (
    .a(_0166_),
    .b(_0130_),
    .c(io_out_5_)
  );
  and_bi _2555_ (
    .a(io_adder_out_6_),
    .b(_1121_),
    .c(_0167_)
  );
  and_bi _2556_ (
    .a(_0764_),
    .b(_1471_),
    .c(_0168_)
  );
  and_bi _2557_ (
    .a(_1362_),
    .b(_0168_),
    .c(_0169_)
  );
  and_bi _2558_ (
    .a(_1141_),
    .b(_0169_),
    .c(_0170_)
  );
  and_bi _2559_ (
    .a(_1361_),
    .b(_0170_),
    .c(_0171_)
  );
  and_bi _2560_ (
    .a(_1336_),
    .b(_0171_),
    .c(_0172_)
  );
  and_bb _2561_ (
    .a(_1343_),
    .b(io_in2_6_),
    .c(_0173_)
  );
  or_bb _2562_ (
    .a(_0173_),
    .b(io_in1_6_),
    .c(_0174_)
  );
  and_bb _2563_ (
    .a(io_in2_6_),
    .b(io_in1_6_),
    .c(_0175_)
  );
  and_bb _2564_ (
    .a(_0175_),
    .b(_1341_),
    .c(_0176_)
  );
  and_bi _2565_ (
    .a(_0174_),
    .b(_0176_),
    .c(_0177_)
  );
  or_bb _2566_ (
    .a(_0177_),
    .b(_1345_),
    .c(_0178_)
  );
  and_bi _2567_ (
    .a(_1345_),
    .b(_0175_),
    .c(_0179_)
  );
  or_bb _2568_ (
    .a(_0179_),
    .b(_1336_),
    .c(_0180_)
  );
  and_bi _2569_ (
    .a(_0178_),
    .b(_0180_),
    .c(_0181_)
  );
  or_bb _2570_ (
    .a(_0181_),
    .b(_1140_),
    .c(_0182_)
  );
  or_bb _2571_ (
    .a(_0182_),
    .b(_0172_),
    .c(_0183_)
  );
  or_bb _2572_ (
    .a(_1505_),
    .b(io_in2_2_),
    .c(_0184_)
  );
  and_bi _2573_ (
    .a(io_in2_2_),
    .b(_1511_),
    .c(_0185_)
  );
  and_bi _2574_ (
    .a(_0184_),
    .b(_0185_),
    .c(_0186_)
  );
  and_bi _2575_ (
    .a(_0764_),
    .b(_0186_),
    .c(_0187_)
  );
  and_bi _2576_ (
    .a(_0383_),
    .b(_1515_),
    .c(_0188_)
  );
  and_bi _2577_ (
    .a(io_in2_2_),
    .b(_0005_),
    .c(_0189_)
  );
  or_bb _2578_ (
    .a(_0189_),
    .b(_0188_),
    .c(_0190_)
  );
  and_bi _2579_ (
    .a(io_in2_3_),
    .b(_0190_),
    .c(_0191_)
  );
  or_bb _2580_ (
    .a(_0191_),
    .b(_0187_),
    .c(_0192_)
  );
  and_bi _2581_ (
    .a(_1141_),
    .b(_0192_),
    .c(_0193_)
  );
  and_bi _2582_ (
    .a(_1369_),
    .b(_0764_),
    .c(_0194_)
  );
  and_bi _2583_ (
    .a(_0383_),
    .b(_0009_),
    .c(_0195_)
  );
  and_bi _2584_ (
    .a(_0016_),
    .b(_0383_),
    .c(_0196_)
  );
  or_bb _2585_ (
    .a(_0196_),
    .b(_0195_),
    .c(_0197_)
  );
  and_bi _2586_ (
    .a(_0764_),
    .b(_0197_),
    .c(_0198_)
  );
  or_bb _2587_ (
    .a(_0198_),
    .b(_0194_),
    .c(_0199_)
  );
  and_bi _2588_ (
    .a(io_in2_4_),
    .b(_0199_),
    .c(_0200_)
  );
  or_bb _2589_ (
    .a(_0200_),
    .b(_0193_),
    .c(_0201_)
  );
  and_bi _2590_ (
    .a(_1140_),
    .b(_0201_),
    .c(_0202_)
  );
  or_bb _2591_ (
    .a(_0202_),
    .b(_1477_),
    .c(_0203_)
  );
  and_bi _2592_ (
    .a(_0183_),
    .b(_0203_),
    .c(_0204_)
  );
  or_bb _2593_ (
    .a(_0204_),
    .b(_0167_),
    .c(io_out_6_)
  );
  and_bi _2594_ (
    .a(io_adder_out_7_),
    .b(_1121_),
    .c(_0205_)
  );
  and_bi _2595_ (
    .a(_0764_),
    .b(_1330_),
    .c(_0206_)
  );
  and_bi _2596_ (
    .a(_1362_),
    .b(_0206_),
    .c(_0207_)
  );
  and_bi _2597_ (
    .a(_1141_),
    .b(_0207_),
    .c(_0208_)
  );
  and_bi _2598_ (
    .a(_1361_),
    .b(_0208_),
    .c(_0209_)
  );
  and_bi _2599_ (
    .a(_1336_),
    .b(_0209_),
    .c(_0210_)
  );
  or_bb _2600_ (
    .a(_1345_),
    .b(_0741_),
    .c(_0211_)
  );
  and_bi _2601_ (
    .a(_0741_),
    .b(_1343_),
    .c(_0212_)
  );
  or_bb _2602_ (
    .a(_0212_),
    .b(_0803_),
    .c(_0213_)
  );
  or_ii _2603_ (
    .a(_0213_),
    .b(_0211_),
    .c(_0214_)
  );
  and_bi _2604_ (
    .a(_1341_),
    .b(_0803_),
    .c(_0215_)
  );
  and_bi _2605_ (
    .a(_0215_),
    .b(_0211_),
    .c(_0216_)
  );
  or_bb _2606_ (
    .a(_0216_),
    .b(_1336_),
    .c(_0217_)
  );
  and_bi _2607_ (
    .a(_0214_),
    .b(_0217_),
    .c(_0218_)
  );
  or_bb _2608_ (
    .a(_0218_),
    .b(_1140_),
    .c(_0219_)
  );
  or_bb _2609_ (
    .a(_0219_),
    .b(_0210_),
    .c(_0220_)
  );
  or_bb _2610_ (
    .a(_0051_),
    .b(io_in2_2_),
    .c(_0221_)
  );
  and_bi _2611_ (
    .a(io_in2_2_),
    .b(_0057_),
    .c(_0222_)
  );
  and_bi _2612_ (
    .a(_0221_),
    .b(_0222_),
    .c(_0223_)
  );
  and_bi _2613_ (
    .a(_0764_),
    .b(_0223_),
    .c(_0224_)
  );
  and_bi _2614_ (
    .a(_0383_),
    .b(_0061_),
    .c(_0225_)
  );
  and_bi _2615_ (
    .a(io_in2_2_),
    .b(_0069_),
    .c(_0226_)
  );
  or_bb _2616_ (
    .a(_0226_),
    .b(_0225_),
    .c(_0227_)
  );
  and_bi _2617_ (
    .a(_0227_),
    .b(_0764_),
    .c(_0228_)
  );
  or_bb _2618_ (
    .a(_0228_),
    .b(_0224_),
    .c(_0229_)
  );
  and_bi _2619_ (
    .a(_1141_),
    .b(_0229_),
    .c(_0230_)
  );
  or_bb _2620_ (
    .a(_0073_),
    .b(io_in2_2_),
    .c(_0231_)
  );
  and_bi _2621_ (
    .a(_0082_),
    .b(_0383_),
    .c(_0232_)
  );
  and_bi _2622_ (
    .a(_0231_),
    .b(_0232_),
    .c(_0233_)
  );
  and_bi _2623_ (
    .a(_0764_),
    .b(_0233_),
    .c(_0234_)
  );
  and_bi _2624_ (
    .a(_0352_),
    .b(_0394_),
    .c(_0235_)
  );
  or_bb _2625_ (
    .a(_0235_),
    .b(_0764_),
    .c(_0236_)
  );
  and_bi _2626_ (
    .a(_1324_),
    .b(_0236_),
    .c(_0237_)
  );
  or_bb _2627_ (
    .a(_0237_),
    .b(_0234_),
    .c(_0238_)
  );
  and_bi _2628_ (
    .a(io_in2_4_),
    .b(_0238_),
    .c(_0239_)
  );
  or_bb _2629_ (
    .a(_0239_),
    .b(_0230_),
    .c(_0240_)
  );
  and_bb _2630_ (
    .a(_0240_),
    .b(_1140_),
    .c(_0241_)
  );
  or_bb _2631_ (
    .a(_0241_),
    .b(_1477_),
    .c(_0242_)
  );
  and_bi _2632_ (
    .a(_0220_),
    .b(_0242_),
    .c(_0243_)
  );
  or_bb _2633_ (
    .a(_0243_),
    .b(_0205_),
    .c(io_out_7_)
  );
  and_bi _2634_ (
    .a(io_adder_out_8_),
    .b(_1121_),
    .c(_0244_)
  );
  and_bi _2635_ (
    .a(_0238_),
    .b(io_in2_4_),
    .c(_0245_)
  );
  and_bi _2636_ (
    .a(_1361_),
    .b(_0245_),
    .c(_0246_)
  );
  and_bi _2637_ (
    .a(_1336_),
    .b(_0246_),
    .c(_0247_)
  );
  and_bi _2638_ (
    .a(io_in1_8_),
    .b(_1345_),
    .c(_0248_)
  );
  and_bi _2639_ (
    .a(_0812_),
    .b(_1343_),
    .c(_0249_)
  );
  and_bi _2640_ (
    .a(io_in2_8_),
    .b(_0249_),
    .c(_0250_)
  );
  or_bb _2641_ (
    .a(_0250_),
    .b(_0248_),
    .c(_0251_)
  );
  and_bb _2642_ (
    .a(_1341_),
    .b(io_in2_8_),
    .c(_0252_)
  );
  and_bb _2643_ (
    .a(_0252_),
    .b(_0248_),
    .c(_0253_)
  );
  or_bb _2644_ (
    .a(_0253_),
    .b(_1336_),
    .c(_0254_)
  );
  and_bi _2645_ (
    .a(_0251_),
    .b(_0254_),
    .c(_0255_)
  );
  or_bb _2646_ (
    .a(_0255_),
    .b(_1140_),
    .c(_0256_)
  );
  or_bb _2647_ (
    .a(_0256_),
    .b(_0247_),
    .c(_0257_)
  );
  and_bi _2648_ (
    .a(_0764_),
    .b(_1188_),
    .c(_0258_)
  );
  and_bi _2649_ (
    .a(io_in2_3_),
    .b(_1284_),
    .c(_0259_)
  );
  or_bb _2650_ (
    .a(_0259_),
    .b(_0258_),
    .c(_0260_)
  );
  and_bi _2651_ (
    .a(_1141_),
    .b(_0260_),
    .c(_0261_)
  );
  and_bi _2652_ (
    .a(io_in2_4_),
    .b(_0207_),
    .c(_0262_)
  );
  or_bb _2653_ (
    .a(_0262_),
    .b(_0261_),
    .c(_0263_)
  );
  and_bi _2654_ (
    .a(_1140_),
    .b(_0263_),
    .c(_0264_)
  );
  or_bb _2655_ (
    .a(_0264_),
    .b(_1477_),
    .c(_0265_)
  );
  and_bi _2656_ (
    .a(_0257_),
    .b(_0265_),
    .c(_0266_)
  );
  or_bb _2657_ (
    .a(_0266_),
    .b(_0244_),
    .c(io_out_8_)
  );
  and_bi _2658_ (
    .a(io_adder_out_9_),
    .b(_1121_),
    .c(_0267_)
  );
  and_bi _2659_ (
    .a(_1141_),
    .b(_0199_),
    .c(_0268_)
  );
  and_bi _2660_ (
    .a(_1361_),
    .b(_0268_),
    .c(_0269_)
  );
  and_bi _2661_ (
    .a(_1336_),
    .b(_0269_),
    .c(_0270_)
  );
  and_bi _2662_ (
    .a(_0821_),
    .b(_1343_),
    .c(_0271_)
  );
  and_bi _2663_ (
    .a(io_in1_9_),
    .b(_1345_),
    .c(_0272_)
  );
  or_bb _2664_ (
    .a(_0272_),
    .b(_0823_),
    .c(_0273_)
  );
  or_bb _2665_ (
    .a(_0273_),
    .b(_0271_),
    .c(_0274_)
  );
  and_bi _2666_ (
    .a(_1341_),
    .b(_0823_),
    .c(_0275_)
  );
  and_bi _2667_ (
    .a(_0272_),
    .b(_0275_),
    .c(_0276_)
  );
  and_bi _2668_ (
    .a(_0274_),
    .b(_0276_),
    .c(_0277_)
  );
  and_bi _2669_ (
    .a(_1337_),
    .b(_0277_),
    .c(_0278_)
  );
  or_bb _2670_ (
    .a(_0278_),
    .b(_1140_),
    .c(_0279_)
  );
  or_bb _2671_ (
    .a(_0279_),
    .b(_0270_),
    .c(_0280_)
  );
  and_bi _2672_ (
    .a(_0764_),
    .b(_1406_),
    .c(_0281_)
  );
  and_bi _2673_ (
    .a(io_in2_3_),
    .b(_1451_),
    .c(_0282_)
  );
  or_bb _2674_ (
    .a(_0282_),
    .b(io_in2_4_),
    .c(_0283_)
  );
  or_bb _2675_ (
    .a(_0283_),
    .b(_0281_),
    .c(_0284_)
  );
  and_bi _2676_ (
    .a(_0169_),
    .b(_1141_),
    .c(_0285_)
  );
  or_bi _2677_ (
    .a(_0285_),
    .b(_0284_),
    .c(_0286_)
  );
  and_bb _2678_ (
    .a(_0286_),
    .b(_1140_),
    .c(_0287_)
  );
  or_bb _2679_ (
    .a(_0287_),
    .b(_1477_),
    .c(_0288_)
  );
  and_bi _2680_ (
    .a(_0280_),
    .b(_0288_),
    .c(_0289_)
  );
  or_bb _2681_ (
    .a(_0289_),
    .b(_0267_),
    .c(io_out_9_)
  );
  and_bi _2682_ (
    .a(io_adder_out_10_),
    .b(_1121_),
    .c(_0290_)
  );
  and_bi _2683_ (
    .a(_1141_),
    .b(_0161_),
    .c(_0291_)
  );
  and_bi _2684_ (
    .a(_1361_),
    .b(_0291_),
    .c(_0292_)
  );
  and_bi _2685_ (
    .a(_1336_),
    .b(_0292_),
    .c(_0293_)
  );
  and_bi _2686_ (
    .a(_0832_),
    .b(_1343_),
    .c(_0294_)
  );
  inv _2687_ (
    .din(io_in2_10_),
    .dout(_0295_)
  );
  and_bi _2688_ (
    .a(io_in1_10_),
    .b(_1345_),
    .c(_0296_)
  );
  or_bb _2689_ (
    .a(_0296_),
    .b(_0295_),
    .c(_0297_)
  );
  or_bb _2690_ (
    .a(_0297_),
    .b(_0294_),
    .c(_0298_)
  );
  and_bi _2691_ (
    .a(_1341_),
    .b(_0295_),
    .c(_0299_)
  );
  and_bi _2692_ (
    .a(_0296_),
    .b(_0299_),
    .c(_0300_)
  );
  and_bi _2693_ (
    .a(_0298_),
    .b(_0300_),
    .c(_0301_)
  );
  and_bi _2694_ (
    .a(_1337_),
    .b(_0301_),
    .c(_0302_)
  );
  or_bb _2695_ (
    .a(_0302_),
    .b(_1140_),
    .c(_0303_)
  );
  or_bb _2696_ (
    .a(_0303_),
    .b(_0293_),
    .c(_0304_)
  );
  and_bi _2697_ (
    .a(_0764_),
    .b(_1517_),
    .c(_0305_)
  );
  and_bi _2698_ (
    .a(io_in2_3_),
    .b(_0011_),
    .c(_0306_)
  );
  or_bb _2699_ (
    .a(_0306_),
    .b(io_in2_4_),
    .c(_0307_)
  );
  or_bb _2700_ (
    .a(_0307_),
    .b(_0305_),
    .c(_0308_)
  );
  and_bi _2701_ (
    .a(_0132_),
    .b(_1141_),
    .c(_0309_)
  );
  or_bi _2702_ (
    .a(_0309_),
    .b(_0308_),
    .c(_0310_)
  );
  and_bb _2703_ (
    .a(_0310_),
    .b(_1140_),
    .c(_0311_)
  );
  or_bb _2704_ (
    .a(_0311_),
    .b(_1477_),
    .c(_0312_)
  );
  and_bi _2705_ (
    .a(_0304_),
    .b(_0312_),
    .c(_0313_)
  );
  or_bb _2706_ (
    .a(_0313_),
    .b(_0290_),
    .c(io_out_10_)
  );
  and_bi _2707_ (
    .a(io_adder_out_11_),
    .b(_1121_),
    .c(_0314_)
  );
  and_bi _2708_ (
    .a(_0114_),
    .b(io_in2_4_),
    .c(_0315_)
  );
  and_bi _2709_ (
    .a(_1361_),
    .b(_0315_),
    .c(_0316_)
  );
  and_bi _2710_ (
    .a(_1336_),
    .b(_0316_),
    .c(_0317_)
  );
  and_bi _2711_ (
    .a(io_in1_11_),
    .b(_1345_),
    .c(_0318_)
  );
  and_bi _2712_ (
    .a(_0740_),
    .b(_1343_),
    .c(_0319_)
  );
  and_bi _2713_ (
    .a(io_in2_11_),
    .b(_0319_),
    .c(_0320_)
  );
  or_bb _2714_ (
    .a(_0320_),
    .b(_0318_),
    .c(_0321_)
  );
  and_bi _2715_ (
    .a(_1341_),
    .b(_0844_),
    .c(_0322_)
  );
  and_bb _2716_ (
    .a(_0322_),
    .b(_0318_),
    .c(_0323_)
  );
  or_bb _2717_ (
    .a(_0323_),
    .b(_1336_),
    .c(_0324_)
  );
  and_bi _2718_ (
    .a(_0321_),
    .b(_0324_),
    .c(_0325_)
  );
  or_bb _2719_ (
    .a(_0325_),
    .b(_1140_),
    .c(_0326_)
  );
  or_bb _2720_ (
    .a(_0326_),
    .b(_0317_),
    .c(_0327_)
  );
  and_bi _2721_ (
    .a(_0764_),
    .b(_0063_),
    .c(_0328_)
  );
  and_bi _2722_ (
    .a(io_in2_3_),
    .b(_0075_),
    .c(_0329_)
  );
  or_bb _2723_ (
    .a(_0329_),
    .b(io_in2_4_),
    .c(_0330_)
  );
  or_bb _2724_ (
    .a(_0330_),
    .b(_0328_),
    .c(_0331_)
  );
  and_bi _2725_ (
    .a(_0094_),
    .b(_1141_),
    .c(_0332_)
  );
  or_bi _2726_ (
    .a(_0332_),
    .b(_0331_),
    .c(_0333_)
  );
  and_bb _2727_ (
    .a(_0333_),
    .b(_1140_),
    .c(_0334_)
  );
  or_bb _2728_ (
    .a(_0334_),
    .b(_1477_),
    .c(_0335_)
  );
  and_bi _2729_ (
    .a(_0327_),
    .b(_0335_),
    .c(_0336_)
  );
  or_bb _2730_ (
    .a(_0336_),
    .b(_0314_),
    .c(io_out_11_)
  );
  and_bi _2731_ (
    .a(_1141_),
    .b(_0086_),
    .c(_0337_)
  );
  and_bi _2732_ (
    .a(_1361_),
    .b(_0337_),
    .c(_0338_)
  );
  and_bi _2733_ (
    .a(_1336_),
    .b(_0338_),
    .c(_0339_)
  );
  and_bi _2734_ (
    .a(io_in1_12_),
    .b(_1345_),
    .c(_0342_)
  );
  and_bi _2735_ (
    .a(_0850_),
    .b(_1343_),
    .c(_0343_)
  );
  and_bi _2736_ (
    .a(io_in2_12_),
    .b(_0343_),
    .c(_0344_)
  );
  or_bb _2737_ (
    .a(_0344_),
    .b(_0342_),
    .c(_0345_)
  );
  and_bb _2738_ (
    .a(_1341_),
    .b(io_in2_12_),
    .c(_0346_)
  );
  and_bb _2739_ (
    .a(_0346_),
    .b(_0342_),
    .c(_0347_)
  );
  or_bb _2740_ (
    .a(_0347_),
    .b(_1336_),
    .c(_0348_)
  );
  and_bi _2741_ (
    .a(_0345_),
    .b(_0348_),
    .c(_0349_)
  );
  or_bb _2742_ (
    .a(_0349_),
    .b(_1140_),
    .c(_0350_)
  );
  or_bb _2743_ (
    .a(_0350_),
    .b(_0339_),
    .c(_0351_)
  );
  and_bi _2744_ (
    .a(_0764_),
    .b(_0122_),
    .c(_0353_)
  );
  and_bi _2745_ (
    .a(io_in2_3_),
    .b(_0112_),
    .c(_0354_)
  );
  or_bb _2746_ (
    .a(_0354_),
    .b(_0353_),
    .c(_0355_)
  );
  and_bi _2747_ (
    .a(_1141_),
    .b(_0355_),
    .c(_0356_)
  );
  and_bi _2748_ (
    .a(io_in2_4_),
    .b(_0030_),
    .c(_0357_)
  );
  or_bb _2749_ (
    .a(_0357_),
    .b(_0356_),
    .c(_0358_)
  );
  and_bi _2750_ (
    .a(_1140_),
    .b(_0358_),
    .c(_0359_)
  );
  or_bb _2751_ (
    .a(_0359_),
    .b(_1477_),
    .c(_0360_)
  );
  and_bi _2752_ (
    .a(_0351_),
    .b(_0360_),
    .c(_0361_)
  );
  and_bi _2753_ (
    .a(io_adder_out_12_),
    .b(_1121_),
    .c(_0362_)
  );
  or_bb _2754_ (
    .a(_0362_),
    .b(_0361_),
    .c(io_out_12_)
  );
  and_bi _2755_ (
    .a(io_adder_out_13_),
    .b(_1121_),
    .c(_0364_)
  );
  and_bi _2756_ (
    .a(_0020_),
    .b(io_in2_4_),
    .c(_0365_)
  );
  and_bi _2757_ (
    .a(_1361_),
    .b(_0365_),
    .c(_0366_)
  );
  and_bi _2758_ (
    .a(_1336_),
    .b(_0366_),
    .c(_0367_)
  );
  or_bb _2759_ (
    .a(_1345_),
    .b(_0739_),
    .c(_0368_)
  );
  and_bi _2760_ (
    .a(_0739_),
    .b(_1343_),
    .c(_0369_)
  );
  or_bb _2761_ (
    .a(_0369_),
    .b(_0862_),
    .c(_0370_)
  );
  or_ii _2762_ (
    .a(_0370_),
    .b(_0368_),
    .c(_0371_)
  );
  and_bi _2763_ (
    .a(_1341_),
    .b(_0862_),
    .c(_0372_)
  );
  and_bi _2764_ (
    .a(_0372_),
    .b(_0368_),
    .c(_0373_)
  );
  or_bb _2765_ (
    .a(_0373_),
    .b(_1336_),
    .c(_0374_)
  );
  and_bi _2766_ (
    .a(_0371_),
    .b(_0374_),
    .c(_0375_)
  );
  or_bb _2767_ (
    .a(_0375_),
    .b(_1140_),
    .c(_0376_)
  );
  or_bb _2768_ (
    .a(_0376_),
    .b(_0367_),
    .c(_0377_)
  );
  and_bi _2769_ (
    .a(_0764_),
    .b(_0152_),
    .c(_0378_)
  );
  and_bi _2770_ (
    .a(io_in2_3_),
    .b(_0159_),
    .c(_0379_)
  );
  or_bb _2771_ (
    .a(_0379_),
    .b(_0378_),
    .c(_0380_)
  );
  and_bi _2772_ (
    .a(_1141_),
    .b(_0380_),
    .c(_0381_)
  );
  and_bi _2773_ (
    .a(io_in2_4_),
    .b(_1484_),
    .c(_0382_)
  );
  or_bb _2774_ (
    .a(_0382_),
    .b(_0381_),
    .c(_0385_)
  );
  and_bi _2775_ (
    .a(_1140_),
    .b(_0385_),
    .c(_0386_)
  );
  or_bb _2776_ (
    .a(_0386_),
    .b(_1477_),
    .c(_0387_)
  );
  and_bi _2777_ (
    .a(_0377_),
    .b(_0387_),
    .c(_0388_)
  );
  or_bb _2778_ (
    .a(_0388_),
    .b(_0364_),
    .c(io_out_13_)
  );
  and_bi _2779_ (
    .a(io_adder_out_14_),
    .b(_1121_),
    .c(_0389_)
  );
  and_bi _2780_ (
    .a(_1141_),
    .b(_1473_),
    .c(_0390_)
  );
  and_bi _2781_ (
    .a(_1361_),
    .b(_0390_),
    .c(_0391_)
  );
  and_bi _2782_ (
    .a(_1336_),
    .b(_0391_),
    .c(_0392_)
  );
  and_bb _2783_ (
    .a(_1343_),
    .b(io_in2_14_),
    .c(_0393_)
  );
  or_bb _2784_ (
    .a(_0393_),
    .b(io_in1_14_),
    .c(_0395_)
  );
  and_bb _2785_ (
    .a(io_in2_14_),
    .b(io_in1_14_),
    .c(_0396_)
  );
  and_bb _2786_ (
    .a(_0396_),
    .b(_1341_),
    .c(_0397_)
  );
  and_bi _2787_ (
    .a(_0395_),
    .b(_0397_),
    .c(_0398_)
  );
  or_bb _2788_ (
    .a(_0398_),
    .b(_1345_),
    .c(_0399_)
  );
  and_bi _2789_ (
    .a(_1345_),
    .b(_0396_),
    .c(_0400_)
  );
  or_bb _2790_ (
    .a(_0400_),
    .b(_1336_),
    .c(_0401_)
  );
  and_bi _2791_ (
    .a(_0399_),
    .b(_0401_),
    .c(_0402_)
  );
  or_bb _2792_ (
    .a(_0402_),
    .b(_1140_),
    .c(_0403_)
  );
  or_bb _2793_ (
    .a(_0403_),
    .b(_0392_),
    .c(_0404_)
  );
  and_bi _2794_ (
    .a(_0764_),
    .b(_0190_),
    .c(_0406_)
  );
  and_bi _2795_ (
    .a(io_in2_3_),
    .b(_0197_),
    .c(_0407_)
  );
  or_bb _2796_ (
    .a(_0407_),
    .b(_0406_),
    .c(_0408_)
  );
  and_bi _2797_ (
    .a(_1141_),
    .b(_0408_),
    .c(_0409_)
  );
  and_bi _2798_ (
    .a(io_in2_4_),
    .b(_1371_),
    .c(_0410_)
  );
  or_bb _2799_ (
    .a(_0410_),
    .b(_0409_),
    .c(_0411_)
  );
  and_bi _2800_ (
    .a(_1140_),
    .b(_0411_),
    .c(_0412_)
  );
  or_bb _2801_ (
    .a(_0412_),
    .b(_1477_),
    .c(_0413_)
  );
  and_bi _2802_ (
    .a(_0404_),
    .b(_0413_),
    .c(_0414_)
  );
  or_bb _2803_ (
    .a(_0414_),
    .b(_0389_),
    .c(io_out_14_)
  );
  and_bi _2804_ (
    .a(io_adder_out_15_),
    .b(_1121_),
    .c(_0416_)
  );
  and_bi _2805_ (
    .a(_1141_),
    .b(_1332_),
    .c(_0417_)
  );
  and_bi _2806_ (
    .a(_1361_),
    .b(_0417_),
    .c(_0418_)
  );
  and_bi _2807_ (
    .a(_1336_),
    .b(_0418_),
    .c(_0419_)
  );
  and_bi _2808_ (
    .a(_0877_),
    .b(_1343_),
    .c(_0420_)
  );
  and_bi _2809_ (
    .a(io_in1_15_),
    .b(_1345_),
    .c(_0421_)
  );
  or_bb _2810_ (
    .a(_0421_),
    .b(_0879_),
    .c(_0422_)
  );
  or_bb _2811_ (
    .a(_0422_),
    .b(_0420_),
    .c(_0423_)
  );
  and_bi _2812_ (
    .a(_1341_),
    .b(_0879_),
    .c(_0424_)
  );
  and_bi _2813_ (
    .a(_0421_),
    .b(_0424_),
    .c(_0425_)
  );
  and_bi _2814_ (
    .a(_0423_),
    .b(_0425_),
    .c(_0426_)
  );
  and_bi _2815_ (
    .a(_1337_),
    .b(_0426_),
    .c(_0427_)
  );
  or_bb _2816_ (
    .a(_0427_),
    .b(_1140_),
    .c(_0428_)
  );
  or_bb _2817_ (
    .a(_0428_),
    .b(_0419_),
    .c(_0429_)
  );
  and_bi _2818_ (
    .a(_0352_),
    .b(_0405_),
    .c(_0430_)
  );
  and_bi _2819_ (
    .a(io_in2_4_),
    .b(_0430_),
    .c(_0431_)
  );
  or_ii _2820_ (
    .a(_0431_),
    .b(_1324_),
    .c(_0432_)
  );
  or_ii _2821_ (
    .a(_0233_),
    .b(io_in2_3_),
    .c(_0433_)
  );
  and_bi _2822_ (
    .a(_0764_),
    .b(_0227_),
    .c(_0434_)
  );
  or_bb _2823_ (
    .a(_0434_),
    .b(io_in2_4_),
    .c(_0435_)
  );
  and_bi _2824_ (
    .a(_0433_),
    .b(_0435_),
    .c(_0438_)
  );
  and_bi _2825_ (
    .a(_0432_),
    .b(_0438_),
    .c(_0439_)
  );
  and_bb _2826_ (
    .a(_0439_),
    .b(_1140_),
    .c(_0440_)
  );
  or_bb _2827_ (
    .a(_0440_),
    .b(_1477_),
    .c(_0441_)
  );
  and_bi _2828_ (
    .a(_0429_),
    .b(_0441_),
    .c(_0442_)
  );
  or_bb _2829_ (
    .a(_0442_),
    .b(_0416_),
    .c(io_out_15_)
  );
  and_bi _2830_ (
    .a(io_adder_out_16_),
    .b(_1121_),
    .c(_0443_)
  );
  and_bi _2831_ (
    .a(_1336_),
    .b(_0439_),
    .c(_0444_)
  );
  and_bb _2832_ (
    .a(_1343_),
    .b(io_in2_16_),
    .c(_0445_)
  );
  or_bb _2833_ (
    .a(_0445_),
    .b(io_in1_16_),
    .c(_0446_)
  );
  and_bb _2834_ (
    .a(io_in2_16_),
    .b(io_in1_16_),
    .c(_0448_)
  );
  and_bb _2835_ (
    .a(_0448_),
    .b(_1341_),
    .c(_0449_)
  );
  and_bi _2836_ (
    .a(_0446_),
    .b(_0449_),
    .c(_0450_)
  );
  or_bb _2837_ (
    .a(_0450_),
    .b(_1345_),
    .c(_0451_)
  );
  and_bi _2838_ (
    .a(_1345_),
    .b(_0448_),
    .c(_0452_)
  );
  or_bb _2839_ (
    .a(_0452_),
    .b(_1336_),
    .c(_0453_)
  );
  and_bi _2840_ (
    .a(_0451_),
    .b(_0453_),
    .c(_0454_)
  );
  or_bb _2841_ (
    .a(_0454_),
    .b(_1140_),
    .c(_0455_)
  );
  or_bb _2842_ (
    .a(_0455_),
    .b(_0444_),
    .c(_0456_)
  );
  and_bb _2843_ (
    .a(_0418_),
    .b(_1140_),
    .c(_0457_)
  );
  or_bb _2844_ (
    .a(_0457_),
    .b(_1477_),
    .c(_0459_)
  );
  and_bi _2845_ (
    .a(_0456_),
    .b(_0459_),
    .c(_0460_)
  );
  or_bb _2846_ (
    .a(_0460_),
    .b(_0443_),
    .c(io_out_16_)
  );
  and_bi _2847_ (
    .a(io_adder_out_17_),
    .b(_1121_),
    .c(_0461_)
  );
  and_bi _2848_ (
    .a(_0411_),
    .b(_1337_),
    .c(_0462_)
  );
  and_bi _2849_ (
    .a(_1343_),
    .b(_0898_),
    .c(_0463_)
  );
  or_bb _2850_ (
    .a(_0463_),
    .b(io_in1_17_),
    .c(_0464_)
  );
  and_bb _2851_ (
    .a(io_in2_17_),
    .b(io_in1_17_),
    .c(_0465_)
  );
  and_bb _2852_ (
    .a(_0465_),
    .b(_1341_),
    .c(_0466_)
  );
  and_bi _2853_ (
    .a(_0464_),
    .b(_0466_),
    .c(_0467_)
  );
  or_bb _2854_ (
    .a(_0467_),
    .b(_1345_),
    .c(_0468_)
  );
  and_bi _2855_ (
    .a(_1345_),
    .b(_0465_),
    .c(_0469_)
  );
  or_bb _2856_ (
    .a(_0469_),
    .b(_1336_),
    .c(_0470_)
  );
  and_bi _2857_ (
    .a(_0468_),
    .b(_0470_),
    .c(_0471_)
  );
  or_bb _2858_ (
    .a(_0471_),
    .b(_1140_),
    .c(_0472_)
  );
  or_bb _2859_ (
    .a(_0472_),
    .b(_0462_),
    .c(_0473_)
  );
  and_bb _2860_ (
    .a(_0391_),
    .b(_1140_),
    .c(_0474_)
  );
  or_bb _2861_ (
    .a(_0474_),
    .b(_1477_),
    .c(_0475_)
  );
  and_bi _2862_ (
    .a(_0473_),
    .b(_0475_),
    .c(_0476_)
  );
  or_bb _2863_ (
    .a(_0476_),
    .b(_0461_),
    .c(io_out_17_)
  );
  and_bi _2864_ (
    .a(io_adder_out_18_),
    .b(_1121_),
    .c(_0479_)
  );
  and_bi _2865_ (
    .a(_0385_),
    .b(_1337_),
    .c(_0480_)
  );
  and_bb _2866_ (
    .a(_1343_),
    .b(io_in2_18_),
    .c(_0481_)
  );
  or_bb _2867_ (
    .a(_0481_),
    .b(io_in1_18_),
    .c(_0482_)
  );
  and_bb _2868_ (
    .a(io_in2_18_),
    .b(io_in1_18_),
    .c(_0483_)
  );
  and_bb _2869_ (
    .a(_0483_),
    .b(_1341_),
    .c(_0484_)
  );
  and_bi _2870_ (
    .a(_0482_),
    .b(_0484_),
    .c(_0485_)
  );
  or_bb _2871_ (
    .a(_0485_),
    .b(_1345_),
    .c(_0486_)
  );
  and_bi _2872_ (
    .a(_1345_),
    .b(_0483_),
    .c(_0487_)
  );
  or_bb _2873_ (
    .a(_0487_),
    .b(_1336_),
    .c(_0488_)
  );
  and_bi _2874_ (
    .a(_0486_),
    .b(_0488_),
    .c(_0490_)
  );
  or_bb _2875_ (
    .a(_0490_),
    .b(_1140_),
    .c(_0491_)
  );
  or_bb _2876_ (
    .a(_0491_),
    .b(_0480_),
    .c(_0492_)
  );
  and_bb _2877_ (
    .a(_0366_),
    .b(_1140_),
    .c(_0493_)
  );
  or_bb _2878_ (
    .a(_0493_),
    .b(_1477_),
    .c(_0494_)
  );
  and_bi _2879_ (
    .a(_0492_),
    .b(_0494_),
    .c(_0495_)
  );
  or_bb _2880_ (
    .a(_0495_),
    .b(_0479_),
    .c(io_out_18_)
  );
  and_bi _2881_ (
    .a(io_adder_out_19_),
    .b(_1121_),
    .c(_0496_)
  );
  and_bi _2882_ (
    .a(_0358_),
    .b(_1337_),
    .c(_0497_)
  );
  and_bi _2883_ (
    .a(_1343_),
    .b(_0916_),
    .c(_0498_)
  );
  or_bb _2884_ (
    .a(_0498_),
    .b(io_in1_19_),
    .c(_0500_)
  );
  and_bb _2885_ (
    .a(io_in2_19_),
    .b(io_in1_19_),
    .c(_0501_)
  );
  and_bb _2886_ (
    .a(_0501_),
    .b(_1341_),
    .c(_0502_)
  );
  and_bi _2887_ (
    .a(_0500_),
    .b(_0502_),
    .c(_0503_)
  );
  or_bb _2888_ (
    .a(_0503_),
    .b(_1345_),
    .c(_0504_)
  );
  and_bi _2889_ (
    .a(_1345_),
    .b(_0501_),
    .c(_0505_)
  );
  or_bb _2890_ (
    .a(_0505_),
    .b(_1336_),
    .c(_0506_)
  );
  and_bi _2891_ (
    .a(_0504_),
    .b(_0506_),
    .c(_0507_)
  );
  or_bb _2892_ (
    .a(_0507_),
    .b(_1140_),
    .c(_0508_)
  );
  or_bb _2893_ (
    .a(_0508_),
    .b(_0497_),
    .c(_0509_)
  );
  and_bb _2894_ (
    .a(_0338_),
    .b(_1140_),
    .c(_0511_)
  );
  or_bb _2895_ (
    .a(_0511_),
    .b(_1477_),
    .c(_0512_)
  );
  and_bi _2896_ (
    .a(_0509_),
    .b(_0512_),
    .c(_0513_)
  );
  or_bb _2897_ (
    .a(_0513_),
    .b(_0496_),
    .c(io_out_19_)
  );
  and_bi _2898_ (
    .a(io_adder_out_20_),
    .b(_1121_),
    .c(_0514_)
  );
  and_bi _2899_ (
    .a(_1336_),
    .b(_0333_),
    .c(_0515_)
  );
  and_bb _2900_ (
    .a(_1343_),
    .b(io_in2_20_),
    .c(_0516_)
  );
  or_bb _2901_ (
    .a(_0516_),
    .b(io_in1_20_),
    .c(_0517_)
  );
  and_bb _2902_ (
    .a(io_in2_20_),
    .b(io_in1_20_),
    .c(_0518_)
  );
  and_bb _2903_ (
    .a(_0518_),
    .b(_1341_),
    .c(_0519_)
  );
  and_bi _2904_ (
    .a(_0517_),
    .b(_0519_),
    .c(_0520_)
  );
  or_bb _2905_ (
    .a(_0520_),
    .b(_1345_),
    .c(_0521_)
  );
  and_bi _2906_ (
    .a(_1345_),
    .b(_0518_),
    .c(_0522_)
  );
  or_bb _2907_ (
    .a(_0522_),
    .b(_1336_),
    .c(_0523_)
  );
  and_bi _2908_ (
    .a(_0521_),
    .b(_0523_),
    .c(_0524_)
  );
  or_bb _2909_ (
    .a(_0524_),
    .b(_1140_),
    .c(_0525_)
  );
  or_bb _2910_ (
    .a(_0525_),
    .b(_0515_),
    .c(_0526_)
  );
  and_bb _2911_ (
    .a(_0316_),
    .b(_1140_),
    .c(_0527_)
  );
  or_bb _2912_ (
    .a(_0527_),
    .b(_1477_),
    .c(_0528_)
  );
  and_bi _2913_ (
    .a(_0526_),
    .b(_0528_),
    .c(_0529_)
  );
  or_bb _2914_ (
    .a(_0529_),
    .b(_0514_),
    .c(io_out_20_)
  );
  and_bi _2915_ (
    .a(io_adder_out_21_),
    .b(_1121_),
    .c(_0532_)
  );
  and_bi _2916_ (
    .a(_1336_),
    .b(_0310_),
    .c(_0533_)
  );
  and_bi _2917_ (
    .a(_1343_),
    .b(_0936_),
    .c(_0534_)
  );
  or_bb _2918_ (
    .a(_0534_),
    .b(io_in1_21_),
    .c(_0535_)
  );
  and_bb _2919_ (
    .a(io_in2_21_),
    .b(io_in1_21_),
    .c(_0536_)
  );
  and_bb _2920_ (
    .a(_0536_),
    .b(_1341_),
    .c(_0537_)
  );
  and_bi _2921_ (
    .a(_0535_),
    .b(_0537_),
    .c(_0538_)
  );
  or_bb _2922_ (
    .a(_0538_),
    .b(_1345_),
    .c(_0539_)
  );
  and_bi _2923_ (
    .a(_1345_),
    .b(_0536_),
    .c(_0540_)
  );
  or_bb _2924_ (
    .a(_0540_),
    .b(_1336_),
    .c(_0542_)
  );
  and_bi _2925_ (
    .a(_0539_),
    .b(_0542_),
    .c(_0543_)
  );
  or_bb _2926_ (
    .a(_0543_),
    .b(_1140_),
    .c(_0544_)
  );
  or_bb _2927_ (
    .a(_0544_),
    .b(_0533_),
    .c(_0545_)
  );
  and_bb _2928_ (
    .a(_0292_),
    .b(_1140_),
    .c(_0546_)
  );
  or_bb _2929_ (
    .a(_0546_),
    .b(_1477_),
    .c(_0547_)
  );
  and_bi _2930_ (
    .a(_0545_),
    .b(_0547_),
    .c(_0548_)
  );
  or_bb _2931_ (
    .a(_0548_),
    .b(_0532_),
    .c(io_out_21_)
  );
  and_bi _2932_ (
    .a(io_adder_out_22_),
    .b(_1121_),
    .c(_0549_)
  );
  and_bi _2933_ (
    .a(_1336_),
    .b(_0286_),
    .c(_0550_)
  );
  or_bb _2934_ (
    .a(_1345_),
    .b(_0945_),
    .c(_0552_)
  );
  inv _2935_ (
    .din(io_in2_22_),
    .dout(_0553_)
  );
  and_bi _2936_ (
    .a(_0945_),
    .b(_1343_),
    .c(_0554_)
  );
  or_bb _2937_ (
    .a(_0554_),
    .b(_0553_),
    .c(_0555_)
  );
  or_ii _2938_ (
    .a(_0555_),
    .b(_0552_),
    .c(_0556_)
  );
  and_bi _2939_ (
    .a(_1341_),
    .b(_0553_),
    .c(_0557_)
  );
  and_bi _2940_ (
    .a(_0557_),
    .b(_0552_),
    .c(_0558_)
  );
  or_bb _2941_ (
    .a(_0558_),
    .b(_1336_),
    .c(_0559_)
  );
  and_bi _2942_ (
    .a(_0556_),
    .b(_0559_),
    .c(_0560_)
  );
  or_bb _2943_ (
    .a(_0560_),
    .b(_1140_),
    .c(_0561_)
  );
  or_bb _2944_ (
    .a(_0561_),
    .b(_0550_),
    .c(_0562_)
  );
  and_bb _2945_ (
    .a(_0269_),
    .b(_1140_),
    .c(_0563_)
  );
  or_bb _2946_ (
    .a(_0563_),
    .b(_1477_),
    .c(_0564_)
  );
  and_bi _2947_ (
    .a(_0562_),
    .b(_0564_),
    .c(_0565_)
  );
  or_bb _2948_ (
    .a(_0565_),
    .b(_0549_),
    .c(io_out_22_)
  );
  and_bi _2949_ (
    .a(io_adder_out_23_),
    .b(_1121_),
    .c(_0566_)
  );
  and_bi _2950_ (
    .a(_0263_),
    .b(_1337_),
    .c(_0567_)
  );
  and_bi _2951_ (
    .a(_1343_),
    .b(_0955_),
    .c(_0568_)
  );
  or_bb _2952_ (
    .a(_0568_),
    .b(io_in1_23_),
    .c(_0569_)
  );
  and_bb _2953_ (
    .a(io_in2_23_),
    .b(io_in1_23_),
    .c(_0570_)
  );
  and_bb _2954_ (
    .a(_0570_),
    .b(_1341_),
    .c(_0573_)
  );
  and_bi _2955_ (
    .a(_0569_),
    .b(_0573_),
    .c(_0574_)
  );
  or_bb _2956_ (
    .a(_0574_),
    .b(_1345_),
    .c(_0575_)
  );
  and_bi _2957_ (
    .a(_1345_),
    .b(_0570_),
    .c(_0576_)
  );
  or_bb _2958_ (
    .a(_0576_),
    .b(_1336_),
    .c(_0577_)
  );
  and_bi _2959_ (
    .a(_0575_),
    .b(_0577_),
    .c(_0578_)
  );
  or_bb _2960_ (
    .a(_0578_),
    .b(_1140_),
    .c(_0579_)
  );
  or_bb _2961_ (
    .a(_0579_),
    .b(_0567_),
    .c(_0580_)
  );
  and_bb _2962_ (
    .a(_0246_),
    .b(_1140_),
    .c(_0581_)
  );
  or_bb _2963_ (
    .a(_0581_),
    .b(_1477_),
    .c(_0582_)
  );
  and_bi _2964_ (
    .a(_0580_),
    .b(_0582_),
    .c(_0584_)
  );
  or_bb _2965_ (
    .a(_0584_),
    .b(_0566_),
    .c(io_out_23_)
  );
  and_bi _2966_ (
    .a(_1336_),
    .b(_0240_),
    .c(_0585_)
  );
  and_bb _2967_ (
    .a(_1343_),
    .b(io_in2_24_),
    .c(_0586_)
  );
  or_bb _2968_ (
    .a(_0586_),
    .b(io_in1_24_),
    .c(_0587_)
  );
  and_bb _2969_ (
    .a(io_in2_24_),
    .b(io_in1_24_),
    .c(_0588_)
  );
  and_bb _2970_ (
    .a(_0588_),
    .b(_1341_),
    .c(_0589_)
  );
  and_bi _2971_ (
    .a(_0587_),
    .b(_0589_),
    .c(_0590_)
  );
  or_bb _2972_ (
    .a(_0590_),
    .b(_1345_),
    .c(_0591_)
  );
  and_bi _2973_ (
    .a(_1345_),
    .b(_0588_),
    .c(_0592_)
  );
  or_bb _2974_ (
    .a(_0592_),
    .b(_1336_),
    .c(_0594_)
  );
  and_bi _2975_ (
    .a(_0591_),
    .b(_0594_),
    .c(_0595_)
  );
  or_bb _2976_ (
    .a(_0595_),
    .b(_1140_),
    .c(_0596_)
  );
  or_bb _2977_ (
    .a(_0596_),
    .b(_0585_),
    .c(_0597_)
  );
  and_bb _2978_ (
    .a(_0209_),
    .b(_1140_),
    .c(_0598_)
  );
  or_bb _2979_ (
    .a(_0598_),
    .b(_1477_),
    .c(_0599_)
  );
  and_bi _2980_ (
    .a(_0597_),
    .b(_0599_),
    .c(_0600_)
  );
  and_bi _2981_ (
    .a(io_adder_out_24_),
    .b(_1121_),
    .c(_0601_)
  );
  or_bb _2982_ (
    .a(_0601_),
    .b(_0600_),
    .c(io_out_24_)
  );
  and_bi _2983_ (
    .a(io_adder_out_25_),
    .b(_1121_),
    .c(_0602_)
  );
  and_bi _2984_ (
    .a(_0201_),
    .b(_1337_),
    .c(_0604_)
  );
  and_bb _2985_ (
    .a(_1343_),
    .b(io_in2_25_),
    .c(_0605_)
  );
  or_bb _2986_ (
    .a(_0605_),
    .b(io_in1_25_),
    .c(_0606_)
  );
  and_bb _2987_ (
    .a(io_in2_25_),
    .b(io_in1_25_),
    .c(_0607_)
  );
  and_bb _2988_ (
    .a(_0607_),
    .b(_1341_),
    .c(_0608_)
  );
  and_bi _2989_ (
    .a(_0606_),
    .b(_0608_),
    .c(_0609_)
  );
  or_bb _2990_ (
    .a(_0609_),
    .b(_1345_),
    .c(_0610_)
  );
  and_bi _2991_ (
    .a(_1345_),
    .b(_0607_),
    .c(_0611_)
  );
  or_bb _2992_ (
    .a(_0611_),
    .b(_1336_),
    .c(_0612_)
  );
  and_bi _2993_ (
    .a(_0610_),
    .b(_0612_),
    .c(_0613_)
  );
  or_bb _2994_ (
    .a(_0613_),
    .b(_1140_),
    .c(_0614_)
  );
  or_bb _2995_ (
    .a(_0614_),
    .b(_0604_),
    .c(_0615_)
  );
  and_bb _2996_ (
    .a(_0171_),
    .b(_1140_),
    .c(_0616_)
  );
  or_bb _2997_ (
    .a(_0616_),
    .b(_1477_),
    .c(_0617_)
  );
  and_bi _2998_ (
    .a(_0615_),
    .b(_0617_),
    .c(_0618_)
  );
  or_bb _2999_ (
    .a(_0618_),
    .b(_0602_),
    .c(io_out_25_)
  );
  and_bi _3000_ (
    .a(io_adder_out_26_),
    .b(_1121_),
    .c(_0619_)
  );
  and_bi _3001_ (
    .a(_0163_),
    .b(_1337_),
    .c(_0620_)
  );
  or_bb _3002_ (
    .a(_1345_),
    .b(_0735_),
    .c(_0621_)
  );
  inv _3003_ (
    .din(io_in2_26_),
    .dout(_0622_)
  );
  and_bi _3004_ (
    .a(_0735_),
    .b(_1343_),
    .c(_0625_)
  );
  or_bb _3005_ (
    .a(_0625_),
    .b(_0622_),
    .c(_0626_)
  );
  or_ii _3006_ (
    .a(_0626_),
    .b(_0621_),
    .c(_0627_)
  );
  and_bi _3007_ (
    .a(_1341_),
    .b(_0622_),
    .c(_0628_)
  );
  and_bi _3008_ (
    .a(_0628_),
    .b(_0621_),
    .c(_0629_)
  );
  or_bb _3009_ (
    .a(_0629_),
    .b(_1336_),
    .c(_0630_)
  );
  and_bi _3010_ (
    .a(_0627_),
    .b(_0630_),
    .c(_0631_)
  );
  or_bb _3011_ (
    .a(_0631_),
    .b(_1140_),
    .c(_0632_)
  );
  or_bb _3012_ (
    .a(_0632_),
    .b(_0620_),
    .c(_0633_)
  );
  and_bb _3013_ (
    .a(_0134_),
    .b(_1140_),
    .c(_0634_)
  );
  or_bb _3014_ (
    .a(_0634_),
    .b(_1477_),
    .c(_0636_)
  );
  and_bi _3015_ (
    .a(_0633_),
    .b(_0636_),
    .c(_0637_)
  );
  or_bb _3016_ (
    .a(_0637_),
    .b(_0619_),
    .c(io_out_26_)
  );
  and_bi _3017_ (
    .a(io_adder_out_27_),
    .b(_1121_),
    .c(_0638_)
  );
  and_bi _3018_ (
    .a(_1336_),
    .b(_0126_),
    .c(_0639_)
  );
  and_bb _3019_ (
    .a(_1343_),
    .b(io_in2_27_),
    .c(_0640_)
  );
  or_bb _3020_ (
    .a(_0640_),
    .b(io_in1_27_),
    .c(_0641_)
  );
  and_bb _3021_ (
    .a(io_in2_27_),
    .b(io_in1_27_),
    .c(_0642_)
  );
  and_bb _3022_ (
    .a(_0642_),
    .b(_1341_),
    .c(_0643_)
  );
  and_bi _3023_ (
    .a(_0641_),
    .b(_0643_),
    .c(_0644_)
  );
  or_bb _3024_ (
    .a(_0644_),
    .b(_1345_),
    .c(_0646_)
  );
  and_bi _3025_ (
    .a(_1345_),
    .b(_0642_),
    .c(_0647_)
  );
  or_bb _3026_ (
    .a(_0647_),
    .b(_1336_),
    .c(_0648_)
  );
  and_bi _3027_ (
    .a(_0646_),
    .b(_0648_),
    .c(_0649_)
  );
  or_bb _3028_ (
    .a(_0649_),
    .b(_1140_),
    .c(_0650_)
  );
  or_bb _3029_ (
    .a(_0650_),
    .b(_0639_),
    .c(_0651_)
  );
  and_bb _3030_ (
    .a(_0096_),
    .b(_1140_),
    .c(_0652_)
  );
  or_bb _3031_ (
    .a(_0652_),
    .b(_1477_),
    .c(_0653_)
  );
  and_bi _3032_ (
    .a(_0651_),
    .b(_0653_),
    .c(_0654_)
  );
  or_bb _3033_ (
    .a(_0654_),
    .b(_0638_),
    .c(io_out_27_)
  );
  and_bi _3034_ (
    .a(io_adder_out_28_),
    .b(_1121_),
    .c(_0655_)
  );
  and_bi _3035_ (
    .a(_0088_),
    .b(_1337_),
    .c(_0656_)
  );
  and_bb _3036_ (
    .a(_1343_),
    .b(io_in2_28_),
    .c(_0657_)
  );
  or_bb _3037_ (
    .a(_0657_),
    .b(io_in1_28_),
    .c(_0658_)
  );
  and_bb _3038_ (
    .a(io_in2_28_),
    .b(io_in1_28_),
    .c(_0659_)
  );
  and_bb _3039_ (
    .a(_0659_),
    .b(_1341_),
    .c(_0660_)
  );
  and_bi _3040_ (
    .a(_0658_),
    .b(_0660_),
    .c(_0661_)
  );
  or_bb _3041_ (
    .a(_0661_),
    .b(_1345_),
    .c(_0662_)
  );
  and_bi _3042_ (
    .a(_1345_),
    .b(_0659_),
    .c(_0663_)
  );
  or_bb _3043_ (
    .a(_0663_),
    .b(_1336_),
    .c(_0664_)
  );
  and_bi _3044_ (
    .a(_0662_),
    .b(_0664_),
    .c(_0667_)
  );
  or_bb _3045_ (
    .a(_0667_),
    .b(_1140_),
    .c(_0668_)
  );
  or_bb _3046_ (
    .a(_0668_),
    .b(_0656_),
    .c(_0669_)
  );
  and_bb _3047_ (
    .a(_0032_),
    .b(_1140_),
    .c(_0670_)
  );
  or_bb _3048_ (
    .a(_0670_),
    .b(_1477_),
    .c(_0671_)
  );
  and_bi _3049_ (
    .a(_0669_),
    .b(_0671_),
    .c(_0672_)
  );
  or_bb _3050_ (
    .a(_0672_),
    .b(_0655_),
    .c(io_out_28_)
  );
  and_bi _3051_ (
    .a(_1336_),
    .b(_0022_),
    .c(_0673_)
  );
  and_bi _3052_ (
    .a(_1343_),
    .b(_0363_),
    .c(_0674_)
  );
  or_bb _3053_ (
    .a(_0674_),
    .b(io_in1_29_),
    .c(_0675_)
  );
  and_bb _3054_ (
    .a(io_in2_29_),
    .b(io_in1_29_),
    .c(_0677_)
  );
  and_bb _3055_ (
    .a(_0677_),
    .b(_1341_),
    .c(_0678_)
  );
  and_bi _3056_ (
    .a(_0675_),
    .b(_0678_),
    .c(_0679_)
  );
  or_bb _3057_ (
    .a(_0679_),
    .b(_1345_),
    .c(_0680_)
  );
  and_bi _3058_ (
    .a(_1345_),
    .b(_0677_),
    .c(_0681_)
  );
  or_bb _3059_ (
    .a(_0681_),
    .b(_1336_),
    .c(_0682_)
  );
  and_bi _3060_ (
    .a(_0680_),
    .b(_0682_),
    .c(_0683_)
  );
  or_bb _3061_ (
    .a(_0683_),
    .b(_1140_),
    .c(_0684_)
  );
  or_bb _3062_ (
    .a(_0684_),
    .b(_0673_),
    .c(_0685_)
  );
  and_bb _3063_ (
    .a(_1486_),
    .b(_1140_),
    .c(_0686_)
  );
  or_bb _3064_ (
    .a(_0686_),
    .b(_1477_),
    .c(_0688_)
  );
  and_bi _3065_ (
    .a(_0685_),
    .b(_0688_),
    .c(_0689_)
  );
  and_bi _3066_ (
    .a(io_adder_out_29_),
    .b(_1121_),
    .c(_0690_)
  );
  or_bb _3067_ (
    .a(_0690_),
    .b(_0689_),
    .c(io_out_29_)
  );
  and_bi _3068_ (
    .a(io_adder_out_30_),
    .b(_1121_),
    .c(_0691_)
  );
  and_bi _3069_ (
    .a(_1475_),
    .b(_1337_),
    .c(_0692_)
  );
  and_bi _3070_ (
    .a(_0733_),
    .b(_1343_),
    .c(_0693_)
  );
  inv _3071_ (
    .din(io_in2_30_),
    .dout(_0694_)
  );
  and_bi _3072_ (
    .a(io_in1_30_),
    .b(_1345_),
    .c(_0695_)
  );
  or_bb _3073_ (
    .a(_0695_),
    .b(_0694_),
    .c(_0696_)
  );
  or_bb _3074_ (
    .a(_0696_),
    .b(_0693_),
    .c(_0698_)
  );
  and_bi _3075_ (
    .a(_1341_),
    .b(_0694_),
    .c(_0699_)
  );
  and_bi _3076_ (
    .a(_0695_),
    .b(_0699_),
    .c(_0700_)
  );
  and_bi _3077_ (
    .a(_0698_),
    .b(_0700_),
    .c(_0701_)
  );
  and_bi _3078_ (
    .a(_1337_),
    .b(_0701_),
    .c(_0702_)
  );
  or_bb _3079_ (
    .a(_0702_),
    .b(_1140_),
    .c(_0703_)
  );
  or_bb _3080_ (
    .a(_0703_),
    .b(_0692_),
    .c(_0704_)
  );
  and_bb _3081_ (
    .a(_1373_),
    .b(_1140_),
    .c(_0705_)
  );
  or_bb _3082_ (
    .a(_0705_),
    .b(_1477_),
    .c(_0706_)
  );
  and_bi _3083_ (
    .a(_0704_),
    .b(_0706_),
    .c(_0707_)
  );
  or_bb _3084_ (
    .a(_0707_),
    .b(_0691_),
    .c(io_out_30_)
  );
  and_bi _3085_ (
    .a(io_adder_out_31_),
    .b(_1121_),
    .c(_0708_)
  );
  and_bi _3086_ (
    .a(_1334_),
    .b(_1337_),
    .c(_0709_)
  );
  and_bb _3087_ (
    .a(io_in2_31_),
    .b(io_in1_31_),
    .c(_0710_)
  );
  and_bi _3088_ (
    .a(_1345_),
    .b(_0710_),
    .c(_0711_)
  );
  and_bi _3089_ (
    .a(_1337_),
    .b(_0711_),
    .c(_0712_)
  );
  or_bb _3090_ (
    .a(_1341_),
    .b(_0340_),
    .c(_0713_)
  );
  and_bb _3091_ (
    .a(_1343_),
    .b(_1125_),
    .c(_0714_)
  );
  or_bb _3092_ (
    .a(_0714_),
    .b(_1124_),
    .c(_0715_)
  );
  and_bi _3093_ (
    .a(_0713_),
    .b(_0715_),
    .c(_0716_)
  );
  and_bi _3094_ (
    .a(_0712_),
    .b(_0716_),
    .c(_0719_)
  );
  or_bb _3095_ (
    .a(_0719_),
    .b(_1140_),
    .c(_0720_)
  );
  or_bb _3096_ (
    .a(_0720_),
    .b(_0709_),
    .c(_0721_)
  );
  and_bb _3097_ (
    .a(_1339_),
    .b(_1140_),
    .c(_0722_)
  );
  or_bb _3098_ (
    .a(_0722_),
    .b(_1477_),
    .c(_0723_)
  );
  and_bi _3099_ (
    .a(_0721_),
    .b(_0723_),
    .c(_0724_)
  );
  or_bb _3100_ (
    .a(_0724_),
    .b(_0708_),
    .c(io_out_31_)
  );
endmodule
