module sorter32(a, b);
  input a_0_;
  input a_1_;
  input a_2_;
  input a_3_;
  input a_4_;
  input a_5_;
  input a_6_;
  input a_7_;
  input a_8_;
  input a_9_;
  input a_10_;
  input a_11_;
  input a_12_;
  input a_13_;
  input a_14_;
  input a_15_;
  input a_16_;
  input a_17_;
  input a_18_;
  input a_19_;
  input a_20_;
  input a_21_;
  input a_22_;
  input a_23_;
  input a_24_;
  input a_25_;
  input a_26_;
  input a_27_;
  input a_28_;
  input a_29_;
  input a_30_;
  input a_31_;
  output b_0_;
  output b_1_;
  output b_2_;
  output b_3_;
  output b_4_;
  output b_5_;
  output b_6_;
  output b_7_;
  output b_8_;
  output b_9_;
  output b_10_;
  output b_11_;
  output b_12_;
  output b_13_;
  output b_14_;
  output b_15_;
  output b_16_;
  output b_17_;
  output b_18_;
  output b_19_;
  output b_20_;
  output b_21_;
  output b_22_;
  output b_23_;
  output b_24_;
  output b_25_;
  output b_26_;
  output b_27_;
  output b_28_;
  output b_29_;
  output b_30_;
  output b_31_;
  wire c_0_;
  wire c_1_;
  wire c_2_;
  wire c_3_;
  wire c_4_;
  wire c_5_;
  wire c_6_;
  wire c_7_;
  wire c_8_;
  wire c_9_;
  wire c_10_;
  wire c_11_;
  wire c_12_;
  wire c_13_;
  wire c_14_;
  wire c_15_;
  wire c_16_;
  wire c_17_;
  wire c_18_;
  wire c_19_;
  wire c_20_;
  wire c_21_;
  wire c_22_;
  wire c_23_;
  wire c_24_;
  wire c_25_;
  wire c_26_;
  wire c_27_;
  wire c_28_;
  wire c_29_;
  wire c_30_;
  wire c_31_;
  wire _gdown_c_0_;
  wire _gdown_c_1_;
  wire _gdown_c_2_;
  wire _gdown_c_3_;
  wire _gdown_c_4_;
  wire _gdown_c_5_;
  wire _gdown_c_6_;
  wire _gdown_c_7_;
  wire _gdown_c_8_;
  wire _gdown_c_9_;
  wire _gdown_c_10_;
  wire _gdown_c_11_;
  wire _gdown_c_12_;
  wire _gdown_c_13_;
  wire _gdown_c_14_;
  wire _gdown_c_15_;
  wire _gdown_gdown_c_0_;
  wire _gdown_gdown_c_1_;
  wire _gdown_gdown_c_2_;
  wire _gdown_gdown_c_3_;
  wire _gdown_gdown_c_4_;
  wire _gdown_gdown_c_5_;
  wire _gdown_gdown_c_6_;
  wire _gdown_gdown_c_7_;
  wire _gdown_gdown_gdown_c_0_;
  wire _gdown_gdown_gdown_c_1_;
  wire _gdown_gdown_gdown_c_2_;
  wire _gdown_gdown_gdown_c_3_;
  wire _gdown_gdown_gdown_g_3_c_0_;
  wire _gdown_gdown_gdown_g_3_c_1_;
  wire _gdown_gdown_gdown_g_3_c_2_;
  wire _gdown_gdown_gdown_g_3_c_3_;
  wire _gdown_gdown_gup_c_0_;
  wire _gdown_gdown_gup_c_1_;
  wire _gdown_gdown_gup_c_2_;
  wire _gdown_gdown_gup_c_3_;
  wire _gdown_gdown_gup_g_3_c_0_;
  wire _gdown_gdown_gup_g_3_c_1_;
  wire _gdown_gdown_gup_g_3_c_2_;
  wire _gdown_gdown_gup_g_3_c_3_;
  wire _gdown_gdown_m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_;
  wire _gdown_gdown_m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_;
  wire _gdown_gdown_m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_;
  wire _gdown_gdown_m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_;
  wire _gdown_gdown_m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_;
  wire _gdown_gdown_m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_;
  wire _gdown_gdown_m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_;
  wire _gdown_gdown_m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_;
  wire _gdown_gdown_m_genblock__src_b32s_merger8_v_1333_0__m_c_0_;
  wire _gdown_gdown_m_genblock__src_b32s_merger8_v_1333_0__m_c_1_;
  wire _gdown_gdown_m_genblock__src_b32s_merger8_v_1333_0__m_c_2_;
  wire _gdown_gdown_m_genblock__src_b32s_merger8_v_1333_0__m_c_3_;
  wire _gdown_gdown_m_genblock__src_b32s_merger8_v_1334_1__m_c_0_;
  wire _gdown_gdown_m_genblock__src_b32s_merger8_v_1334_1__m_c_1_;
  wire _gdown_gdown_m_genblock__src_b32s_merger8_v_1334_1__m_c_2_;
  wire _gdown_gdown_m_genblock__src_b32s_merger8_v_1334_1__m_c_3_;
  wire _gdown_gup_c_0_;
  wire _gdown_gup_c_1_;
  wire _gdown_gup_c_2_;
  wire _gdown_gup_c_3_;
  wire _gdown_gup_c_4_;
  wire _gdown_gup_c_5_;
  wire _gdown_gup_c_6_;
  wire _gdown_gup_c_7_;
  wire _gdown_gup_gdown_c_0_;
  wire _gdown_gup_gdown_c_1_;
  wire _gdown_gup_gdown_c_2_;
  wire _gdown_gup_gdown_c_3_;
  wire _gdown_gup_gdown_g_3_c_0_;
  wire _gdown_gup_gdown_g_3_c_1_;
  wire _gdown_gup_gdown_g_3_c_2_;
  wire _gdown_gup_gdown_g_3_c_3_;
  wire _gdown_gup_gup_c_0_;
  wire _gdown_gup_gup_c_1_;
  wire _gdown_gup_gup_c_2_;
  wire _gdown_gup_gup_c_3_;
  wire _gdown_gup_gup_g_3_c_0_;
  wire _gdown_gup_gup_g_3_c_1_;
  wire _gdown_gup_gup_g_3_c_2_;
  wire _gdown_gup_gup_g_3_c_3_;
  wire _gdown_gup_m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_;
  wire _gdown_gup_m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_;
  wire _gdown_gup_m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_;
  wire _gdown_gup_m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_;
  wire _gdown_gup_m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_;
  wire _gdown_gup_m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_;
  wire _gdown_gup_m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_;
  wire _gdown_gup_m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_;
  wire _gdown_gup_m_genblock__src_b32s_merger8_v_1333_0__m_c_0_;
  wire _gdown_gup_m_genblock__src_b32s_merger8_v_1333_0__m_c_1_;
  wire _gdown_gup_m_genblock__src_b32s_merger8_v_1333_0__m_c_2_;
  wire _gdown_gup_m_genblock__src_b32s_merger8_v_1333_0__m_c_3_;
  wire _gdown_gup_m_genblock__src_b32s_merger8_v_1334_1__m_c_0_;
  wire _gdown_gup_m_genblock__src_b32s_merger8_v_1334_1__m_c_1_;
  wire _gdown_gup_m_genblock__src_b32s_merger8_v_1334_1__m_c_2_;
  wire _gdown_gup_m_genblock__src_b32s_merger8_v_1334_1__m_c_3_;
  wire _gdown_m_genblock__src_b32s_merger16_v_101_0__g_ord_0_;
  wire _gdown_m_genblock__src_b32s_merger16_v_101_0__g_ord_1_;
  wire _gdown_m_genblock__src_b32s_merger16_v_102_1__g_ord_0_;
  wire _gdown_m_genblock__src_b32s_merger16_v_102_1__g_ord_1_;
  wire _gdown_m_genblock__src_b32s_merger16_v_103_2__g_ord_0_;
  wire _gdown_m_genblock__src_b32s_merger16_v_103_2__g_ord_1_;
  wire _gdown_m_genblock__src_b32s_merger16_v_104_3__g_ord_0_;
  wire _gdown_m_genblock__src_b32s_merger16_v_104_3__g_ord_1_;
  wire _gdown_m_genblock__src_b32s_merger16_v_105_4__g_ord_0_;
  wire _gdown_m_genblock__src_b32s_merger16_v_105_4__g_ord_1_;
  wire _gdown_m_genblock__src_b32s_merger16_v_106_5__g_ord_0_;
  wire _gdown_m_genblock__src_b32s_merger16_v_106_5__g_ord_1_;
  wire _gdown_m_genblock__src_b32s_merger16_v_107_6__g_ord_0_;
  wire _gdown_m_genblock__src_b32s_merger16_v_107_6__g_ord_1_;
  wire _gdown_m_genblock__src_b32s_merger16_v_108_7__g_ord_0_;
  wire _gdown_m_genblock__src_b32s_merger16_v_108_7__g_ord_1_;
  wire _gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_;
  wire _gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_;
  wire _gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_;
  wire _gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_;
  wire _gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_;
  wire _gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_;
  wire _gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_;
  wire _gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_;
  wire _gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_0_;
  wire _gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_1_;
  wire _gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_2_;
  wire _gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_3_;
  wire _gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_0_;
  wire _gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_1_;
  wire _gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_2_;
  wire _gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_3_;
  wire _gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_;
  wire _gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_;
  wire _gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_;
  wire _gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_;
  wire _gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_;
  wire _gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_;
  wire _gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_;
  wire _gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_;
  wire _gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_0_;
  wire _gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_1_;
  wire _gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_2_;
  wire _gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_3_;
  wire _gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_0_;
  wire _gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_1_;
  wire _gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_2_;
  wire _gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_3_;
  wire _gup_c_0_;
  wire _gup_c_1_;
  wire _gup_c_2_;
  wire _gup_c_3_;
  wire _gup_c_4_;
  wire _gup_c_5_;
  wire _gup_c_6_;
  wire _gup_c_7_;
  wire _gup_c_8_;
  wire _gup_c_9_;
  wire _gup_c_10_;
  wire _gup_c_11_;
  wire _gup_c_12_;
  wire _gup_c_13_;
  wire _gup_c_14_;
  wire _gup_c_15_;
  wire _gup_gdown_c_0_;
  wire _gup_gdown_c_1_;
  wire _gup_gdown_c_2_;
  wire _gup_gdown_c_3_;
  wire _gup_gdown_c_4_;
  wire _gup_gdown_c_5_;
  wire _gup_gdown_c_6_;
  wire _gup_gdown_c_7_;
  wire _gup_gdown_gdown_c_0_;
  wire _gup_gdown_gdown_c_1_;
  wire _gup_gdown_gdown_c_2_;
  wire _gup_gdown_gdown_c_3_;
  wire _gup_gdown_gdown_g_3_c_0_;
  wire _gup_gdown_gdown_g_3_c_1_;
  wire _gup_gdown_gdown_g_3_c_2_;
  wire _gup_gdown_gdown_g_3_c_3_;
  wire _gup_gdown_gup_c_0_;
  wire _gup_gdown_gup_c_1_;
  wire _gup_gdown_gup_c_2_;
  wire _gup_gdown_gup_c_3_;
  wire _gup_gdown_gup_g_3_c_0_;
  wire _gup_gdown_gup_g_3_c_1_;
  wire _gup_gdown_gup_g_3_c_2_;
  wire _gup_gdown_gup_g_3_c_3_;
  wire _gup_gdown_m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_;
  wire _gup_gdown_m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_;
  wire _gup_gdown_m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_;
  wire _gup_gdown_m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_;
  wire _gup_gdown_m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_;
  wire _gup_gdown_m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_;
  wire _gup_gdown_m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_;
  wire _gup_gdown_m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_;
  wire _gup_gdown_m_genblock__src_b32s_merger8_v_1333_0__m_c_0_;
  wire _gup_gdown_m_genblock__src_b32s_merger8_v_1333_0__m_c_1_;
  wire _gup_gdown_m_genblock__src_b32s_merger8_v_1333_0__m_c_2_;
  wire _gup_gdown_m_genblock__src_b32s_merger8_v_1333_0__m_c_3_;
  wire _gup_gdown_m_genblock__src_b32s_merger8_v_1334_1__m_c_0_;
  wire _gup_gdown_m_genblock__src_b32s_merger8_v_1334_1__m_c_1_;
  wire _gup_gdown_m_genblock__src_b32s_merger8_v_1334_1__m_c_2_;
  wire _gup_gdown_m_genblock__src_b32s_merger8_v_1334_1__m_c_3_;
  wire _gup_gup_c_0_;
  wire _gup_gup_c_1_;
  wire _gup_gup_c_2_;
  wire _gup_gup_c_3_;
  wire _gup_gup_c_4_;
  wire _gup_gup_c_5_;
  wire _gup_gup_c_6_;
  wire _gup_gup_c_7_;
  wire _gup_gup_gdown_c_0_;
  wire _gup_gup_gdown_c_1_;
  wire _gup_gup_gdown_c_2_;
  wire _gup_gup_gdown_c_3_;
  wire _gup_gup_gdown_g_3_c_0_;
  wire _gup_gup_gdown_g_3_c_1_;
  wire _gup_gup_gdown_g_3_c_2_;
  wire _gup_gup_gdown_g_3_c_3_;
  wire _gup_gup_gup_c_0_;
  wire _gup_gup_gup_c_1_;
  wire _gup_gup_gup_c_2_;
  wire _gup_gup_gup_c_3_;
  wire _gup_gup_gup_g_3_c_0_;
  wire _gup_gup_gup_g_3_c_1_;
  wire _gup_gup_gup_g_3_c_2_;
  wire _gup_gup_gup_g_3_c_3_;
  wire _gup_gup_m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_;
  wire _gup_gup_m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_;
  wire _gup_gup_m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_;
  wire _gup_gup_m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_;
  wire _gup_gup_m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_;
  wire _gup_gup_m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_;
  wire _gup_gup_m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_;
  wire _gup_gup_m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_;
  wire _gup_gup_m_genblock__src_b32s_merger8_v_1333_0__m_c_0_;
  wire _gup_gup_m_genblock__src_b32s_merger8_v_1333_0__m_c_1_;
  wire _gup_gup_m_genblock__src_b32s_merger8_v_1333_0__m_c_2_;
  wire _gup_gup_m_genblock__src_b32s_merger8_v_1333_0__m_c_3_;
  wire _gup_gup_m_genblock__src_b32s_merger8_v_1334_1__m_c_0_;
  wire _gup_gup_m_genblock__src_b32s_merger8_v_1334_1__m_c_1_;
  wire _gup_gup_m_genblock__src_b32s_merger8_v_1334_1__m_c_2_;
  wire _gup_gup_m_genblock__src_b32s_merger8_v_1334_1__m_c_3_;
  wire _gup_m_genblock__src_b32s_merger16_v_101_0__g_ord_0_;
  wire _gup_m_genblock__src_b32s_merger16_v_101_0__g_ord_1_;
  wire _gup_m_genblock__src_b32s_merger16_v_102_1__g_ord_0_;
  wire _gup_m_genblock__src_b32s_merger16_v_102_1__g_ord_1_;
  wire _gup_m_genblock__src_b32s_merger16_v_103_2__g_ord_0_;
  wire _gup_m_genblock__src_b32s_merger16_v_103_2__g_ord_1_;
  wire _gup_m_genblock__src_b32s_merger16_v_104_3__g_ord_0_;
  wire _gup_m_genblock__src_b32s_merger16_v_104_3__g_ord_1_;
  wire _gup_m_genblock__src_b32s_merger16_v_105_4__g_ord_0_;
  wire _gup_m_genblock__src_b32s_merger16_v_105_4__g_ord_1_;
  wire _gup_m_genblock__src_b32s_merger16_v_106_5__g_ord_0_;
  wire _gup_m_genblock__src_b32s_merger16_v_106_5__g_ord_1_;
  wire _gup_m_genblock__src_b32s_merger16_v_107_6__g_ord_0_;
  wire _gup_m_genblock__src_b32s_merger16_v_107_6__g_ord_1_;
  wire _gup_m_genblock__src_b32s_merger16_v_108_7__g_ord_0_;
  wire _gup_m_genblock__src_b32s_merger16_v_108_7__g_ord_1_;
  wire _gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_;
  wire _gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_;
  wire _gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_;
  wire _gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_;
  wire _gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_;
  wire _gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_;
  wire _gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_;
  wire _gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_;
  wire _gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_0_;
  wire _gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_1_;
  wire _gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_2_;
  wire _gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_3_;
  wire _gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_0_;
  wire _gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_1_;
  wire _gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_2_;
  wire _gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_3_;
  wire _gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_;
  wire _gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_;
  wire _gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_;
  wire _gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_;
  wire _gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_;
  wire _gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_;
  wire _gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_;
  wire _gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_;
  wire _gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_0_;
  wire _gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_1_;
  wire _gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_2_;
  wire _gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_3_;
  wire _gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_0_;
  wire _gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_1_;
  wire _gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_2_;
  wire _gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_3_;
  wire _m_genblock__src_b32s_merger32_v_1011_0__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1011_0__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1012_1__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1012_1__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1013_2__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1013_2__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1014_3__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1014_3__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1015_4__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1015_4__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1016_5__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1016_5__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1017_6__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1017_6__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1018_7__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1018_7__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1019_8__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1019_8__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1020_9__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1020_9__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1021_10__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1021_10__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1022_11__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1022_11__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1023_12__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1023_12__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1024_13__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1024_13__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1025_14__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1025_14__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1026_15__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1026_15__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_101_0__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_101_0__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_102_1__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_102_1__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_103_2__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_103_2__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_104_3__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_104_3__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_105_4__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_105_4__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_106_5__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_106_5__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_107_6__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_107_6__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_108_7__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_108_7__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_0_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_1_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_2_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_3_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_0_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_1_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_2_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_3_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_0_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_1_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_2_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_3_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_0_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_1_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_2_;
  wire _m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_3_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_101_0__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_101_0__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_102_1__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_102_1__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_103_2__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_103_2__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_104_3__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_104_3__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_105_4__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_105_4__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_106_5__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_106_5__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_107_6__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_107_6__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_108_7__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_108_7__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_0_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_1_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_2_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_3_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_0_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_1_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_2_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_3_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_0_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_1_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_2_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_3_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_0_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_1_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_2_;
  wire _m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_3_;
  or_bb _000_ (
    .a(a_30_),
    .b(a_31_),
    .c(_gdown_gdown_gdown_c_3_)
  );
  and_bb _001_ (
    .a(a_30_),
    .b(a_31_),
    .c(_gdown_gdown_gdown_c_2_)
  );
  or_bb _002_ (
    .a(a_28_),
    .b(a_29_),
    .c(_gdown_gdown_gdown_c_0_)
  );
  and_bb _003_ (
    .a(a_28_),
    .b(a_29_),
    .c(_gdown_gdown_gdown_c_1_)
  );
  or_bb _004_ (
    .a(_gdown_gdown_gdown_c_1_),
    .b(_gdown_gdown_gdown_c_3_),
    .c(_gdown_gdown_gdown_g_3_c_3_)
  );
  and_bb _005_ (
    .a(_gdown_gdown_gdown_c_1_),
    .b(_gdown_gdown_gdown_c_3_),
    .c(_gdown_gdown_gdown_g_3_c_1_)
  );
  or_bb _006_ (
    .a(_gdown_gdown_gdown_c_0_),
    .b(_gdown_gdown_gdown_c_2_),
    .c(_gdown_gdown_gdown_g_3_c_2_)
  );
  and_bb _007_ (
    .a(_gdown_gdown_gdown_c_0_),
    .b(_gdown_gdown_gdown_c_2_),
    .c(_gdown_gdown_gdown_g_3_c_0_)
  );
  or_bb _008_ (
    .a(_gdown_gdown_gdown_g_3_c_2_),
    .b(_gdown_gdown_gdown_g_3_c_3_),
    .c(_gdown_gdown_c_7_)
  );
  and_bb _009_ (
    .a(_gdown_gdown_gdown_g_3_c_2_),
    .b(_gdown_gdown_gdown_g_3_c_3_),
    .c(_gdown_gdown_c_6_)
  );
  or_bb _010_ (
    .a(_gdown_gdown_gdown_g_3_c_0_),
    .b(_gdown_gdown_gdown_g_3_c_1_),
    .c(_gdown_gdown_c_5_)
  );
  and_bb _011_ (
    .a(_gdown_gdown_gdown_g_3_c_0_),
    .b(_gdown_gdown_gdown_g_3_c_1_),
    .c(_gdown_gdown_c_4_)
  );
  or_bb _012_ (
    .a(a_26_),
    .b(a_27_),
    .c(_gdown_gdown_gup_c_3_)
  );
  and_bb _013_ (
    .a(a_26_),
    .b(a_27_),
    .c(_gdown_gdown_gup_c_2_)
  );
  or_bb _014_ (
    .a(a_24_),
    .b(a_25_),
    .c(_gdown_gdown_gup_c_0_)
  );
  and_bb _015_ (
    .a(a_24_),
    .b(a_25_),
    .c(_gdown_gdown_gup_c_1_)
  );
  or_bb _016_ (
    .a(_gdown_gdown_gup_c_1_),
    .b(_gdown_gdown_gup_c_3_),
    .c(_gdown_gdown_gup_g_3_c_3_)
  );
  and_bb _017_ (
    .a(_gdown_gdown_gup_c_1_),
    .b(_gdown_gdown_gup_c_3_),
    .c(_gdown_gdown_gup_g_3_c_1_)
  );
  or_bb _018_ (
    .a(_gdown_gdown_gup_c_0_),
    .b(_gdown_gdown_gup_c_2_),
    .c(_gdown_gdown_gup_g_3_c_2_)
  );
  and_bb _019_ (
    .a(_gdown_gdown_gup_c_0_),
    .b(_gdown_gdown_gup_c_2_),
    .c(_gdown_gdown_gup_g_3_c_0_)
  );
  or_bb _020_ (
    .a(_gdown_gdown_gup_g_3_c_2_),
    .b(_gdown_gdown_gup_g_3_c_3_),
    .c(_gdown_gdown_c_0_)
  );
  and_bb _021_ (
    .a(_gdown_gdown_gup_g_3_c_2_),
    .b(_gdown_gdown_gup_g_3_c_3_),
    .c(_gdown_gdown_c_1_)
  );
  or_bb _022_ (
    .a(_gdown_gdown_gup_g_3_c_0_),
    .b(_gdown_gdown_gup_g_3_c_1_),
    .c(_gdown_gdown_c_2_)
  );
  and_bb _023_ (
    .a(_gdown_gdown_gup_g_3_c_0_),
    .b(_gdown_gdown_gup_g_3_c_1_),
    .c(_gdown_gdown_c_3_)
  );
  or_bb _024_ (
    .a(_gdown_gdown_c_0_),
    .b(_gdown_gdown_c_4_),
    .c(_gdown_gdown_m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_)
  );
  and_bb _025_ (
    .a(_gdown_gdown_c_0_),
    .b(_gdown_gdown_c_4_),
    .c(_gdown_gdown_m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_)
  );
  or_bb _026_ (
    .a(_gdown_gdown_c_1_),
    .b(_gdown_gdown_c_5_),
    .c(_gdown_gdown_m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_)
  );
  and_bb _027_ (
    .a(_gdown_gdown_c_1_),
    .b(_gdown_gdown_c_5_),
    .c(_gdown_gdown_m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_)
  );
  or_bb _028_ (
    .a(_gdown_gdown_c_2_),
    .b(_gdown_gdown_c_6_),
    .c(_gdown_gdown_m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_)
  );
  and_bb _029_ (
    .a(_gdown_gdown_c_2_),
    .b(_gdown_gdown_c_6_),
    .c(_gdown_gdown_m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_)
  );
  or_bb _030_ (
    .a(_gdown_gdown_c_3_),
    .b(_gdown_gdown_c_7_),
    .c(_gdown_gdown_m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_)
  );
  and_bb _031_ (
    .a(_gdown_gdown_c_3_),
    .b(_gdown_gdown_c_7_),
    .c(_gdown_gdown_m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_)
  );
  or_bb _032_ (
    .a(_gdown_gdown_m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_),
    .b(_gdown_gdown_m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_),
    .c(_gdown_gdown_m_genblock__src_b32s_merger8_v_1333_0__m_c_3_)
  );
  and_bb _033_ (
    .a(_gdown_gdown_m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_),
    .b(_gdown_gdown_m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_),
    .c(_gdown_gdown_m_genblock__src_b32s_merger8_v_1333_0__m_c_1_)
  );
  or_bb _034_ (
    .a(_gdown_gdown_m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_),
    .b(_gdown_gdown_m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_),
    .c(_gdown_gdown_m_genblock__src_b32s_merger8_v_1333_0__m_c_2_)
  );
  and_bb _035_ (
    .a(_gdown_gdown_m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_),
    .b(_gdown_gdown_m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_),
    .c(_gdown_gdown_m_genblock__src_b32s_merger8_v_1333_0__m_c_0_)
  );
  or_bb _036_ (
    .a(_gdown_gdown_m_genblock__src_b32s_merger8_v_1333_0__m_c_2_),
    .b(_gdown_gdown_m_genblock__src_b32s_merger8_v_1333_0__m_c_3_),
    .c(_gdown_c_11_)
  );
  and_bb _037_ (
    .a(_gdown_gdown_m_genblock__src_b32s_merger8_v_1333_0__m_c_2_),
    .b(_gdown_gdown_m_genblock__src_b32s_merger8_v_1333_0__m_c_3_),
    .c(_gdown_c_10_)
  );
  or_bb _038_ (
    .a(_gdown_gdown_m_genblock__src_b32s_merger8_v_1333_0__m_c_0_),
    .b(_gdown_gdown_m_genblock__src_b32s_merger8_v_1333_0__m_c_1_),
    .c(_gdown_c_9_)
  );
  and_bb _039_ (
    .a(_gdown_gdown_m_genblock__src_b32s_merger8_v_1333_0__m_c_0_),
    .b(_gdown_gdown_m_genblock__src_b32s_merger8_v_1333_0__m_c_1_),
    .c(_gdown_c_8_)
  );
  or_bb _040_ (
    .a(_gdown_gdown_m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_),
    .b(_gdown_gdown_m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_),
    .c(_gdown_gdown_m_genblock__src_b32s_merger8_v_1334_1__m_c_3_)
  );
  and_bb _041_ (
    .a(_gdown_gdown_m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_),
    .b(_gdown_gdown_m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_),
    .c(_gdown_gdown_m_genblock__src_b32s_merger8_v_1334_1__m_c_1_)
  );
  or_bb _042_ (
    .a(_gdown_gdown_m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_),
    .b(_gdown_gdown_m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_),
    .c(_gdown_gdown_m_genblock__src_b32s_merger8_v_1334_1__m_c_2_)
  );
  and_bb _043_ (
    .a(_gdown_gdown_m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_),
    .b(_gdown_gdown_m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_),
    .c(_gdown_gdown_m_genblock__src_b32s_merger8_v_1334_1__m_c_0_)
  );
  or_bb _044_ (
    .a(_gdown_gdown_m_genblock__src_b32s_merger8_v_1334_1__m_c_2_),
    .b(_gdown_gdown_m_genblock__src_b32s_merger8_v_1334_1__m_c_3_),
    .c(_gdown_c_15_)
  );
  and_bb _045_ (
    .a(_gdown_gdown_m_genblock__src_b32s_merger8_v_1334_1__m_c_2_),
    .b(_gdown_gdown_m_genblock__src_b32s_merger8_v_1334_1__m_c_3_),
    .c(_gdown_c_14_)
  );
  or_bb _046_ (
    .a(_gdown_gdown_m_genblock__src_b32s_merger8_v_1334_1__m_c_0_),
    .b(_gdown_gdown_m_genblock__src_b32s_merger8_v_1334_1__m_c_1_),
    .c(_gdown_c_13_)
  );
  and_bb _047_ (
    .a(_gdown_gdown_m_genblock__src_b32s_merger8_v_1334_1__m_c_0_),
    .b(_gdown_gdown_m_genblock__src_b32s_merger8_v_1334_1__m_c_1_),
    .c(_gdown_c_12_)
  );
  or_bb _048_ (
    .a(a_22_),
    .b(a_23_),
    .c(_gdown_gup_gdown_c_3_)
  );
  and_bb _049_ (
    .a(a_22_),
    .b(a_23_),
    .c(_gdown_gup_gdown_c_2_)
  );
  or_bb _050_ (
    .a(a_20_),
    .b(a_21_),
    .c(_gdown_gup_gdown_c_0_)
  );
  and_bb _051_ (
    .a(a_20_),
    .b(a_21_),
    .c(_gdown_gup_gdown_c_1_)
  );
  or_bb _052_ (
    .a(_gdown_gup_gdown_c_1_),
    .b(_gdown_gup_gdown_c_3_),
    .c(_gdown_gup_gdown_g_3_c_3_)
  );
  and_bb _053_ (
    .a(_gdown_gup_gdown_c_1_),
    .b(_gdown_gup_gdown_c_3_),
    .c(_gdown_gup_gdown_g_3_c_1_)
  );
  or_bb _054_ (
    .a(_gdown_gup_gdown_c_0_),
    .b(_gdown_gup_gdown_c_2_),
    .c(_gdown_gup_gdown_g_3_c_2_)
  );
  and_bb _055_ (
    .a(_gdown_gup_gdown_c_0_),
    .b(_gdown_gup_gdown_c_2_),
    .c(_gdown_gup_gdown_g_3_c_0_)
  );
  or_bb _056_ (
    .a(_gdown_gup_gdown_g_3_c_2_),
    .b(_gdown_gup_gdown_g_3_c_3_),
    .c(_gdown_gup_c_7_)
  );
  and_bb _057_ (
    .a(_gdown_gup_gdown_g_3_c_2_),
    .b(_gdown_gup_gdown_g_3_c_3_),
    .c(_gdown_gup_c_6_)
  );
  or_bb _058_ (
    .a(_gdown_gup_gdown_g_3_c_0_),
    .b(_gdown_gup_gdown_g_3_c_1_),
    .c(_gdown_gup_c_5_)
  );
  and_bb _059_ (
    .a(_gdown_gup_gdown_g_3_c_0_),
    .b(_gdown_gup_gdown_g_3_c_1_),
    .c(_gdown_gup_c_4_)
  );
  or_bb _060_ (
    .a(a_18_),
    .b(a_19_),
    .c(_gdown_gup_gup_c_3_)
  );
  and_bb _061_ (
    .a(a_18_),
    .b(a_19_),
    .c(_gdown_gup_gup_c_2_)
  );
  or_bb _062_ (
    .a(a_16_),
    .b(a_17_),
    .c(_gdown_gup_gup_c_0_)
  );
  and_bb _063_ (
    .a(a_16_),
    .b(a_17_),
    .c(_gdown_gup_gup_c_1_)
  );
  or_bb _064_ (
    .a(_gdown_gup_gup_c_1_),
    .b(_gdown_gup_gup_c_3_),
    .c(_gdown_gup_gup_g_3_c_3_)
  );
  and_bb _065_ (
    .a(_gdown_gup_gup_c_1_),
    .b(_gdown_gup_gup_c_3_),
    .c(_gdown_gup_gup_g_3_c_1_)
  );
  or_bb _066_ (
    .a(_gdown_gup_gup_c_0_),
    .b(_gdown_gup_gup_c_2_),
    .c(_gdown_gup_gup_g_3_c_2_)
  );
  and_bb _067_ (
    .a(_gdown_gup_gup_c_0_),
    .b(_gdown_gup_gup_c_2_),
    .c(_gdown_gup_gup_g_3_c_0_)
  );
  or_bb _068_ (
    .a(_gdown_gup_gup_g_3_c_2_),
    .b(_gdown_gup_gup_g_3_c_3_),
    .c(_gdown_gup_c_0_)
  );
  and_bb _069_ (
    .a(_gdown_gup_gup_g_3_c_2_),
    .b(_gdown_gup_gup_g_3_c_3_),
    .c(_gdown_gup_c_1_)
  );
  or_bb _070_ (
    .a(_gdown_gup_gup_g_3_c_0_),
    .b(_gdown_gup_gup_g_3_c_1_),
    .c(_gdown_gup_c_2_)
  );
  and_bb _071_ (
    .a(_gdown_gup_gup_g_3_c_0_),
    .b(_gdown_gup_gup_g_3_c_1_),
    .c(_gdown_gup_c_3_)
  );
  or_bb _072_ (
    .a(_gdown_gup_c_0_),
    .b(_gdown_gup_c_4_),
    .c(_gdown_gup_m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_)
  );
  and_bb _073_ (
    .a(_gdown_gup_c_0_),
    .b(_gdown_gup_c_4_),
    .c(_gdown_gup_m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_)
  );
  or_bb _074_ (
    .a(_gdown_gup_c_1_),
    .b(_gdown_gup_c_5_),
    .c(_gdown_gup_m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_)
  );
  and_bb _075_ (
    .a(_gdown_gup_c_1_),
    .b(_gdown_gup_c_5_),
    .c(_gdown_gup_m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_)
  );
  or_bb _076_ (
    .a(_gdown_gup_c_2_),
    .b(_gdown_gup_c_6_),
    .c(_gdown_gup_m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_)
  );
  and_bb _077_ (
    .a(_gdown_gup_c_2_),
    .b(_gdown_gup_c_6_),
    .c(_gdown_gup_m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_)
  );
  or_bb _078_ (
    .a(_gdown_gup_c_3_),
    .b(_gdown_gup_c_7_),
    .c(_gdown_gup_m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_)
  );
  and_bb _079_ (
    .a(_gdown_gup_c_3_),
    .b(_gdown_gup_c_7_),
    .c(_gdown_gup_m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_)
  );
  or_bb _080_ (
    .a(_gdown_gup_m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_),
    .b(_gdown_gup_m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_),
    .c(_gdown_gup_m_genblock__src_b32s_merger8_v_1333_0__m_c_3_)
  );
  and_bb _081_ (
    .a(_gdown_gup_m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_),
    .b(_gdown_gup_m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_),
    .c(_gdown_gup_m_genblock__src_b32s_merger8_v_1333_0__m_c_1_)
  );
  or_bb _082_ (
    .a(_gdown_gup_m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_),
    .b(_gdown_gup_m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_),
    .c(_gdown_gup_m_genblock__src_b32s_merger8_v_1333_0__m_c_2_)
  );
  and_bb _083_ (
    .a(_gdown_gup_m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_),
    .b(_gdown_gup_m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_),
    .c(_gdown_gup_m_genblock__src_b32s_merger8_v_1333_0__m_c_0_)
  );
  or_bb _084_ (
    .a(_gdown_gup_m_genblock__src_b32s_merger8_v_1333_0__m_c_2_),
    .b(_gdown_gup_m_genblock__src_b32s_merger8_v_1333_0__m_c_3_),
    .c(_gdown_c_4_)
  );
  and_bb _085_ (
    .a(_gdown_gup_m_genblock__src_b32s_merger8_v_1333_0__m_c_2_),
    .b(_gdown_gup_m_genblock__src_b32s_merger8_v_1333_0__m_c_3_),
    .c(_gdown_c_5_)
  );
  or_bb _086_ (
    .a(_gdown_gup_m_genblock__src_b32s_merger8_v_1333_0__m_c_0_),
    .b(_gdown_gup_m_genblock__src_b32s_merger8_v_1333_0__m_c_1_),
    .c(_gdown_c_6_)
  );
  and_bb _087_ (
    .a(_gdown_gup_m_genblock__src_b32s_merger8_v_1333_0__m_c_0_),
    .b(_gdown_gup_m_genblock__src_b32s_merger8_v_1333_0__m_c_1_),
    .c(_gdown_c_7_)
  );
  or_bb _088_ (
    .a(_gdown_gup_m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_),
    .b(_gdown_gup_m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_),
    .c(_gdown_gup_m_genblock__src_b32s_merger8_v_1334_1__m_c_3_)
  );
  and_bb _089_ (
    .a(_gdown_gup_m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_),
    .b(_gdown_gup_m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_),
    .c(_gdown_gup_m_genblock__src_b32s_merger8_v_1334_1__m_c_1_)
  );
  or_bb _090_ (
    .a(_gdown_gup_m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_),
    .b(_gdown_gup_m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_),
    .c(_gdown_gup_m_genblock__src_b32s_merger8_v_1334_1__m_c_2_)
  );
  and_bb _091_ (
    .a(_gdown_gup_m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_),
    .b(_gdown_gup_m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_),
    .c(_gdown_gup_m_genblock__src_b32s_merger8_v_1334_1__m_c_0_)
  );
  or_bb _092_ (
    .a(_gdown_gup_m_genblock__src_b32s_merger8_v_1334_1__m_c_2_),
    .b(_gdown_gup_m_genblock__src_b32s_merger8_v_1334_1__m_c_3_),
    .c(_gdown_c_0_)
  );
  and_bb _093_ (
    .a(_gdown_gup_m_genblock__src_b32s_merger8_v_1334_1__m_c_2_),
    .b(_gdown_gup_m_genblock__src_b32s_merger8_v_1334_1__m_c_3_),
    .c(_gdown_c_1_)
  );
  or_bb _094_ (
    .a(_gdown_gup_m_genblock__src_b32s_merger8_v_1334_1__m_c_0_),
    .b(_gdown_gup_m_genblock__src_b32s_merger8_v_1334_1__m_c_1_),
    .c(_gdown_c_2_)
  );
  and_bb _095_ (
    .a(_gdown_gup_m_genblock__src_b32s_merger8_v_1334_1__m_c_0_),
    .b(_gdown_gup_m_genblock__src_b32s_merger8_v_1334_1__m_c_1_),
    .c(_gdown_c_3_)
  );
  or_bb _096_ (
    .a(_gdown_c_0_),
    .b(_gdown_c_8_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_101_0__g_ord_1_)
  );
  and_bb _097_ (
    .a(_gdown_c_0_),
    .b(_gdown_c_8_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_101_0__g_ord_0_)
  );
  or_bb _098_ (
    .a(_gdown_c_1_),
    .b(_gdown_c_9_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_102_1__g_ord_1_)
  );
  and_bb _099_ (
    .a(_gdown_c_1_),
    .b(_gdown_c_9_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_102_1__g_ord_0_)
  );
  or_bb _100_ (
    .a(_gdown_c_2_),
    .b(_gdown_c_10_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_103_2__g_ord_1_)
  );
  and_bb _101_ (
    .a(_gdown_c_2_),
    .b(_gdown_c_10_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_103_2__g_ord_0_)
  );
  or_bb _102_ (
    .a(_gdown_c_3_),
    .b(_gdown_c_11_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_104_3__g_ord_1_)
  );
  and_bb _103_ (
    .a(_gdown_c_3_),
    .b(_gdown_c_11_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_104_3__g_ord_0_)
  );
  or_bb _104_ (
    .a(_gdown_c_4_),
    .b(_gdown_c_12_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_105_4__g_ord_1_)
  );
  and_bb _105_ (
    .a(_gdown_c_4_),
    .b(_gdown_c_12_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_105_4__g_ord_0_)
  );
  or_bb _106_ (
    .a(_gdown_c_5_),
    .b(_gdown_c_13_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_106_5__g_ord_1_)
  );
  and_bb _107_ (
    .a(_gdown_c_5_),
    .b(_gdown_c_13_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_106_5__g_ord_0_)
  );
  or_bb _108_ (
    .a(_gdown_c_6_),
    .b(_gdown_c_14_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_107_6__g_ord_1_)
  );
  and_bb _109_ (
    .a(_gdown_c_6_),
    .b(_gdown_c_14_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_107_6__g_ord_0_)
  );
  or_bb _110_ (
    .a(_gdown_c_7_),
    .b(_gdown_c_15_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_108_7__g_ord_1_)
  );
  and_bb _111_ (
    .a(_gdown_c_7_),
    .b(_gdown_c_15_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_108_7__g_ord_0_)
  );
  or_bb _112_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_101_0__g_ord_1_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_105_4__g_ord_1_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_)
  );
  and_bb _113_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_101_0__g_ord_1_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_105_4__g_ord_1_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_)
  );
  or_bb _114_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_102_1__g_ord_1_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_106_5__g_ord_1_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_)
  );
  and_bb _115_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_102_1__g_ord_1_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_106_5__g_ord_1_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_)
  );
  or_bb _116_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_103_2__g_ord_1_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_107_6__g_ord_1_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_)
  );
  and_bb _117_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_103_2__g_ord_1_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_107_6__g_ord_1_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_)
  );
  or_bb _118_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_104_3__g_ord_1_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_108_7__g_ord_1_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_)
  );
  and_bb _119_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_104_3__g_ord_1_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_108_7__g_ord_1_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_)
  );
  or_bb _120_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_3_)
  );
  and_bb _121_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_1_)
  );
  or_bb _122_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_2_)
  );
  and_bb _123_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_0_)
  );
  or_bb _124_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_2_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_3_),
    .c(c_27_)
  );
  and_bb _125_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_2_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_3_),
    .c(c_26_)
  );
  or_bb _126_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_0_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_1_),
    .c(c_25_)
  );
  and_bb _127_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_0_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_1_),
    .c(c_24_)
  );
  or_bb _128_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_3_)
  );
  and_bb _129_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_1_)
  );
  or_bb _130_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_2_)
  );
  and_bb _131_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_0_)
  );
  or_bb _132_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_2_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_3_),
    .c(c_31_)
  );
  and_bb _133_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_2_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_3_),
    .c(c_30_)
  );
  or_bb _134_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_0_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_1_),
    .c(c_29_)
  );
  and_bb _135_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_0_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_1_),
    .c(c_28_)
  );
  or_bb _136_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_101_0__g_ord_0_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_105_4__g_ord_0_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_)
  );
  and_bb _137_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_101_0__g_ord_0_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_105_4__g_ord_0_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_)
  );
  or_bb _138_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_102_1__g_ord_0_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_106_5__g_ord_0_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_)
  );
  and_bb _139_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_102_1__g_ord_0_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_106_5__g_ord_0_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_)
  );
  or_bb _140_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_103_2__g_ord_0_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_107_6__g_ord_0_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_)
  );
  and_bb _141_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_103_2__g_ord_0_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_107_6__g_ord_0_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_)
  );
  or_bb _142_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_104_3__g_ord_0_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_108_7__g_ord_0_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_)
  );
  and_bb _143_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_104_3__g_ord_0_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_108_7__g_ord_0_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_)
  );
  or_bb _144_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_3_)
  );
  and_bb _145_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_1_)
  );
  or_bb _146_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_2_)
  );
  and_bb _147_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_0_)
  );
  or_bb _148_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_2_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_3_),
    .c(c_19_)
  );
  and_bb _149_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_2_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_3_),
    .c(c_18_)
  );
  or_bb _150_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_0_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_1_),
    .c(c_17_)
  );
  and_bb _151_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_0_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_1_),
    .c(c_16_)
  );
  or_bb _152_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_3_)
  );
  and_bb _153_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_1_)
  );
  or_bb _154_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_2_)
  );
  and_bb _155_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_),
    .c(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_0_)
  );
  or_bb _156_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_2_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_3_),
    .c(c_23_)
  );
  and_bb _157_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_2_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_3_),
    .c(c_22_)
  );
  or_bb _158_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_0_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_1_),
    .c(c_21_)
  );
  and_bb _159_ (
    .a(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_0_),
    .b(_gdown_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_1_),
    .c(c_20_)
  );
  or_bb _160_ (
    .a(a_14_),
    .b(a_15_),
    .c(_gup_gdown_gdown_c_3_)
  );
  and_bb _161_ (
    .a(a_14_),
    .b(a_15_),
    .c(_gup_gdown_gdown_c_2_)
  );
  or_bb _162_ (
    .a(a_12_),
    .b(a_13_),
    .c(_gup_gdown_gdown_c_0_)
  );
  and_bb _163_ (
    .a(a_12_),
    .b(a_13_),
    .c(_gup_gdown_gdown_c_1_)
  );
  or_bb _164_ (
    .a(_gup_gdown_gdown_c_1_),
    .b(_gup_gdown_gdown_c_3_),
    .c(_gup_gdown_gdown_g_3_c_3_)
  );
  and_bb _165_ (
    .a(_gup_gdown_gdown_c_1_),
    .b(_gup_gdown_gdown_c_3_),
    .c(_gup_gdown_gdown_g_3_c_1_)
  );
  or_bb _166_ (
    .a(_gup_gdown_gdown_c_0_),
    .b(_gup_gdown_gdown_c_2_),
    .c(_gup_gdown_gdown_g_3_c_2_)
  );
  and_bb _167_ (
    .a(_gup_gdown_gdown_c_0_),
    .b(_gup_gdown_gdown_c_2_),
    .c(_gup_gdown_gdown_g_3_c_0_)
  );
  or_bb _168_ (
    .a(_gup_gdown_gdown_g_3_c_2_),
    .b(_gup_gdown_gdown_g_3_c_3_),
    .c(_gup_gdown_c_7_)
  );
  and_bb _169_ (
    .a(_gup_gdown_gdown_g_3_c_2_),
    .b(_gup_gdown_gdown_g_3_c_3_),
    .c(_gup_gdown_c_6_)
  );
  or_bb _170_ (
    .a(_gup_gdown_gdown_g_3_c_0_),
    .b(_gup_gdown_gdown_g_3_c_1_),
    .c(_gup_gdown_c_5_)
  );
  and_bb _171_ (
    .a(_gup_gdown_gdown_g_3_c_0_),
    .b(_gup_gdown_gdown_g_3_c_1_),
    .c(_gup_gdown_c_4_)
  );
  or_bb _172_ (
    .a(a_10_),
    .b(a_11_),
    .c(_gup_gdown_gup_c_3_)
  );
  and_bb _173_ (
    .a(a_10_),
    .b(a_11_),
    .c(_gup_gdown_gup_c_2_)
  );
  or_bb _174_ (
    .a(a_8_),
    .b(a_9_),
    .c(_gup_gdown_gup_c_0_)
  );
  and_bb _175_ (
    .a(a_8_),
    .b(a_9_),
    .c(_gup_gdown_gup_c_1_)
  );
  or_bb _176_ (
    .a(_gup_gdown_gup_c_1_),
    .b(_gup_gdown_gup_c_3_),
    .c(_gup_gdown_gup_g_3_c_3_)
  );
  and_bb _177_ (
    .a(_gup_gdown_gup_c_1_),
    .b(_gup_gdown_gup_c_3_),
    .c(_gup_gdown_gup_g_3_c_1_)
  );
  or_bb _178_ (
    .a(_gup_gdown_gup_c_0_),
    .b(_gup_gdown_gup_c_2_),
    .c(_gup_gdown_gup_g_3_c_2_)
  );
  and_bb _179_ (
    .a(_gup_gdown_gup_c_0_),
    .b(_gup_gdown_gup_c_2_),
    .c(_gup_gdown_gup_g_3_c_0_)
  );
  or_bb _180_ (
    .a(_gup_gdown_gup_g_3_c_2_),
    .b(_gup_gdown_gup_g_3_c_3_),
    .c(_gup_gdown_c_0_)
  );
  and_bb _181_ (
    .a(_gup_gdown_gup_g_3_c_2_),
    .b(_gup_gdown_gup_g_3_c_3_),
    .c(_gup_gdown_c_1_)
  );
  or_bb _182_ (
    .a(_gup_gdown_gup_g_3_c_0_),
    .b(_gup_gdown_gup_g_3_c_1_),
    .c(_gup_gdown_c_2_)
  );
  and_bb _183_ (
    .a(_gup_gdown_gup_g_3_c_0_),
    .b(_gup_gdown_gup_g_3_c_1_),
    .c(_gup_gdown_c_3_)
  );
  or_bb _184_ (
    .a(_gup_gdown_c_0_),
    .b(_gup_gdown_c_4_),
    .c(_gup_gdown_m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_)
  );
  and_bb _185_ (
    .a(_gup_gdown_c_0_),
    .b(_gup_gdown_c_4_),
    .c(_gup_gdown_m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_)
  );
  or_bb _186_ (
    .a(_gup_gdown_c_1_),
    .b(_gup_gdown_c_5_),
    .c(_gup_gdown_m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_)
  );
  and_bb _187_ (
    .a(_gup_gdown_c_1_),
    .b(_gup_gdown_c_5_),
    .c(_gup_gdown_m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_)
  );
  or_bb _188_ (
    .a(_gup_gdown_c_2_),
    .b(_gup_gdown_c_6_),
    .c(_gup_gdown_m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_)
  );
  and_bb _189_ (
    .a(_gup_gdown_c_2_),
    .b(_gup_gdown_c_6_),
    .c(_gup_gdown_m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_)
  );
  or_bb _190_ (
    .a(_gup_gdown_c_3_),
    .b(_gup_gdown_c_7_),
    .c(_gup_gdown_m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_)
  );
  and_bb _191_ (
    .a(_gup_gdown_c_3_),
    .b(_gup_gdown_c_7_),
    .c(_gup_gdown_m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_)
  );
  or_bb _192_ (
    .a(_gup_gdown_m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_),
    .b(_gup_gdown_m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_),
    .c(_gup_gdown_m_genblock__src_b32s_merger8_v_1333_0__m_c_3_)
  );
  and_bb _193_ (
    .a(_gup_gdown_m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_),
    .b(_gup_gdown_m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_),
    .c(_gup_gdown_m_genblock__src_b32s_merger8_v_1333_0__m_c_1_)
  );
  or_bb _194_ (
    .a(_gup_gdown_m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_),
    .b(_gup_gdown_m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_),
    .c(_gup_gdown_m_genblock__src_b32s_merger8_v_1333_0__m_c_2_)
  );
  and_bb _195_ (
    .a(_gup_gdown_m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_),
    .b(_gup_gdown_m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_),
    .c(_gup_gdown_m_genblock__src_b32s_merger8_v_1333_0__m_c_0_)
  );
  or_bb _196_ (
    .a(_gup_gdown_m_genblock__src_b32s_merger8_v_1333_0__m_c_2_),
    .b(_gup_gdown_m_genblock__src_b32s_merger8_v_1333_0__m_c_3_),
    .c(_gup_c_11_)
  );
  and_bb _197_ (
    .a(_gup_gdown_m_genblock__src_b32s_merger8_v_1333_0__m_c_2_),
    .b(_gup_gdown_m_genblock__src_b32s_merger8_v_1333_0__m_c_3_),
    .c(_gup_c_10_)
  );
  or_bb _198_ (
    .a(_gup_gdown_m_genblock__src_b32s_merger8_v_1333_0__m_c_0_),
    .b(_gup_gdown_m_genblock__src_b32s_merger8_v_1333_0__m_c_1_),
    .c(_gup_c_9_)
  );
  and_bb _199_ (
    .a(_gup_gdown_m_genblock__src_b32s_merger8_v_1333_0__m_c_0_),
    .b(_gup_gdown_m_genblock__src_b32s_merger8_v_1333_0__m_c_1_),
    .c(_gup_c_8_)
  );
  or_bb _200_ (
    .a(_gup_gdown_m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_),
    .b(_gup_gdown_m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_),
    .c(_gup_gdown_m_genblock__src_b32s_merger8_v_1334_1__m_c_3_)
  );
  and_bb _201_ (
    .a(_gup_gdown_m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_),
    .b(_gup_gdown_m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_),
    .c(_gup_gdown_m_genblock__src_b32s_merger8_v_1334_1__m_c_1_)
  );
  or_bb _202_ (
    .a(_gup_gdown_m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_),
    .b(_gup_gdown_m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_),
    .c(_gup_gdown_m_genblock__src_b32s_merger8_v_1334_1__m_c_2_)
  );
  and_bb _203_ (
    .a(_gup_gdown_m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_),
    .b(_gup_gdown_m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_),
    .c(_gup_gdown_m_genblock__src_b32s_merger8_v_1334_1__m_c_0_)
  );
  or_bb _204_ (
    .a(_gup_gdown_m_genblock__src_b32s_merger8_v_1334_1__m_c_2_),
    .b(_gup_gdown_m_genblock__src_b32s_merger8_v_1334_1__m_c_3_),
    .c(_gup_c_15_)
  );
  and_bb _205_ (
    .a(_gup_gdown_m_genblock__src_b32s_merger8_v_1334_1__m_c_2_),
    .b(_gup_gdown_m_genblock__src_b32s_merger8_v_1334_1__m_c_3_),
    .c(_gup_c_14_)
  );
  or_bb _206_ (
    .a(_gup_gdown_m_genblock__src_b32s_merger8_v_1334_1__m_c_0_),
    .b(_gup_gdown_m_genblock__src_b32s_merger8_v_1334_1__m_c_1_),
    .c(_gup_c_13_)
  );
  and_bb _207_ (
    .a(_gup_gdown_m_genblock__src_b32s_merger8_v_1334_1__m_c_0_),
    .b(_gup_gdown_m_genblock__src_b32s_merger8_v_1334_1__m_c_1_),
    .c(_gup_c_12_)
  );
  or_bb _208_ (
    .a(a_6_),
    .b(a_7_),
    .c(_gup_gup_gdown_c_3_)
  );
  and_bb _209_ (
    .a(a_6_),
    .b(a_7_),
    .c(_gup_gup_gdown_c_2_)
  );
  or_bb _210_ (
    .a(a_4_),
    .b(a_5_),
    .c(_gup_gup_gdown_c_0_)
  );
  and_bb _211_ (
    .a(a_4_),
    .b(a_5_),
    .c(_gup_gup_gdown_c_1_)
  );
  or_bb _212_ (
    .a(_gup_gup_gdown_c_1_),
    .b(_gup_gup_gdown_c_3_),
    .c(_gup_gup_gdown_g_3_c_3_)
  );
  and_bb _213_ (
    .a(_gup_gup_gdown_c_1_),
    .b(_gup_gup_gdown_c_3_),
    .c(_gup_gup_gdown_g_3_c_1_)
  );
  or_bb _214_ (
    .a(_gup_gup_gdown_c_0_),
    .b(_gup_gup_gdown_c_2_),
    .c(_gup_gup_gdown_g_3_c_2_)
  );
  and_bb _215_ (
    .a(_gup_gup_gdown_c_0_),
    .b(_gup_gup_gdown_c_2_),
    .c(_gup_gup_gdown_g_3_c_0_)
  );
  or_bb _216_ (
    .a(_gup_gup_gdown_g_3_c_2_),
    .b(_gup_gup_gdown_g_3_c_3_),
    .c(_gup_gup_c_7_)
  );
  and_bb _217_ (
    .a(_gup_gup_gdown_g_3_c_2_),
    .b(_gup_gup_gdown_g_3_c_3_),
    .c(_gup_gup_c_6_)
  );
  or_bb _218_ (
    .a(_gup_gup_gdown_g_3_c_0_),
    .b(_gup_gup_gdown_g_3_c_1_),
    .c(_gup_gup_c_5_)
  );
  and_bb _219_ (
    .a(_gup_gup_gdown_g_3_c_0_),
    .b(_gup_gup_gdown_g_3_c_1_),
    .c(_gup_gup_c_4_)
  );
  or_bb _220_ (
    .a(a_2_),
    .b(a_3_),
    .c(_gup_gup_gup_c_3_)
  );
  and_bb _221_ (
    .a(a_2_),
    .b(a_3_),
    .c(_gup_gup_gup_c_2_)
  );
  or_bb _222_ (
    .a(a_0_),
    .b(a_1_),
    .c(_gup_gup_gup_c_0_)
  );
  and_bb _223_ (
    .a(a_0_),
    .b(a_1_),
    .c(_gup_gup_gup_c_1_)
  );
  or_bb _224_ (
    .a(_gup_gup_gup_c_1_),
    .b(_gup_gup_gup_c_3_),
    .c(_gup_gup_gup_g_3_c_3_)
  );
  and_bb _225_ (
    .a(_gup_gup_gup_c_1_),
    .b(_gup_gup_gup_c_3_),
    .c(_gup_gup_gup_g_3_c_1_)
  );
  or_bb _226_ (
    .a(_gup_gup_gup_c_0_),
    .b(_gup_gup_gup_c_2_),
    .c(_gup_gup_gup_g_3_c_2_)
  );
  and_bb _227_ (
    .a(_gup_gup_gup_c_0_),
    .b(_gup_gup_gup_c_2_),
    .c(_gup_gup_gup_g_3_c_0_)
  );
  or_bb _228_ (
    .a(_gup_gup_gup_g_3_c_2_),
    .b(_gup_gup_gup_g_3_c_3_),
    .c(_gup_gup_c_0_)
  );
  and_bb _229_ (
    .a(_gup_gup_gup_g_3_c_2_),
    .b(_gup_gup_gup_g_3_c_3_),
    .c(_gup_gup_c_1_)
  );
  or_bb _230_ (
    .a(_gup_gup_gup_g_3_c_0_),
    .b(_gup_gup_gup_g_3_c_1_),
    .c(_gup_gup_c_2_)
  );
  and_bb _231_ (
    .a(_gup_gup_gup_g_3_c_0_),
    .b(_gup_gup_gup_g_3_c_1_),
    .c(_gup_gup_c_3_)
  );
  or_bb _232_ (
    .a(_gup_gup_c_0_),
    .b(_gup_gup_c_4_),
    .c(_gup_gup_m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_)
  );
  and_bb _233_ (
    .a(_gup_gup_c_0_),
    .b(_gup_gup_c_4_),
    .c(_gup_gup_m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_)
  );
  or_bb _234_ (
    .a(_gup_gup_c_1_),
    .b(_gup_gup_c_5_),
    .c(_gup_gup_m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_)
  );
  and_bb _235_ (
    .a(_gup_gup_c_1_),
    .b(_gup_gup_c_5_),
    .c(_gup_gup_m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_)
  );
  or_bb _236_ (
    .a(_gup_gup_c_2_),
    .b(_gup_gup_c_6_),
    .c(_gup_gup_m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_)
  );
  and_bb _237_ (
    .a(_gup_gup_c_2_),
    .b(_gup_gup_c_6_),
    .c(_gup_gup_m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_)
  );
  or_bb _238_ (
    .a(_gup_gup_c_3_),
    .b(_gup_gup_c_7_),
    .c(_gup_gup_m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_)
  );
  and_bb _239_ (
    .a(_gup_gup_c_3_),
    .b(_gup_gup_c_7_),
    .c(_gup_gup_m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_)
  );
  or_bb _240_ (
    .a(_gup_gup_m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_),
    .b(_gup_gup_m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_),
    .c(_gup_gup_m_genblock__src_b32s_merger8_v_1333_0__m_c_3_)
  );
  and_bb _241_ (
    .a(_gup_gup_m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_),
    .b(_gup_gup_m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_),
    .c(_gup_gup_m_genblock__src_b32s_merger8_v_1333_0__m_c_1_)
  );
  or_bb _242_ (
    .a(_gup_gup_m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_),
    .b(_gup_gup_m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_),
    .c(_gup_gup_m_genblock__src_b32s_merger8_v_1333_0__m_c_2_)
  );
  and_bb _243_ (
    .a(_gup_gup_m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_),
    .b(_gup_gup_m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_),
    .c(_gup_gup_m_genblock__src_b32s_merger8_v_1333_0__m_c_0_)
  );
  or_bb _244_ (
    .a(_gup_gup_m_genblock__src_b32s_merger8_v_1333_0__m_c_2_),
    .b(_gup_gup_m_genblock__src_b32s_merger8_v_1333_0__m_c_3_),
    .c(_gup_c_4_)
  );
  and_bb _245_ (
    .a(_gup_gup_m_genblock__src_b32s_merger8_v_1333_0__m_c_2_),
    .b(_gup_gup_m_genblock__src_b32s_merger8_v_1333_0__m_c_3_),
    .c(_gup_c_5_)
  );
  or_bb _246_ (
    .a(_gup_gup_m_genblock__src_b32s_merger8_v_1333_0__m_c_0_),
    .b(_gup_gup_m_genblock__src_b32s_merger8_v_1333_0__m_c_1_),
    .c(_gup_c_6_)
  );
  and_bb _247_ (
    .a(_gup_gup_m_genblock__src_b32s_merger8_v_1333_0__m_c_0_),
    .b(_gup_gup_m_genblock__src_b32s_merger8_v_1333_0__m_c_1_),
    .c(_gup_c_7_)
  );
  or_bb _248_ (
    .a(_gup_gup_m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_),
    .b(_gup_gup_m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_),
    .c(_gup_gup_m_genblock__src_b32s_merger8_v_1334_1__m_c_3_)
  );
  and_bb _249_ (
    .a(_gup_gup_m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_),
    .b(_gup_gup_m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_),
    .c(_gup_gup_m_genblock__src_b32s_merger8_v_1334_1__m_c_1_)
  );
  or_bb _250_ (
    .a(_gup_gup_m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_),
    .b(_gup_gup_m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_),
    .c(_gup_gup_m_genblock__src_b32s_merger8_v_1334_1__m_c_2_)
  );
  and_bb _251_ (
    .a(_gup_gup_m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_),
    .b(_gup_gup_m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_),
    .c(_gup_gup_m_genblock__src_b32s_merger8_v_1334_1__m_c_0_)
  );
  or_bb _252_ (
    .a(_gup_gup_m_genblock__src_b32s_merger8_v_1334_1__m_c_2_),
    .b(_gup_gup_m_genblock__src_b32s_merger8_v_1334_1__m_c_3_),
    .c(_gup_c_0_)
  );
  and_bb _253_ (
    .a(_gup_gup_m_genblock__src_b32s_merger8_v_1334_1__m_c_2_),
    .b(_gup_gup_m_genblock__src_b32s_merger8_v_1334_1__m_c_3_),
    .c(_gup_c_1_)
  );
  or_bb _254_ (
    .a(_gup_gup_m_genblock__src_b32s_merger8_v_1334_1__m_c_0_),
    .b(_gup_gup_m_genblock__src_b32s_merger8_v_1334_1__m_c_1_),
    .c(_gup_c_2_)
  );
  and_bb _255_ (
    .a(_gup_gup_m_genblock__src_b32s_merger8_v_1334_1__m_c_0_),
    .b(_gup_gup_m_genblock__src_b32s_merger8_v_1334_1__m_c_1_),
    .c(_gup_c_3_)
  );
  or_bb _256_ (
    .a(_gup_c_0_),
    .b(_gup_c_8_),
    .c(_gup_m_genblock__src_b32s_merger16_v_101_0__g_ord_1_)
  );
  and_bb _257_ (
    .a(_gup_c_0_),
    .b(_gup_c_8_),
    .c(_gup_m_genblock__src_b32s_merger16_v_101_0__g_ord_0_)
  );
  or_bb _258_ (
    .a(_gup_c_1_),
    .b(_gup_c_9_),
    .c(_gup_m_genblock__src_b32s_merger16_v_102_1__g_ord_1_)
  );
  and_bb _259_ (
    .a(_gup_c_1_),
    .b(_gup_c_9_),
    .c(_gup_m_genblock__src_b32s_merger16_v_102_1__g_ord_0_)
  );
  or_bb _260_ (
    .a(_gup_c_2_),
    .b(_gup_c_10_),
    .c(_gup_m_genblock__src_b32s_merger16_v_103_2__g_ord_1_)
  );
  and_bb _261_ (
    .a(_gup_c_2_),
    .b(_gup_c_10_),
    .c(_gup_m_genblock__src_b32s_merger16_v_103_2__g_ord_0_)
  );
  or_bb _262_ (
    .a(_gup_c_3_),
    .b(_gup_c_11_),
    .c(_gup_m_genblock__src_b32s_merger16_v_104_3__g_ord_1_)
  );
  and_bb _263_ (
    .a(_gup_c_3_),
    .b(_gup_c_11_),
    .c(_gup_m_genblock__src_b32s_merger16_v_104_3__g_ord_0_)
  );
  or_bb _264_ (
    .a(_gup_c_4_),
    .b(_gup_c_12_),
    .c(_gup_m_genblock__src_b32s_merger16_v_105_4__g_ord_1_)
  );
  and_bb _265_ (
    .a(_gup_c_4_),
    .b(_gup_c_12_),
    .c(_gup_m_genblock__src_b32s_merger16_v_105_4__g_ord_0_)
  );
  or_bb _266_ (
    .a(_gup_c_5_),
    .b(_gup_c_13_),
    .c(_gup_m_genblock__src_b32s_merger16_v_106_5__g_ord_1_)
  );
  and_bb _267_ (
    .a(_gup_c_5_),
    .b(_gup_c_13_),
    .c(_gup_m_genblock__src_b32s_merger16_v_106_5__g_ord_0_)
  );
  or_bb _268_ (
    .a(_gup_c_6_),
    .b(_gup_c_14_),
    .c(_gup_m_genblock__src_b32s_merger16_v_107_6__g_ord_1_)
  );
  and_bb _269_ (
    .a(_gup_c_6_),
    .b(_gup_c_14_),
    .c(_gup_m_genblock__src_b32s_merger16_v_107_6__g_ord_0_)
  );
  or_bb _270_ (
    .a(_gup_c_7_),
    .b(_gup_c_15_),
    .c(_gup_m_genblock__src_b32s_merger16_v_108_7__g_ord_1_)
  );
  and_bb _271_ (
    .a(_gup_c_7_),
    .b(_gup_c_15_),
    .c(_gup_m_genblock__src_b32s_merger16_v_108_7__g_ord_0_)
  );
  or_bb _272_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_101_0__g_ord_1_),
    .b(_gup_m_genblock__src_b32s_merger16_v_105_4__g_ord_1_),
    .c(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_)
  );
  and_bb _273_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_101_0__g_ord_1_),
    .b(_gup_m_genblock__src_b32s_merger16_v_105_4__g_ord_1_),
    .c(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_)
  );
  or_bb _274_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_102_1__g_ord_1_),
    .b(_gup_m_genblock__src_b32s_merger16_v_106_5__g_ord_1_),
    .c(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_)
  );
  and_bb _275_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_102_1__g_ord_1_),
    .b(_gup_m_genblock__src_b32s_merger16_v_106_5__g_ord_1_),
    .c(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_)
  );
  or_bb _276_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_103_2__g_ord_1_),
    .b(_gup_m_genblock__src_b32s_merger16_v_107_6__g_ord_1_),
    .c(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_)
  );
  and_bb _277_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_103_2__g_ord_1_),
    .b(_gup_m_genblock__src_b32s_merger16_v_107_6__g_ord_1_),
    .c(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_)
  );
  or_bb _278_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_104_3__g_ord_1_),
    .b(_gup_m_genblock__src_b32s_merger16_v_108_7__g_ord_1_),
    .c(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_)
  );
  and_bb _279_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_104_3__g_ord_1_),
    .b(_gup_m_genblock__src_b32s_merger16_v_108_7__g_ord_1_),
    .c(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_)
  );
  or_bb _280_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_),
    .b(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_),
    .c(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_3_)
  );
  and_bb _281_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_),
    .b(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_),
    .c(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_1_)
  );
  or_bb _282_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_),
    .b(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_),
    .c(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_2_)
  );
  and_bb _283_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_),
    .b(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_),
    .c(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_0_)
  );
  or_bb _284_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_2_),
    .b(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_3_),
    .c(c_4_)
  );
  and_bb _285_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_2_),
    .b(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_3_),
    .c(c_5_)
  );
  or_bb _286_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_0_),
    .b(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_1_),
    .c(c_6_)
  );
  and_bb _287_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_0_),
    .b(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_1_),
    .c(c_7_)
  );
  or_bb _288_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_),
    .b(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_),
    .c(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_3_)
  );
  and_bb _289_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_),
    .b(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_),
    .c(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_1_)
  );
  or_bb _290_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_),
    .b(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_),
    .c(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_2_)
  );
  and_bb _291_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_),
    .b(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_),
    .c(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_0_)
  );
  or_bb _292_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_2_),
    .b(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_3_),
    .c(c_0_)
  );
  and_bb _293_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_2_),
    .b(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_3_),
    .c(c_1_)
  );
  or_bb _294_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_0_),
    .b(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_1_),
    .c(c_2_)
  );
  and_bb _295_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_0_),
    .b(_gup_m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_1_),
    .c(c_3_)
  );
  or_bb _296_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_101_0__g_ord_0_),
    .b(_gup_m_genblock__src_b32s_merger16_v_105_4__g_ord_0_),
    .c(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_)
  );
  and_bb _297_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_101_0__g_ord_0_),
    .b(_gup_m_genblock__src_b32s_merger16_v_105_4__g_ord_0_),
    .c(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_)
  );
  or_bb _298_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_102_1__g_ord_0_),
    .b(_gup_m_genblock__src_b32s_merger16_v_106_5__g_ord_0_),
    .c(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_)
  );
  and_bb _299_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_102_1__g_ord_0_),
    .b(_gup_m_genblock__src_b32s_merger16_v_106_5__g_ord_0_),
    .c(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_)
  );
  or_bb _300_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_103_2__g_ord_0_),
    .b(_gup_m_genblock__src_b32s_merger16_v_107_6__g_ord_0_),
    .c(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_)
  );
  and_bb _301_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_103_2__g_ord_0_),
    .b(_gup_m_genblock__src_b32s_merger16_v_107_6__g_ord_0_),
    .c(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_)
  );
  or_bb _302_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_104_3__g_ord_0_),
    .b(_gup_m_genblock__src_b32s_merger16_v_108_7__g_ord_0_),
    .c(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_)
  );
  and_bb _303_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_104_3__g_ord_0_),
    .b(_gup_m_genblock__src_b32s_merger16_v_108_7__g_ord_0_),
    .c(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_)
  );
  or_bb _304_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_),
    .b(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_),
    .c(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_3_)
  );
  and_bb _305_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_),
    .b(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_),
    .c(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_1_)
  );
  or_bb _306_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_),
    .b(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_),
    .c(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_2_)
  );
  and_bb _307_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_),
    .b(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_),
    .c(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_0_)
  );
  or_bb _308_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_2_),
    .b(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_3_),
    .c(c_12_)
  );
  and_bb _309_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_2_),
    .b(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_3_),
    .c(c_13_)
  );
  or_bb _310_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_0_),
    .b(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_1_),
    .c(c_14_)
  );
  and_bb _311_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_0_),
    .b(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_1_),
    .c(c_15_)
  );
  or_bb _312_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_),
    .b(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_),
    .c(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_3_)
  );
  and_bb _313_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_),
    .b(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_),
    .c(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_1_)
  );
  or_bb _314_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_),
    .b(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_),
    .c(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_2_)
  );
  and_bb _315_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_),
    .b(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_),
    .c(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_0_)
  );
  or_bb _316_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_2_),
    .b(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_3_),
    .c(c_8_)
  );
  and_bb _317_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_2_),
    .b(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_3_),
    .c(c_9_)
  );
  or_bb _318_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_0_),
    .b(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_1_),
    .c(c_10_)
  );
  and_bb _319_ (
    .a(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_0_),
    .b(_gup_m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_1_),
    .c(c_11_)
  );
  or_bb _320_ (
    .a(c_0_),
    .b(c_16_),
    .c(_m_genblock__src_b32s_merger32_v_1011_0__g_ord_1_)
  );
  and_bb _321_ (
    .a(c_0_),
    .b(c_16_),
    .c(_m_genblock__src_b32s_merger32_v_1011_0__g_ord_0_)
  );
  or_bb _322_ (
    .a(c_1_),
    .b(c_17_),
    .c(_m_genblock__src_b32s_merger32_v_1012_1__g_ord_1_)
  );
  and_bb _323_ (
    .a(c_1_),
    .b(c_17_),
    .c(_m_genblock__src_b32s_merger32_v_1012_1__g_ord_0_)
  );
  or_bb _324_ (
    .a(c_2_),
    .b(c_18_),
    .c(_m_genblock__src_b32s_merger32_v_1013_2__g_ord_1_)
  );
  and_bb _325_ (
    .a(c_2_),
    .b(c_18_),
    .c(_m_genblock__src_b32s_merger32_v_1013_2__g_ord_0_)
  );
  or_bb _326_ (
    .a(c_3_),
    .b(c_19_),
    .c(_m_genblock__src_b32s_merger32_v_1014_3__g_ord_1_)
  );
  and_bb _327_ (
    .a(c_3_),
    .b(c_19_),
    .c(_m_genblock__src_b32s_merger32_v_1014_3__g_ord_0_)
  );
  or_bb _328_ (
    .a(c_4_),
    .b(c_20_),
    .c(_m_genblock__src_b32s_merger32_v_1015_4__g_ord_1_)
  );
  and_bb _329_ (
    .a(c_4_),
    .b(c_20_),
    .c(_m_genblock__src_b32s_merger32_v_1015_4__g_ord_0_)
  );
  or_bb _330_ (
    .a(c_5_),
    .b(c_21_),
    .c(_m_genblock__src_b32s_merger32_v_1016_5__g_ord_1_)
  );
  and_bb _331_ (
    .a(c_5_),
    .b(c_21_),
    .c(_m_genblock__src_b32s_merger32_v_1016_5__g_ord_0_)
  );
  or_bb _332_ (
    .a(c_6_),
    .b(c_22_),
    .c(_m_genblock__src_b32s_merger32_v_1017_6__g_ord_1_)
  );
  and_bb _333_ (
    .a(c_6_),
    .b(c_22_),
    .c(_m_genblock__src_b32s_merger32_v_1017_6__g_ord_0_)
  );
  or_bb _334_ (
    .a(c_7_),
    .b(c_23_),
    .c(_m_genblock__src_b32s_merger32_v_1018_7__g_ord_1_)
  );
  and_bb _335_ (
    .a(c_7_),
    .b(c_23_),
    .c(_m_genblock__src_b32s_merger32_v_1018_7__g_ord_0_)
  );
  or_bb _336_ (
    .a(c_8_),
    .b(c_24_),
    .c(_m_genblock__src_b32s_merger32_v_1019_8__g_ord_1_)
  );
  and_bb _337_ (
    .a(c_8_),
    .b(c_24_),
    .c(_m_genblock__src_b32s_merger32_v_1019_8__g_ord_0_)
  );
  or_bb _338_ (
    .a(c_9_),
    .b(c_25_),
    .c(_m_genblock__src_b32s_merger32_v_1020_9__g_ord_1_)
  );
  and_bb _339_ (
    .a(c_9_),
    .b(c_25_),
    .c(_m_genblock__src_b32s_merger32_v_1020_9__g_ord_0_)
  );
  or_bb _340_ (
    .a(c_10_),
    .b(c_26_),
    .c(_m_genblock__src_b32s_merger32_v_1021_10__g_ord_1_)
  );
  and_bb _341_ (
    .a(c_10_),
    .b(c_26_),
    .c(_m_genblock__src_b32s_merger32_v_1021_10__g_ord_0_)
  );
  or_bb _342_ (
    .a(c_11_),
    .b(c_27_),
    .c(_m_genblock__src_b32s_merger32_v_1022_11__g_ord_1_)
  );
  and_bb _343_ (
    .a(c_11_),
    .b(c_27_),
    .c(_m_genblock__src_b32s_merger32_v_1022_11__g_ord_0_)
  );
  or_bb _344_ (
    .a(c_12_),
    .b(c_28_),
    .c(_m_genblock__src_b32s_merger32_v_1023_12__g_ord_1_)
  );
  and_bb _345_ (
    .a(c_12_),
    .b(c_28_),
    .c(_m_genblock__src_b32s_merger32_v_1023_12__g_ord_0_)
  );
  or_bb _346_ (
    .a(c_13_),
    .b(c_29_),
    .c(_m_genblock__src_b32s_merger32_v_1024_13__g_ord_1_)
  );
  and_bb _347_ (
    .a(c_13_),
    .b(c_29_),
    .c(_m_genblock__src_b32s_merger32_v_1024_13__g_ord_0_)
  );
  or_bb _348_ (
    .a(c_14_),
    .b(c_30_),
    .c(_m_genblock__src_b32s_merger32_v_1025_14__g_ord_1_)
  );
  and_bb _349_ (
    .a(c_14_),
    .b(c_30_),
    .c(_m_genblock__src_b32s_merger32_v_1025_14__g_ord_0_)
  );
  or_bb _350_ (
    .a(c_15_),
    .b(c_31_),
    .c(_m_genblock__src_b32s_merger32_v_1026_15__g_ord_1_)
  );
  and_bb _351_ (
    .a(c_15_),
    .b(c_31_),
    .c(_m_genblock__src_b32s_merger32_v_1026_15__g_ord_0_)
  );
  or_bb _352_ (
    .a(_m_genblock__src_b32s_merger32_v_1011_0__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1019_8__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_101_0__g_ord_1_)
  );
  and_bb _353_ (
    .a(_m_genblock__src_b32s_merger32_v_1011_0__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1019_8__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_101_0__g_ord_0_)
  );
  or_bb _354_ (
    .a(_m_genblock__src_b32s_merger32_v_1012_1__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1020_9__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_102_1__g_ord_1_)
  );
  and_bb _355_ (
    .a(_m_genblock__src_b32s_merger32_v_1012_1__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1020_9__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_102_1__g_ord_0_)
  );
  or_bb _356_ (
    .a(_m_genblock__src_b32s_merger32_v_1013_2__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1021_10__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_103_2__g_ord_1_)
  );
  and_bb _357_ (
    .a(_m_genblock__src_b32s_merger32_v_1013_2__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1021_10__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_103_2__g_ord_0_)
  );
  or_bb _358_ (
    .a(_m_genblock__src_b32s_merger32_v_1014_3__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1022_11__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_104_3__g_ord_1_)
  );
  and_bb _359_ (
    .a(_m_genblock__src_b32s_merger32_v_1014_3__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1022_11__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_104_3__g_ord_0_)
  );
  or_bb _360_ (
    .a(_m_genblock__src_b32s_merger32_v_1015_4__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1023_12__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_105_4__g_ord_1_)
  );
  and_bb _361_ (
    .a(_m_genblock__src_b32s_merger32_v_1015_4__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1023_12__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_105_4__g_ord_0_)
  );
  or_bb _362_ (
    .a(_m_genblock__src_b32s_merger32_v_1016_5__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1024_13__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_106_5__g_ord_1_)
  );
  and_bb _363_ (
    .a(_m_genblock__src_b32s_merger32_v_1016_5__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1024_13__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_106_5__g_ord_0_)
  );
  or_bb _364_ (
    .a(_m_genblock__src_b32s_merger32_v_1017_6__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1025_14__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_107_6__g_ord_1_)
  );
  and_bb _365_ (
    .a(_m_genblock__src_b32s_merger32_v_1017_6__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1025_14__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_107_6__g_ord_0_)
  );
  or_bb _366_ (
    .a(_m_genblock__src_b32s_merger32_v_1018_7__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1026_15__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_108_7__g_ord_1_)
  );
  and_bb _367_ (
    .a(_m_genblock__src_b32s_merger32_v_1018_7__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1026_15__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_108_7__g_ord_0_)
  );
  or_bb _368_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_101_0__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_105_4__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_)
  );
  and_bb _369_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_101_0__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_105_4__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_)
  );
  or_bb _370_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_102_1__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_106_5__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_)
  );
  and_bb _371_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_102_1__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_106_5__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_)
  );
  or_bb _372_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_103_2__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_107_6__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_)
  );
  and_bb _373_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_103_2__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_107_6__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_)
  );
  or_bb _374_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_104_3__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_108_7__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_)
  );
  and_bb _375_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_104_3__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_108_7__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_)
  );
  or_bb _376_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_3_)
  );
  and_bb _377_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_1_)
  );
  or_bb _378_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_2_)
  );
  and_bb _379_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_0_)
  );
  or_bb _380_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_2_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_3_),
    .c(b_11_)
  );
  and_bb _381_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_2_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_3_),
    .c(b_10_)
  );
  or_bb _382_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_0_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_1_),
    .c(b_9_)
  );
  and_bb _383_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_0_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_1_),
    .c(b_8_)
  );
  or_bb _384_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_3_)
  );
  and_bb _385_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_1_)
  );
  or_bb _386_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_2_)
  );
  and_bb _387_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_0_)
  );
  or_bb _388_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_2_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_3_),
    .c(b_15_)
  );
  and_bb _389_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_2_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_3_),
    .c(b_14_)
  );
  or_bb _390_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_0_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_1_),
    .c(b_13_)
  );
  and_bb _391_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_0_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_1_),
    .c(b_12_)
  );
  or_bb _392_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_101_0__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_105_4__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_)
  );
  and_bb _393_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_101_0__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_105_4__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_)
  );
  or_bb _394_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_102_1__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_106_5__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_)
  );
  and_bb _395_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_102_1__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_106_5__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_)
  );
  or_bb _396_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_103_2__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_107_6__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_)
  );
  and_bb _397_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_103_2__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_107_6__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_)
  );
  or_bb _398_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_104_3__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_108_7__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_)
  );
  and_bb _399_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_104_3__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_108_7__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_)
  );
  or_bb _400_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_3_)
  );
  and_bb _401_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_1_)
  );
  or_bb _402_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_2_)
  );
  and_bb _403_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_0_)
  );
  or_bb _404_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_2_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_3_),
    .c(b_3_)
  );
  and_bb _405_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_2_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_3_),
    .c(b_2_)
  );
  or_bb _406_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_0_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_1_),
    .c(b_1_)
  );
  and_bb _407_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_0_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_1_),
    .c(b_0_)
  );
  or_bb _408_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_3_)
  );
  and_bb _409_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_1_)
  );
  or_bb _410_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_2_)
  );
  and_bb _411_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_0_)
  );
  or_bb _412_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_2_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_3_),
    .c(b_7_)
  );
  and_bb _413_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_2_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_3_),
    .c(b_6_)
  );
  or_bb _414_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_0_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_1_),
    .c(b_5_)
  );
  and_bb _415_ (
    .a(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_0_),
    .b(_m_genblock__src_b32s_merger32_v_1327_0__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_1_),
    .c(b_4_)
  );
  or_bb _416_ (
    .a(_m_genblock__src_b32s_merger32_v_1011_0__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1019_8__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_101_0__g_ord_1_)
  );
  and_bb _417_ (
    .a(_m_genblock__src_b32s_merger32_v_1011_0__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1019_8__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_101_0__g_ord_0_)
  );
  or_bb _418_ (
    .a(_m_genblock__src_b32s_merger32_v_1012_1__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1020_9__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_102_1__g_ord_1_)
  );
  and_bb _419_ (
    .a(_m_genblock__src_b32s_merger32_v_1012_1__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1020_9__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_102_1__g_ord_0_)
  );
  or_bb _420_ (
    .a(_m_genblock__src_b32s_merger32_v_1013_2__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1021_10__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_103_2__g_ord_1_)
  );
  and_bb _421_ (
    .a(_m_genblock__src_b32s_merger32_v_1013_2__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1021_10__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_103_2__g_ord_0_)
  );
  or_bb _422_ (
    .a(_m_genblock__src_b32s_merger32_v_1014_3__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1022_11__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_104_3__g_ord_1_)
  );
  and_bb _423_ (
    .a(_m_genblock__src_b32s_merger32_v_1014_3__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1022_11__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_104_3__g_ord_0_)
  );
  or_bb _424_ (
    .a(_m_genblock__src_b32s_merger32_v_1015_4__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1023_12__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_105_4__g_ord_1_)
  );
  and_bb _425_ (
    .a(_m_genblock__src_b32s_merger32_v_1015_4__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1023_12__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_105_4__g_ord_0_)
  );
  or_bb _426_ (
    .a(_m_genblock__src_b32s_merger32_v_1016_5__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1024_13__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_106_5__g_ord_1_)
  );
  and_bb _427_ (
    .a(_m_genblock__src_b32s_merger32_v_1016_5__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1024_13__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_106_5__g_ord_0_)
  );
  or_bb _428_ (
    .a(_m_genblock__src_b32s_merger32_v_1017_6__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1025_14__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_107_6__g_ord_1_)
  );
  and_bb _429_ (
    .a(_m_genblock__src_b32s_merger32_v_1017_6__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1025_14__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_107_6__g_ord_0_)
  );
  or_bb _430_ (
    .a(_m_genblock__src_b32s_merger32_v_1018_7__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1026_15__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_108_7__g_ord_1_)
  );
  and_bb _431_ (
    .a(_m_genblock__src_b32s_merger32_v_1018_7__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1026_15__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_108_7__g_ord_0_)
  );
  or_bb _432_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_101_0__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_105_4__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_)
  );
  and_bb _433_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_101_0__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_105_4__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_)
  );
  or_bb _434_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_102_1__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_106_5__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_)
  );
  and_bb _435_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_102_1__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_106_5__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_)
  );
  or_bb _436_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_103_2__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_107_6__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_)
  );
  and_bb _437_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_103_2__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_107_6__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_)
  );
  or_bb _438_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_104_3__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_108_7__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_)
  );
  and_bb _439_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_104_3__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_108_7__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_)
  );
  or_bb _440_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_3_)
  );
  and_bb _441_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_1_)
  );
  or_bb _442_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_2_)
  );
  and_bb _443_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_0_)
  );
  or_bb _444_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_2_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_3_),
    .c(b_27_)
  );
  and_bb _445_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_2_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_3_),
    .c(b_26_)
  );
  or_bb _446_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_0_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_1_),
    .c(b_25_)
  );
  and_bb _447_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_0_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1333_0__m_c_1_),
    .c(b_24_)
  );
  or_bb _448_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_3_)
  );
  and_bb _449_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_1_)
  );
  or_bb _450_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_2_)
  );
  and_bb _451_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_0_)
  );
  or_bb _452_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_2_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_3_),
    .c(b_31_)
  );
  and_bb _453_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_2_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_3_),
    .c(b_30_)
  );
  or_bb _454_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_0_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_1_),
    .c(b_29_)
  );
  and_bb _455_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_0_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_1310_1__m_genblock__src_b32s_merger8_v_1334_1__m_c_1_),
    .c(b_28_)
  );
  or_bb _456_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_101_0__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_105_4__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_)
  );
  and_bb _457_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_101_0__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_105_4__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_)
  );
  or_bb _458_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_102_1__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_106_5__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_)
  );
  and_bb _459_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_102_1__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_106_5__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_)
  );
  or_bb _460_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_103_2__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_107_6__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_)
  );
  and_bb _461_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_103_2__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_107_6__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_)
  );
  or_bb _462_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_104_3__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_108_7__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_)
  );
  and_bb _463_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_104_3__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_108_7__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_)
  );
  or_bb _464_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_3_)
  );
  and_bb _465_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1030_1__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1032_3__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_1_)
  );
  or_bb _466_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_2_)
  );
  and_bb _467_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1029_0__g_ord_0_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1031_2__g_ord_0_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_0_)
  );
  or_bb _468_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_2_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_3_),
    .c(b_19_)
  );
  and_bb _469_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_2_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_3_),
    .c(b_18_)
  );
  or_bb _470_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_0_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_1_),
    .c(b_17_)
  );
  and_bb _471_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_0_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1333_0__m_c_1_),
    .c(b_16_)
  );
  or_bb _472_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_3_)
  );
  and_bb _473_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1030_1__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1032_3__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_1_)
  );
  or_bb _474_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_2_)
  );
  and_bb _475_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1029_0__g_ord_1_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1031_2__g_ord_1_),
    .c(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_0_)
  );
  or_bb _476_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_2_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_3_),
    .c(b_23_)
  );
  and_bb _477_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_2_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_3_),
    .c(b_22_)
  );
  or_bb _478_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_0_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_1_),
    .c(b_21_)
  );
  and_bb _479_ (
    .a(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_0_),
    .b(_m_genblock__src_b32s_merger32_v_1328_1__m_genblock__src_b32s_merger16_v_139_0__m_genblock__src_b32s_merger8_v_1334_1__m_c_1_),
    .c(b_20_)
  );
endmodule
