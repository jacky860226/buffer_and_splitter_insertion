module c432(N86,N69,N34,N92,N27,N43,N47,N79,N73,N24,N108,N1,N82,N56,N102,N17,N50,N63,N76,N99,N8,N11,N21,N30,N66,N89,N40,N53,N115,N14,N105,N60,N4,N95,N37,N112);
    wire new_Jinkela_wire_254;
    wire new_Jinkela_wire_644;
    wire new_Jinkela_wire_573;
    wire new_Jinkela_wire_364;
    wire new_Jinkela_wire_854;
    wire new_Jinkela_wire_269;
    wire new_Jinkela_wire_108;
    wire new_Jinkela_wire_904;
    wire new_Jinkela_wire_958;
    wire new_Jinkela_wire_328;
    wire new_Jinkela_wire_658;
    wire new_Jinkela_wire_182;
    wire new_Jinkela_wire_725;
    wire new_Jinkela_wire_925;
    wire new_Jinkela_wire_597;
    wire _112_;
    wire new_Jinkela_wire_397;
    wire new_Jinkela_wire_533;
    wire _041_;
    wire new_Jinkela_wire_957;
    wire new_Jinkela_wire_494;
    wire new_Jinkela_wire_888;
    wire new_Jinkela_wire_783;
    wire new_Jinkela_wire_80;
    wire new_Jinkela_wire_546;
    wire new_Jinkela_wire_319;
    wire new_Jinkela_wire_273;
    wire new_Jinkela_wire_286;
    wire new_Jinkela_wire_418;
    wire new_Jinkela_wire_799;
    wire new_Jinkela_wire_471;
    wire new_Jinkela_wire_860;
    wire new_Jinkela_wire_363;
    wire new_Jinkela_wire_464;
    wire new_Jinkela_wire_40;
    wire new_net_192;
    wire new_Jinkela_wire_83;
    wire new_Jinkela_wire_838;
    wire new_Jinkela_wire_604;
    wire new_Jinkela_wire_687;
    wire new_Jinkela_wire_707;
    wire new_Jinkela_wire_245;
    wire new_Jinkela_wire_519;
    wire new_Jinkela_wire_149;
    wire new_Jinkela_wire_753;
    wire _060_;
    wire _047_;
    wire new_Jinkela_wire_745;
    wire _088_;
    wire _002_;
    wire new_Jinkela_wire_715;
    wire new_Jinkela_wire_350;
    wire new_Jinkela_wire_259;
    wire new_Jinkela_wire_85;
    wire new_Jinkela_wire_105;
    wire new_Jinkela_wire_967;
    wire new_Jinkela_wire_884;
    wire new_Jinkela_wire_963;
    wire _013_;
    wire new_Jinkela_wire_613;
    wire new_Jinkela_wire_923;
    wire new_Jinkela_wire_822;
    wire new_Jinkela_wire_36;
    wire new_Jinkela_wire_557;
    wire new_Jinkela_wire_377;
    wire new_Jinkela_wire_316;
    wire new_Jinkela_wire_820;
    wire new_Jinkela_wire_812;
    wire new_Jinkela_wire_863;
    wire new_Jinkela_wire_736;
    wire _102_;
    wire new_Jinkela_wire_502;
    wire new_Jinkela_wire_551;
    wire new_Jinkela_wire_642;
    wire new_Jinkela_wire_94;
    wire new_Jinkela_wire_137;
    wire new_Jinkela_wire_620;
    wire new_Jinkela_wire_412;
    wire new_Jinkela_wire_44;
    wire new_Jinkela_wire_496;
    wire new_Jinkela_wire_910;
    wire new_Jinkela_wire_61;
    wire new_Jinkela_wire_279;
    wire new_Jinkela_wire_780;
    wire new_Jinkela_wire_91;
    wire new_Jinkela_wire_486;
    wire new_Jinkela_wire_384;
    wire new_Jinkela_wire_973;
    wire new_Jinkela_wire_585;
    wire _096_;
    wire new_Jinkela_wire_299;
    wire new_Jinkela_wire_101;
    wire new_Jinkela_wire_664;
    wire new_Jinkela_wire_26;
    wire new_Jinkela_wire_666;
    wire new_Jinkela_wire_897;
    wire new_Jinkela_wire_547;
    wire new_Jinkela_wire_775;
    wire new_Jinkela_wire_928;
    wire new_Jinkela_wire_442;
    wire new_Jinkela_wire_869;
    wire new_Jinkela_wire_883;
    wire new_Jinkela_wire_296;
    wire new_Jinkela_wire_488;
    wire new_Jinkela_wire_595;
    wire new_Jinkela_wire_968;
    wire new_Jinkela_wire_970;
    wire new_Jinkela_wire_437;
    wire new_Jinkela_wire_62;
    wire new_Jinkela_wire_726;
    wire new_Jinkela_wire_571;
    wire new_Jinkela_wire_383;
    wire new_Jinkela_wire_335;
    wire new_Jinkela_wire_554;
    wire new_Jinkela_wire_825;
    wire new_Jinkela_wire_95;
    wire _093_;
    wire new_Jinkela_wire_294;
    wire _083_;
    wire new_Jinkela_wire_565;
    wire new_Jinkela_wire_435;
    wire new_Jinkela_wire_460;
    wire _059_;
    wire new_Jinkela_wire_684;
    wire _070_;
    wire new_Jinkela_wire_141;
    wire new_Jinkela_wire_317;
    wire new_Jinkela_wire_416;
    wire _069_;
    wire new_Jinkela_wire_25;
    wire new_Jinkela_wire_12;
    wire new_Jinkela_wire_476;
    wire _100_;
    wire new_Jinkela_wire_24;
    wire new_Jinkela_wire_168;
    wire new_Jinkela_wire_256;
    wire new_Jinkela_wire_683;
    wire _005_;
    wire new_Jinkela_wire_42;
    wire _034_;
    wire new_Jinkela_wire_638;
    wire new_Jinkela_wire_929;
    wire new_Jinkela_wire_621;
    wire new_Jinkela_wire_371;
    wire new_Jinkela_wire_179;
    wire new_Jinkela_wire_19;
    wire new_Jinkela_wire_730;
    wire new_Jinkela_wire_750;
    wire _025_;
    wire new_Jinkela_wire_443;
    wire new_Jinkela_wire_81;
    wire new_Jinkela_wire_912;
    wire new_Jinkela_wire_506;
    wire new_Jinkela_wire_67;
    wire new_Jinkela_wire_239;
    wire new_Jinkela_wire_543;
    wire new_Jinkela_wire_826;
    wire new_Jinkela_wire_865;
    wire new_Jinkela_wire_537;
    wire new_Jinkela_wire_837;
    wire new_Jinkela_wire_47;
    wire _022_;
    wire new_Jinkela_wire_440;
    wire new_Jinkela_wire_807;
    wire new_Jinkela_wire_705;
    wire new_Jinkela_wire_461;
    wire new_Jinkela_wire_176;
    wire new_Jinkela_wire_670;
    wire new_Jinkela_wire_153;
    wire _103_;
    wire new_Jinkela_wire_829;
    wire new_Jinkela_wire_614;
    wire new_Jinkela_wire_352;
    wire new_Jinkela_wire_560;
    wire new_Jinkela_wire_173;
    wire new_Jinkela_wire_951;
    wire new_Jinkela_wire_722;
    wire new_Jinkela_wire_311;
    wire new_Jinkela_wire_667;
    wire new_Jinkela_wire_765;
    wire new_Jinkela_wire_616;
    wire new_Jinkela_wire_142;
    wire new_Jinkela_wire_470;
    wire new_Jinkela_wire_439;
    wire new_Jinkela_wire_107;
    wire new_Jinkela_wire_937;
    wire _055_;
    wire new_Jinkela_wire_728;
    wire new_Jinkela_wire_28;
    wire _004_;
    wire new_Jinkela_wire_9;
    wire _029_;
    wire new_Jinkela_wire_490;
    wire new_Jinkela_wire_767;
    wire new_Jinkela_wire_971;
    wire new_Jinkela_wire_277;
    wire new_Jinkela_wire_600;
    wire new_Jinkela_wire_760;
    wire new_Jinkela_wire_73;
    wire new_Jinkela_wire_20;
    wire new_Jinkela_wire_4;
    wire new_Jinkela_wire_698;
    wire _104_;
    wire new_Jinkela_wire_313;
    wire _049_;
    wire new_Jinkela_wire_399;
    wire new_Jinkela_wire_692;
    wire new_Jinkela_wire_743;
    wire new_Jinkela_wire_157;
    wire new_Jinkela_wire_732;
    wire new_Jinkela_wire_322;
    wire new_Jinkela_wire_300;
    wire new_Jinkela_wire_934;
    wire new_Jinkela_wire_729;
    wire new_Jinkela_wire_493;
    wire new_Jinkela_wire_394;
    wire new_Jinkela_wire_668;
    wire new_Jinkela_wire_257;
    wire new_Jinkela_wire_2;
    wire new_Jinkela_wire_669;
    wire new_Jinkela_wire_909;
    wire new_Jinkela_wire_931;
    wire new_Jinkela_wire_124;
    wire new_Jinkela_wire_131;
    wire _015_;
    wire new_Jinkela_wire_927;
    wire new_Jinkela_wire_233;
    wire new_Jinkela_wire_22;
    wire new_Jinkela_wire_230;
    wire new_Jinkela_wire_824;
    wire _099_;
    wire new_Jinkela_wire_754;
    wire new_Jinkela_wire_991;
    wire new_Jinkela_wire_481;
    wire new_Jinkela_wire_288;
    wire new_Jinkela_wire_526;
    wire new_Jinkela_wire_431;
    wire new_Jinkela_wire_813;
    wire _028_;
    wire new_Jinkela_wire_579;
    wire new_Jinkela_wire_129;
    wire new_Jinkela_wire_497;
    wire new_Jinkela_wire_539;
    wire new_Jinkela_wire_156;
    wire new_Jinkela_wire_167;
    wire new_Jinkela_wire_321;
    wire new_Jinkela_wire_241;
    wire new_Jinkela_wire_78;
    wire new_Jinkela_wire_160;
    wire _061_;
    wire new_Jinkela_wire_276;
    wire new_Jinkela_wire_771;
    wire new_Jinkela_wire_665;
    wire new_Jinkela_wire_814;
    wire new_Jinkela_wire_741;
    wire new_Jinkela_wire_366;
    wire new_Jinkela_wire_877;
    wire new_Jinkela_wire_672;
    wire new_Jinkela_wire_886;
    wire new_Jinkela_wire_336;
    wire new_Jinkela_wire_649;
    wire new_Jinkela_wire_333;
    wire new_Jinkela_wire_5;
    wire new_Jinkela_wire_37;
    wire new_Jinkela_wire_369;
    wire new_Jinkela_wire_862;
    wire _033_;
    wire new_Jinkela_wire_201;
    wire new_Jinkela_wire_529;
    wire new_Jinkela_wire_466;
    wire new_Jinkela_wire_287;
    wire _105_;
    wire _046_;
    wire _064_;
    wire new_Jinkela_wire_779;
    wire _074_;
    wire new_Jinkela_wire_680;
    wire _027_;
    wire new_Jinkela_wire_757;
    wire new_Jinkela_wire_940;
    wire new_Jinkela_wire_514;
    wire new_Jinkela_wire_441;
    wire new_Jinkela_wire_203;
    wire new_Jinkela_wire_425;
    wire new_Jinkela_wire_33;
    wire new_Jinkela_wire_892;
    wire new_Jinkela_wire_656;
    wire new_Jinkela_wire_298;
    wire new_Jinkela_wire_411;
    wire new_Jinkela_wire_778;
    wire new_Jinkela_wire_641;
    wire new_Jinkela_wire_103;
    wire new_Jinkela_wire_719;
    wire new_Jinkela_wire_663;
    wire _019_;
    wire _114_;
    wire new_Jinkela_wire_458;
    wire new_Jinkela_wire_362;
    wire new_Jinkela_wire_845;
    wire new_Jinkela_wire_15;
    wire new_Jinkela_wire_463;
    wire new_Jinkela_wire_893;
    wire new_Jinkela_wire_240;
    wire new_Jinkela_wire_122;
    wire new_Jinkela_wire_184;
    wire new_Jinkela_wire_657;
    wire new_Jinkela_wire_903;
    wire new_Jinkela_wire_320;
    wire new_Jinkela_wire_501;
    wire _076_;
    wire new_Jinkela_wire_652;
    wire new_Jinkela_wire_208;
    wire new_Jinkela_wire_868;
    wire new_Jinkela_wire_889;
    wire _018_;
    wire _116_;
    wire new_Jinkela_wire_111;
    wire new_Jinkela_wire_206;
    wire new_Jinkela_wire_54;
    wire new_net_0;
    wire new_Jinkela_wire_408;
    wire new_Jinkela_wire_341;
    wire _073_;
    wire _052_;
    wire _021_;
    wire new_Jinkela_wire_358;
    wire new_Jinkela_wire_782;
    wire new_Jinkela_wire_52;
    wire new_Jinkela_wire_563;
    wire new_Jinkela_wire_651;
    wire new_Jinkela_wire_249;
    wire new_Jinkela_wire_21;
    wire new_Jinkela_wire_438;
    wire new_Jinkela_wire_224;
    wire new_Jinkela_wire_500;
    wire new_Jinkela_wire_661;
    wire new_Jinkela_wire_267;
    wire new_Jinkela_wire_354;
    wire new_Jinkela_wire_818;
    wire new_Jinkela_wire_283;
    wire new_Jinkela_wire_290;
    wire new_Jinkela_wire_473;
    wire new_Jinkela_wire_836;
    wire new_Jinkela_wire_784;
    wire new_Jinkela_wire_590;
    wire _051_;
    wire new_Jinkela_wire_855;
    wire new_Jinkela_wire_218;
    wire new_Jinkela_wire_39;
    wire new_Jinkela_wire_534;
    wire new_Jinkela_wire_787;
    wire new_Jinkela_wire_289;
    wire new_Jinkela_wire_152;
    wire new_Jinkela_wire_615;
    wire new_Jinkela_wire_27;
    wire new_Jinkela_wire_197;
    wire new_Jinkela_wire_297;
    wire new_Jinkela_wire_704;
    wire new_Jinkela_wire_878;
    wire new_Jinkela_wire_856;
    wire new_Jinkela_wire_980;
    wire _068_;
    wire new_Jinkela_wire_177;
    wire new_Jinkela_wire_365;
    wire new_Jinkela_wire_517;
    wire new_Jinkela_wire_98;
    wire new_Jinkela_wire_71;
    wire new_Jinkela_wire_35;
    wire _075_;
    wire new_Jinkela_wire_811;
    wire new_Jinkela_wire_516;
    wire new_Jinkela_wire_242;
    wire new_Jinkela_wire_381;
    wire new_Jinkela_wire_395;
    wire new_Jinkela_wire_647;
    wire new_Jinkela_wire_400;
    wire new_Jinkela_wire_776;
    wire _030_;
    wire new_Jinkela_wire_405;
    wire new_Jinkela_wire_181;
    wire new_Jinkela_wire_550;
    wire new_Jinkela_wire_467;
    wire new_Jinkela_wire_885;
    wire new_Jinkela_wire_188;
    wire new_Jinkela_wire_907;
    wire new_Jinkela_wire_274;
    wire _084_;
    wire new_Jinkela_wire_57;
    wire new_Jinkela_wire_404;
    wire new_Jinkela_wire_752;
    wire _063_;
    wire new_Jinkela_wire_653;
    wire new_Jinkela_wire_433;
    wire new_Jinkela_wire_75;
    wire new_Jinkela_wire_415;
    wire new_Jinkela_wire_356;
    wire new_Jinkela_wire_452;
    wire new_Jinkela_wire_988;
    wire new_Jinkela_wire_150;
    wire new_Jinkela_wire_66;
    wire new_Jinkela_wire_549;
    wire new_Jinkela_wire_342;
    wire new_Jinkela_wire_520;
    wire new_Jinkela_wire_881;
    wire new_Jinkela_wire_527;
    wire new_Jinkela_wire_43;
    wire new_Jinkela_wire_270;
    wire new_Jinkela_wire_675;
    wire new_Jinkela_wire_828;
    wire new_Jinkela_wire_401;
    wire _078_;
    wire new_Jinkela_wire_890;
    wire new_Jinkela_wire_749;
    wire new_Jinkela_wire_16;
    wire new_Jinkela_wire_899;
    wire new_Jinkela_wire_55;
    wire new_Jinkela_wire_576;
    wire new_Jinkela_wire_449;
    wire new_Jinkela_wire_739;
    wire new_Jinkela_wire_718;
    wire new_Jinkela_wire_528;
    wire new_Jinkela_wire_268;
    wire new_Jinkela_wire_234;
    wire new_Jinkela_wire_121;
    wire new_Jinkela_wire_872;
    wire _086_;
    wire new_Jinkela_wire_632;
    wire new_Jinkela_wire_275;
    wire _016_;
    wire new_Jinkela_wire_391;
    wire new_Jinkela_wire_53;
    wire new_Jinkela_wire_413;
    wire new_Jinkela_wire_211;
    wire new_Jinkela_wire_717;
    wire new_Jinkela_wire_567;
    wire new_Jinkela_wire_232;
    wire new_Jinkela_wire_262;
    wire new_Jinkela_wire_174;
    wire new_Jinkela_wire_450;
    wire new_Jinkela_wire_330;
    wire new_Jinkela_wire_186;
    wire new_Jinkela_wire_694;
    wire new_Jinkela_wire_627;
    wire new_Jinkela_wire_504;
    wire new_Jinkela_wire_617;
    wire new_Jinkela_wire_523;
    wire new_Jinkela_wire_355;
    wire new_Jinkela_wire_695;
    wire new_Jinkela_wire_582;
    wire new_Jinkela_wire_236;
    wire new_Jinkela_wire_212;
    wire new_Jinkela_wire_591;
    wire _008_;
    wire new_Jinkela_wire_357;
    wire new_Jinkela_wire_746;
    wire new_Jinkela_wire_662;
    wire new_Jinkela_wire_307;
    wire new_Jinkela_wire_90;
    wire new_Jinkela_wire_637;
    wire new_Jinkela_wire_802;
    wire _035_;
    wire new_Jinkela_wire_938;
    wire new_Jinkela_wire_915;
    wire new_Jinkela_wire_324;
    wire new_Jinkela_wire_610;
    wire new_Jinkela_wire_34;
    wire new_Jinkela_wire_524;
    wire _042_;
    wire new_Jinkela_wire_788;
    wire new_Jinkela_wire_594;
    wire new_Jinkela_wire_110;
    wire new_Jinkela_wire_960;
    wire new_Jinkela_wire_309;
    wire new_Jinkela_wire_629;
    wire new_Jinkela_wire_612;
    wire _062_;
    wire new_Jinkela_wire_712;
    wire new_Jinkela_wire_636;
    wire new_Jinkela_wire_329;
    wire new_Jinkela_wire_162;
    wire new_Jinkela_wire_990;
    wire new_Jinkela_wire_99;
    wire new_Jinkela_wire_193;
    wire new_Jinkela_wire_45;
    wire new_Jinkela_wire_260;
    wire new_Jinkela_wire_271;
    wire new_Jinkela_wire_195;
    wire new_Jinkela_wire_966;
    wire new_Jinkela_wire_608;
    wire new_Jinkela_wire_281;
    wire new_Jinkela_wire_936;
    wire new_Jinkela_wire_180;
    wire new_Jinkela_wire_301;
    wire new_Jinkela_wire_390;
    wire new_Jinkela_wire_564;
    wire new_Jinkela_wire_225;
    wire new_Jinkela_wire_100;
    wire new_Jinkela_wire_92;
    wire new_Jinkela_wire_902;
    wire new_Jinkela_wire_633;
    wire new_Jinkela_wire_685;
    wire new_Jinkela_wire_426;
    wire new_net_198;
    wire _095_;
    wire new_Jinkela_wire_766;
    wire new_Jinkela_wire_138;
    wire new_Jinkela_wire_983;
    wire new_Jinkela_wire_200;
    wire new_Jinkela_wire_86;
    wire new_Jinkela_wire_46;
    wire new_Jinkela_wire_378;
    wire new_Jinkela_wire_688;
    wire new_Jinkela_wire_791;
    wire new_Jinkela_wire_130;
    wire new_Jinkela_wire_145;
    wire new_Jinkela_wire_387;
    wire new_Jinkela_wire_974;
    wire new_Jinkela_wire_265;
    wire new_Jinkela_wire_941;
    wire new_Jinkela_wire_382;
    wire new_Jinkela_wire_172;
    wire new_Jinkela_wire_148;
    wire new_Jinkela_wire_104;
    wire new_Jinkela_wire_136;
    wire new_Jinkela_wire_584;
    wire new_Jinkela_wire_723;
    wire new_Jinkela_wire_536;
    wire new_Jinkela_wire_898;
    wire new_Jinkela_wire_199;
    wire new_Jinkela_wire_674;
    wire new_Jinkela_wire_38;
    wire new_Jinkela_wire_511;
    wire new_Jinkela_wire_918;
    wire _012_;
    wire new_Jinkela_wire_375;
    wire new_Jinkela_wire_926;
    wire new_Jinkela_wire_492;
    wire new_Jinkela_wire_981;
    wire new_Jinkela_wire_247;
    wire new_Jinkela_wire_727;
    wire new_Jinkela_wire_79;
    wire new_Jinkela_wire_556;
    wire new_Jinkela_wire_593;
    wire _072_;
    wire new_Jinkela_wire_650;
    wire new_Jinkela_wire_163;
    wire new_Jinkela_wire_919;
    wire new_Jinkela_wire_304;
    wire new_Jinkela_wire_815;
    wire new_Jinkela_wire_733;
    wire new_Jinkela_wire_522;
    wire new_Jinkela_wire_396;
    wire new_Jinkela_wire_572;
    wire new_Jinkela_wire_558;
    wire new_Jinkela_wire_59;
    wire new_Jinkela_wire_69;
    wire new_Jinkela_wire_171;
    wire new_Jinkela_wire_459;
    wire new_Jinkela_wire_348;
    wire new_Jinkela_wire_204;
    wire new_Jinkela_wire_315;
    wire new_Jinkela_wire_830;
    wire new_Jinkela_wire_166;
    wire new_Jinkela_wire_468;
    wire new_Jinkela_wire_89;
    wire new_Jinkela_wire_821;
    wire new_Jinkela_wire_731;
    wire new_Jinkela_wire_18;
    wire new_Jinkela_wire_796;
    wire _020_;
    wire new_Jinkela_wire_589;
    wire new_Jinkela_wire_427;
    wire new_Jinkela_wire_834;
    wire new_Jinkela_wire_606;
    wire new_Jinkela_wire_559;
    wire new_Jinkela_wire_871;
    wire new_Jinkela_wire_693;
    wire new_Jinkela_wire_303;
    wire new_Jinkela_wire_624;
    wire new_Jinkela_wire_291;
    wire new_Jinkela_wire_535;
    wire new_Jinkela_wire_388;
    wire new_Jinkela_wire_487;
    wire new_Jinkela_wire_510;
    wire new_Jinkela_wire_456;
    wire new_Jinkela_wire_607;
    wire new_Jinkela_wire_192;
    wire new_Jinkela_wire_102;
    wire _003_;
    wire new_Jinkela_wire_223;
    wire new_Jinkela_wire_975;
    wire new_Jinkela_wire_920;
    wire new_Jinkela_wire_93;
    wire new_Jinkela_wire_602;
    wire new_Jinkela_wire_202;
    wire new_Jinkela_wire_993;
    wire new_Jinkela_wire_774;
    wire _071_;
    wire _024_;
    wire new_Jinkela_wire_346;
    wire _031_;
    wire new_Jinkela_wire_841;
    wire _054_;
    wire new_Jinkela_wire_772;
    wire new_Jinkela_wire_697;
    wire new_Jinkela_wire_88;
    wire _111_;
    wire new_Jinkela_wire_552;
    wire new_Jinkela_wire_842;
    wire _066_;
    wire _045_;
    wire new_Jinkela_wire_942;
    wire new_Jinkela_wire_143;
    wire new_Jinkela_wire_962;
    wire _011_;
    wire new_Jinkela_wire_263;
    wire _097_;
    wire _050_;
    wire _038_;
    wire new_Jinkela_wire_803;
    wire new_Jinkela_wire_58;
    wire new_Jinkela_wire_513;
    wire new_Jinkela_wire_790;
    wire new_Jinkela_wire_716;
    wire new_Jinkela_wire_380;
    wire new_Jinkela_wire_611;
    wire new_Jinkela_wire_943;
    wire new_Jinkela_wire_569;
    wire new_net_196;
    wire new_Jinkela_wire_161;
    wire new_Jinkela_wire_338;
    wire new_Jinkela_wire_3;
    wire new_Jinkela_wire_489;
    wire _082_;
    wire new_Jinkela_wire_495;
    wire new_Jinkela_wire_959;
    wire new_Jinkela_wire_849;
    wire new_Jinkela_wire_508;
    wire new_Jinkela_wire_965;
    wire new_Jinkela_wire_955;
    wire new_Jinkela_wire_389;
    wire new_Jinkela_wire_701;
    wire new_Jinkela_wire_708;
    wire _053_;
    wire new_Jinkela_wire_798;
    wire new_Jinkela_wire_630;
    wire new_Jinkela_wire_374;
    wire new_Jinkela_wire_419;
    wire new_Jinkela_wire_994;
    wire new_Jinkela_wire_68;
    wire _087_;
    wire new_Jinkela_wire_954;
    wire new_Jinkela_wire_911;
    wire new_Jinkela_wire_407;
    wire new_Jinkela_wire_785;
    wire new_Jinkela_wire_72;
    wire new_Jinkela_wire_169;
    wire new_Jinkela_wire_671;
    wire new_Jinkela_wire_677;
    wire new_Jinkela_wire_77;
    wire new_Jinkela_wire_220;
    wire new_Jinkela_wire_221;
    wire new_Jinkela_wire_545;
    wire new_Jinkela_wire_222;
    wire new_Jinkela_wire_454;
    wire new_Jinkela_wire_312;
    wire new_Jinkela_wire_231;
    wire new_Jinkela_wire_499;
    wire new_Jinkela_wire_158;
    wire new_Jinkela_wire_525;
    wire new_Jinkela_wire_343;
    wire new_Jinkela_wire_14;
    wire new_Jinkela_wire_462;
    wire new_Jinkela_wire_905;
    wire new_Jinkela_wire_740;
    wire new_Jinkela_wire_844;
    wire new_Jinkela_wire_972;
    wire new_Jinkela_wire_659;
    wire new_Jinkela_wire_882;
    wire new_Jinkela_wire_410;
    wire new_Jinkela_wire_906;
    wire new_Jinkela_wire_846;
    wire new_Jinkela_wire_518;
    wire new_Jinkela_wire_568;
    wire new_Jinkela_wire_566;
    wire new_Jinkela_wire_424;
    wire new_net_194;
    wire new_Jinkela_wire_429;
    wire new_Jinkela_wire_474;
    wire new_Jinkela_wire_989;
    wire new_Jinkela_wire_323;
    wire new_Jinkela_wire_503;
    wire new_Jinkela_wire_592;
    wire new_Jinkela_wire_453;
    wire new_Jinkela_wire_742;
    wire new_Jinkela_wire_952;
    wire new_Jinkela_wire_540;
    wire new_Jinkela_wire_485;
    wire new_Jinkela_wire_605;
    wire new_Jinkela_wire_118;
    wire new_Jinkela_wire_116;
    wire new_Jinkela_wire_331;
    wire new_Jinkela_wire_961;
    wire new_Jinkela_wire_689;
    wire new_Jinkela_wire_367;
    wire new_Jinkela_wire_370;
    wire new_Jinkela_wire_479;
    wire new_Jinkela_wire_120;
    wire new_Jinkela_wire_953;
    wire _081_;
    wire new_Jinkela_wire_714;
    wire new_Jinkela_wire_808;
    wire new_Jinkela_wire_574;
    wire new_Jinkela_wire_155;
    wire new_Jinkela_wire_702;
    wire _023_;
    wire new_Jinkela_wire_340;
    wire new_Jinkela_wire_251;
    wire new_Jinkela_wire_762;
    wire new_Jinkela_wire_544;
    wire new_Jinkela_wire_678;
    wire new_Jinkela_wire_421;
    wire _014_;
    wire new_Jinkela_wire_134;
    wire new_Jinkela_wire_924;
    wire new_Jinkela_wire_521;
    wire new_Jinkela_wire_696;
    wire new_Jinkela_wire_922;
    wire new_Jinkela_wire_840;
    wire new_Jinkela_wire_713;
    wire new_Jinkela_wire_393;
    wire new_Jinkela_wire_709;
    wire new_Jinkela_wire_217;
    wire new_Jinkela_wire_948;
    wire new_Jinkela_wire_337;
    wire new_Jinkela_wire_164;
    wire new_Jinkela_wire_97;
    wire new_Jinkela_wire_229;
    wire new_Jinkela_wire_376;
    wire _043_;
    wire new_Jinkela_wire_209;
    wire new_Jinkela_wire_70;
    wire new_Jinkela_wire_261;
    wire new_Jinkela_wire_690;
    wire new_Jinkela_wire_932;
    wire new_Jinkela_wire_17;
    wire _113_;
    wire _106_;
    wire new_Jinkela_wire_349;
    wire new_Jinkela_wire_41;
    wire new_Jinkela_wire_398;
    wire new_Jinkela_wire_859;
    wire new_Jinkela_wire_843;
    wire new_Jinkela_wire_634;
    wire new_Jinkela_wire_777;
    wire new_Jinkela_wire_625;
    wire _037_;
    wire new_Jinkela_wire_848;
    wire new_Jinkela_wire_686;
    wire new_Jinkela_wire_447;
    wire new_Jinkela_wire_619;
    wire new_Jinkela_wire_248;
    wire new_Jinkela_wire_455;
    wire new_Jinkela_wire_876;
    wire new_Jinkela_wire_29;
    wire new_Jinkela_wire_480;
    wire new_Jinkela_wire_673;
    wire new_Jinkela_wire_509;
    wire new_Jinkela_wire_755;
    wire new_Jinkela_wire_189;
    wire new_Jinkela_wire_244;
    wire new_Jinkela_wire_831;
    wire new_Jinkela_wire_792;
    wire new_Jinkela_wire_930;
    wire new_Jinkela_wire_457;
    wire _115_;
    wire new_Jinkela_wire_475;
    wire new_Jinkela_wire_63;
    wire new_Jinkela_wire_280;
    wire new_Jinkela_wire_850;
    wire _044_;
    wire _089_;
    wire new_Jinkela_wire_361;
    wire new_Jinkela_wire_7;
    wire _067_;
    wire new_Jinkela_wire_596;
    wire new_Jinkela_wire_326;
    wire new_Jinkela_wire_332;
    wire new_Jinkela_wire_507;
    wire new_Jinkela_wire_870;
    wire new_Jinkela_wire_139;
    wire new_Jinkela_wire_618;
    wire new_Jinkela_wire_403;
    wire _017_;
    wire new_Jinkela_wire_979;
    wire _085_;
    wire new_Jinkela_wire_933;
    wire new_Jinkela_wire_159;
    wire new_Jinkela_wire_548;
    wire new_Jinkela_wire_215;
    wire new_Jinkela_wire_916;
    wire new_Jinkela_wire_113;
    wire new_Jinkela_wire_982;
    wire new_Jinkela_wire_964;
    wire new_Jinkela_wire_491;
    wire new_Jinkela_wire_451;
    wire new_Jinkela_wire_278;
    wire new_Jinkela_wire_724;
    wire new_Jinkela_wire_851;
    wire new_Jinkela_wire_420;
    wire new_Jinkela_wire_379;
    wire new_Jinkela_wire_112;
    wire new_Jinkela_wire_805;
    wire new_Jinkela_wire_711;
    wire new_Jinkela_wire_985;
    wire new_Jinkela_wire_465;
    wire new_Jinkela_wire_976;
    wire new_Jinkela_wire_969;
    wire new_Jinkela_wire_921;
    wire new_Jinkela_wire_578;
    wire new_Jinkela_wire_896;
    wire new_Jinkela_wire_703;
    wire new_Jinkela_wire_676;
    wire new_Jinkela_wire_583;
    wire new_Jinkela_wire_417;
    wire new_Jinkela_wire_809;
    wire _092_;
    wire new_Jinkela_wire_827;
    wire new_Jinkela_wire_531;
    wire new_Jinkela_wire_178;
    wire new_Jinkela_wire_235;
    wire new_Jinkela_wire_987;
    wire new_Jinkela_wire_30;
    wire new_Jinkela_wire_735;
    wire new_Jinkela_wire_858;
    wire new_Jinkela_wire_125;
    wire new_Jinkela_wire_561;
    wire new_Jinkela_wire_737;
    wire new_Jinkela_wire_6;
    wire new_Jinkela_wire_839;
    wire new_Jinkela_wire_699;
    wire new_Jinkela_wire_144;
    wire new_Jinkela_wire_945;
    wire _036_;
    wire new_Jinkela_wire_255;
    wire new_Jinkela_wire_901;
    wire _056_;
    wire new_Jinkela_wire_285;
    wire new_Jinkela_wire_243;
    wire new_Jinkela_wire_214;
    wire new_Jinkela_wire_747;
    wire new_Jinkela_wire_853;
    wire new_Jinkela_wire_586;
    wire new_Jinkela_wire_432;
    wire new_Jinkela_wire_655;
    wire new_Jinkela_wire_914;
    wire new_Jinkela_wire_258;
    wire new_Jinkela_wire_402;
    wire new_Jinkela_wire_359;
    wire new_Jinkela_wire_345;
    wire new_Jinkela_wire_132;
    wire new_Jinkela_wire_588;
    wire new_Jinkela_wire_353;
    wire new_Jinkela_wire_334;
    wire new_Jinkela_wire_682;
    wire new_Jinkela_wire_65;
    wire _094_;
    wire _107_;
    wire new_Jinkela_wire_226;
    wire new_Jinkela_wire_64;
    wire new_Jinkela_wire_327;
    wire new_Jinkela_wire_23;
    wire _101_;
    wire new_Jinkela_wire_8;
    wire new_Jinkela_wire_133;
    wire new_Jinkela_wire_681;
    wire new_Jinkela_wire_804;
    wire _026_;
    wire new_Jinkela_wire_306;
    wire new_Jinkela_wire_250;
    wire new_Jinkela_wire_744;
    wire new_Jinkela_wire_873;
    wire _091_;
    wire new_Jinkela_wire_789;
    wire new_Jinkela_wire_700;
    wire new_Jinkela_wire_875;
    wire new_Jinkela_wire_756;
    wire new_Jinkela_wire_833;
    wire new_Jinkela_wire_82;
    wire new_Jinkela_wire_887;
    wire new_Jinkela_wire_764;
    wire new_Jinkela_wire_832;
    wire new_Jinkela_wire_917;
    wire new_Jinkela_wire_623;
    wire new_Jinkela_wire_117;
    wire new_Jinkela_wire_515;
    wire new_Jinkela_wire_154;
    wire new_Jinkela_wire_469;
    wire new_Jinkela_wire_183;
    wire new_Jinkela_wire_984;
    wire new_Jinkela_wire_580;
    wire new_Jinkela_wire_628;
    wire new_Jinkela_wire_165;
    wire new_Jinkela_wire_96;
    wire new_Jinkela_wire_532;
    wire new_Jinkela_wire_422;
    wire new_Jinkela_wire_835;
    wire new_Jinkela_wire_570;
    wire new_Jinkela_wire_227;
    wire new_Jinkela_wire_867;
    wire new_Jinkela_wire_127;
    wire new_Jinkela_wire_126;
    wire new_Jinkela_wire_436;
    wire new_Jinkela_wire_986;
    wire new_Jinkela_wire_196;
    wire new_Jinkela_wire_386;
    wire new_Jinkela_wire_444;
    wire new_Jinkela_wire_228;
    wire new_Jinkela_wire_555;
    wire new_Jinkela_wire_541;
    wire new_Jinkela_wire_360;
    wire _032_;
    wire new_Jinkela_wire_76;
    wire new_Jinkela_wire_119;
    wire new_Jinkela_wire_295;
    wire _057_;
    wire new_Jinkela_wire_446;
    wire new_Jinkela_wire_74;
    wire new_Jinkela_wire_190;
    wire new_Jinkela_wire_87;
    wire new_Jinkela_wire_423;
    wire new_Jinkela_wire_477;
    wire _058_;
    wire new_Jinkela_wire_49;
    wire new_Jinkela_wire_318;
    wire new_Jinkela_wire_368;
    wire _080_;
    wire new_Jinkela_wire_706;
    wire new_Jinkela_wire_562;
    wire new_Jinkela_wire_147;
    wire new_Jinkela_wire_654;
    wire new_Jinkela_wire_880;
    wire new_Jinkela_wire_770;
    wire new_Jinkela_wire_879;
    wire _000_;
    wire new_Jinkela_wire_643;
    wire new_Jinkela_wire_816;
    wire new_Jinkela_wire_106;
    wire new_Jinkela_wire_428;
    wire new_Jinkela_wire_817;
    wire new_Jinkela_wire_763;
    wire new_Jinkela_wire_170;
    wire new_Jinkela_wire_56;
    wire new_Jinkela_wire_645;
    wire new_Jinkela_wire_648;
    wire _006_;
    wire new_Jinkela_wire_852;
    wire new_Jinkela_wire_13;
    wire new_Jinkela_wire_385;
    wire new_Jinkela_wire_373;
    wire new_Jinkela_wire_944;
    wire _039_;
    wire new_Jinkela_wire_115;
    wire new_Jinkela_wire_185;
    wire new_Jinkela_wire_205;
    wire new_Jinkela_wire_140;
    wire new_Jinkela_wire_50;
    wire new_Jinkela_wire_60;
    wire new_Jinkela_wire_891;
    wire new_Jinkela_wire_1;
    wire _048_;
    wire new_Jinkela_wire_31;
    wire new_Jinkela_wire_598;
    wire new_Jinkela_wire_679;
    wire new_Jinkela_wire_175;
    wire new_Jinkela_wire_738;
    wire new_Jinkela_wire_847;
    wire new_Jinkela_wire_587;
    wire new_Jinkela_wire_748;
    wire new_Jinkela_wire_751;
    wire new_Jinkela_wire_32;
    wire new_Jinkela_wire_786;
    wire new_Jinkela_wire_512;
    wire new_Jinkela_wire_325;
    wire new_Jinkela_wire_210;
    wire new_Jinkela_wire_483;
    wire new_Jinkela_wire_484;
    wire new_Jinkela_wire_640;
    wire new_Jinkela_wire_823;
    wire new_Jinkela_wire_913;
    wire new_Jinkela_wire_977;
    wire new_Jinkela_wire_935;
    wire new_Jinkela_wire_794;
    wire new_Jinkela_wire_956;
    wire new_Jinkela_wire_434;
    wire _077_;
    wire new_Jinkela_wire_252;
    wire new_Jinkela_wire_409;
    wire new_Jinkela_wire_603;
    wire new_Jinkela_wire_219;
    wire new_Jinkela_wire_372;
    wire new_Jinkela_wire_448;
    wire new_Jinkela_wire_861;
    wire new_Jinkela_wire_599;
    wire new_Jinkela_wire_710;
    wire new_Jinkela_wire_482;
    wire new_Jinkela_wire_347;
    wire new_Jinkela_wire_761;
    wire new_Jinkela_wire_806;
    wire new_Jinkela_wire_946;
    wire new_Jinkela_wire_768;
    wire new_Jinkela_wire_660;
    wire new_Jinkela_wire_734;
    wire new_Jinkela_wire_308;
    wire new_Jinkela_wire_123;
    wire new_Jinkela_wire_207;
    wire _065_;
    wire new_Jinkela_wire_793;
    wire new_Jinkela_wire_135;
    wire new_Jinkela_wire_264;
    wire new_Jinkela_wire_282;
    wire new_Jinkela_wire_908;
    wire new_Jinkela_wire_48;
    wire new_Jinkela_wire_351;
    wire _009_;
    wire new_Jinkela_wire_128;
    wire new_Jinkela_wire_151;
    wire new_Jinkela_wire_198;
    wire new_Jinkela_wire_109;
    wire new_Jinkela_wire_758;
    wire new_Jinkela_wire_900;
    wire new_Jinkela_wire_978;
    wire new_Jinkela_wire_344;
    wire new_Jinkela_wire_950;
    wire new_Jinkela_wire_314;
    wire new_Jinkela_wire_553;
    wire _098_;
    wire new_Jinkela_wire_310;
    wire new_Jinkela_wire_810;
    wire new_Jinkela_wire_622;
    wire new_Jinkela_wire_542;
    wire new_Jinkela_wire_146;
    wire new_Jinkela_wire_430;
    wire _108_;
    wire new_Jinkela_wire_609;
    wire new_Jinkela_wire_538;
    wire new_Jinkela_wire_769;
    wire new_Jinkela_wire_11;
    wire new_Jinkela_wire_800;
    wire new_Jinkela_wire_114;
    wire new_Jinkela_wire_581;
    wire new_Jinkela_wire_498;
    wire new_Jinkela_wire_601;
    wire new_Jinkela_wire_472;
    wire new_Jinkela_wire_266;
    wire new_Jinkela_wire_414;
    wire new_Jinkela_wire_631;
    wire new_Jinkela_wire_284;
    wire _109_;
    wire new_Jinkela_wire_797;
    wire new_Jinkela_wire_238;
    wire new_Jinkela_wire_194;
    wire new_Jinkela_wire_577;
    wire new_Jinkela_wire_646;
    wire new_Jinkela_wire_478;
    wire new_Jinkela_wire_575;
    wire new_Jinkela_wire_720;
    wire new_Jinkela_wire_773;
    wire new_Jinkela_wire_272;
    wire new_Jinkela_wire_795;
    wire new_Jinkela_wire_293;
    wire _110_;
    wire new_Jinkela_wire_939;
    wire new_Jinkela_wire_801;
    wire new_Jinkela_wire_992;
    wire new_Jinkela_wire_339;
    wire new_Jinkela_wire_947;
    wire new_Jinkela_wire_51;
    wire new_Jinkela_wire_639;
    wire new_Jinkela_wire_0;
    wire new_Jinkela_wire_305;
    wire _079_;
    wire new_Jinkela_wire_691;
    wire new_Jinkela_wire_187;
    wire new_Jinkela_wire_216;
    wire new_Jinkela_wire_759;
    wire new_Jinkela_wire_635;
    wire new_Jinkela_wire_84;
    wire new_Jinkela_wire_246;
    wire new_Jinkela_wire_721;
    wire new_Jinkela_wire_781;
    wire new_Jinkela_wire_191;
    wire new_Jinkela_wire_895;
    wire new_Jinkela_wire_866;
    wire _007_;
    wire _090_;
    wire _010_;
    wire new_Jinkela_wire_10;
    wire new_Jinkela_wire_857;
    wire new_Jinkela_wire_253;
    wire new_Jinkela_wire_894;
    wire new_Jinkela_wire_406;
    wire new_Jinkela_wire_949;
    wire new_Jinkela_wire_237;
    wire new_Jinkela_wire_626;
    wire new_Jinkela_wire_302;
    wire _001_;
    wire new_Jinkela_wire_874;
    wire new_Jinkela_wire_505;
    wire new_Jinkela_wire_213;
    wire new_Jinkela_wire_445;
    wire new_Jinkela_wire_530;
    wire new_Jinkela_wire_819;
    wire _040_;
    wire new_Jinkela_wire_292;
    wire new_Jinkela_wire_392;
    wire new_Jinkela_wire_864;
    input N86;
    input N69;
    input N34;
    input N92;
    input N27;
    input N43;
    input N47;
    input N79;
    input N73;
    input N24;
    input N108;
    input N1;
    input N82;
    input N56;
    input N102;
    input N17;
    input N50;
    input N63;
    input N76;
    input N99;
    input N8;
    input N11;
    input N21;
    input N30;
    input N66;
    input N89;
    input N40;
    input N53;
    input N115;
    input N14;
    input N105;
    input N60;
    input N4;
    input N95;
    input N37;
    input N112;
    output N430;
    output N431;
    output N223;
    output N432;
    output N329;
    output N421;
    output N370;

    bfr new_Jinkela_buffer_683 (
        .din(_016_),
        .dout(new_Jinkela_wire_801)
    );

    spl2 new_Jinkela_splitter_22 (
        .a(N89),
        .b(new_Jinkela_wire_382),
        .c(new_Jinkela_wire_383)
    );

    bfr new_Jinkela_buffer_768 (
        .din(new_Jinkela_wire_905),
        .dout(new_Jinkela_wire_906)
    );

    bfr new_Jinkela_buffer_287 (
        .din(new_Jinkela_wire_326),
        .dout(new_Jinkela_wire_327)
    );

    bfr new_Jinkela_buffer_551 (
        .din(new_Jinkela_wire_616),
        .dout(new_Jinkela_wire_617)
    );

    bfr new_Jinkela_buffer_674 (
        .din(new_Jinkela_wire_791),
        .dout(new_Jinkela_wire_792)
    );

    spl4L new_Jinkela_splitter_52 (
        .a(new_Jinkela_wire_784),
        .b(new_Jinkela_wire_785),
        .d(new_Jinkela_wire_786),
        .e(new_Jinkela_wire_787),
        .c(new_Jinkela_wire_788)
    );

    bfr new_Jinkela_buffer_276 (
        .din(new_Jinkela_wire_313),
        .dout(new_Jinkela_wire_314)
    );

    bfr new_Jinkela_buffer_586 (
        .din(new_Jinkela_wire_668),
        .dout(new_Jinkela_wire_669)
    );

    bfr new_Jinkela_buffer_560 (
        .din(new_Jinkela_wire_638),
        .dout(new_Jinkela_wire_639)
    );

    bfr new_Jinkela_buffer_293 (
        .din(new_Jinkela_wire_332),
        .dout(new_Jinkela_wire_333)
    );

    bfr new_Jinkela_buffer_552 (
        .din(new_Jinkela_wire_617),
        .dout(new_Jinkela_wire_618)
    );

    bfr new_Jinkela_buffer_681 (
        .din(_063_),
        .dout(new_Jinkela_wire_799)
    );

    bfr new_Jinkela_buffer_277 (
        .din(new_Jinkela_wire_314),
        .dout(new_Jinkela_wire_315)
    );

    bfr new_Jinkela_buffer_682 (
        .din(new_Jinkela_wire_799),
        .dout(new_Jinkela_wire_800)
    );

    bfr new_Jinkela_buffer_288 (
        .din(new_Jinkela_wire_327),
        .dout(new_Jinkela_wire_328)
    );

    spl2 new_Jinkela_splitter_40 (
        .a(_025_),
        .b(new_Jinkela_wire_683),
        .c(new_Jinkela_wire_684)
    );

    bfr new_Jinkela_buffer_561 (
        .din(new_Jinkela_wire_639),
        .dout(new_Jinkela_wire_640)
    );

    spl2 new_Jinkela_splitter_54 (
        .a(_008_),
        .b(new_Jinkela_wire_802),
        .c(new_Jinkela_wire_803)
    );

    bfr new_Jinkela_buffer_278 (
        .din(new_Jinkela_wire_315),
        .dout(new_Jinkela_wire_316)
    );

    bfr new_Jinkela_buffer_675 (
        .din(new_Jinkela_wire_792),
        .dout(new_Jinkela_wire_793)
    );

    bfr new_Jinkela_buffer_593 (
        .din(new_Jinkela_wire_677),
        .dout(new_Jinkela_wire_678)
    );

    bfr new_Jinkela_buffer_346 (
        .din(N40),
        .dout(new_Jinkela_wire_392)
    );

    bfr new_Jinkela_buffer_672 (
        .din(_068_),
        .dout(new_Jinkela_wire_775)
    );

    spl2 new_Jinkela_splitter_55 (
        .a(_035_),
        .b(new_Jinkela_wire_813),
        .c(new_Jinkela_wire_814)
    );

    bfr new_Jinkela_buffer_317 (
        .din(new_Jinkela_wire_360),
        .dout(new_Jinkela_wire_361)
    );

    bfr new_Jinkela_buffer_562 (
        .din(new_Jinkela_wire_640),
        .dout(new_Jinkela_wire_641)
    );

    bfr new_Jinkela_buffer_684 (
        .din(new_Jinkela_wire_803),
        .dout(new_Jinkela_wire_804)
    );

    bfr new_Jinkela_buffer_279 (
        .din(new_Jinkela_wire_316),
        .dout(new_Jinkela_wire_317)
    );

    bfr new_Jinkela_buffer_676 (
        .din(new_Jinkela_wire_793),
        .dout(new_Jinkela_wire_794)
    );

    bfr new_Jinkela_buffer_289 (
        .din(new_Jinkela_wire_328),
        .dout(new_Jinkela_wire_329)
    );

    bfr new_Jinkela_buffer_587 (
        .din(new_Jinkela_wire_669),
        .dout(new_Jinkela_wire_670)
    );

    bfr new_Jinkela_buffer_563 (
        .din(new_Jinkela_wire_641),
        .dout(new_Jinkela_wire_642)
    );

    bfr new_Jinkela_buffer_280 (
        .din(new_Jinkela_wire_317),
        .dout(new_Jinkela_wire_318)
    );

    bfr new_Jinkela_buffer_677 (
        .din(new_Jinkela_wire_794),
        .dout(new_Jinkela_wire_795)
    );

    bfr new_Jinkela_buffer_764 (
        .din(new_Jinkela_wire_897),
        .dout(new_Jinkela_wire_898)
    );

    bfr new_Jinkela_buffer_294 (
        .din(new_Jinkela_wire_333),
        .dout(new_Jinkela_wire_334)
    );

    bfr new_Jinkela_buffer_564 (
        .din(new_Jinkela_wire_642),
        .dout(new_Jinkela_wire_643)
    );

    spl2 new_Jinkela_splitter_56 (
        .a(_042_),
        .b(new_Jinkela_wire_816),
        .c(new_Jinkela_wire_817)
    );

    bfr new_Jinkela_buffer_281 (
        .din(new_Jinkela_wire_318),
        .dout(new_Jinkela_wire_319)
    );

    bfr new_Jinkela_buffer_678 (
        .din(new_Jinkela_wire_795),
        .dout(new_Jinkela_wire_796)
    );

    spl2 new_Jinkela_splitter_41 (
        .a(_022_),
        .b(new_Jinkela_wire_694),
        .c(new_Jinkela_wire_695)
    );

    bfr new_Jinkela_buffer_309 (
        .din(new_Jinkela_wire_352),
        .dout(new_Jinkela_wire_353)
    );

    bfr new_Jinkela_buffer_588 (
        .din(new_Jinkela_wire_670),
        .dout(new_Jinkela_wire_671)
    );

    bfr new_Jinkela_buffer_755 (
        .din(new_Jinkela_wire_886),
        .dout(new_Jinkela_wire_887)
    );

    bfr new_Jinkela_buffer_565 (
        .din(new_Jinkela_wire_643),
        .dout(new_Jinkela_wire_644)
    );

    bfr new_Jinkela_buffer_295 (
        .din(new_Jinkela_wire_334),
        .dout(new_Jinkela_wire_335)
    );

    bfr new_Jinkela_buffer_679 (
        .din(new_Jinkela_wire_796),
        .dout(new_Jinkela_wire_797)
    );

    bfr new_Jinkela_buffer_685 (
        .din(new_Jinkela_wire_804),
        .dout(new_Jinkela_wire_805)
    );

    bfr new_Jinkela_buffer_338 (
        .din(new_Jinkela_wire_383),
        .dout(new_Jinkela_wire_384)
    );

    bfr new_Jinkela_buffer_566 (
        .din(new_Jinkela_wire_644),
        .dout(new_Jinkela_wire_645)
    );

    bfr new_Jinkela_buffer_296 (
        .din(new_Jinkela_wire_335),
        .dout(new_Jinkela_wire_336)
    );

    bfr new_Jinkela_buffer_680 (
        .din(new_Jinkela_wire_797),
        .dout(new_Jinkela_wire_798)
    );

    bfr new_Jinkela_buffer_310 (
        .din(new_Jinkela_wire_353),
        .dout(new_Jinkela_wire_354)
    );

    bfr new_Jinkela_buffer_589 (
        .din(new_Jinkela_wire_671),
        .dout(new_Jinkela_wire_672)
    );

    bfr new_Jinkela_buffer_693 (
        .din(new_Jinkela_wire_814),
        .dout(new_Jinkela_wire_815)
    );

    bfr new_Jinkela_buffer_567 (
        .din(new_Jinkela_wire_645),
        .dout(new_Jinkela_wire_646)
    );

    bfr new_Jinkela_buffer_694 (
        .din(_062_),
        .dout(new_Jinkela_wire_818)
    );

    bfr new_Jinkela_buffer_297 (
        .din(new_Jinkela_wire_336),
        .dout(new_Jinkela_wire_337)
    );

    bfr new_Jinkela_buffer_686 (
        .din(new_Jinkela_wire_805),
        .dout(new_Jinkela_wire_806)
    );

    bfr new_Jinkela_buffer_594 (
        .din(new_Jinkela_wire_678),
        .dout(new_Jinkela_wire_679)
    );

    spl2 new_Jinkela_splitter_57 (
        .a(_003_),
        .b(new_Jinkela_wire_827),
        .c(new_Jinkela_wire_828)
    );

    bfr new_Jinkela_buffer_318 (
        .din(new_Jinkela_wire_361),
        .dout(new_Jinkela_wire_362)
    );

    bfr new_Jinkela_buffer_568 (
        .din(new_Jinkela_wire_646),
        .dout(new_Jinkela_wire_647)
    );

    bfr new_Jinkela_buffer_298 (
        .din(new_Jinkela_wire_337),
        .dout(new_Jinkela_wire_338)
    );

    bfr new_Jinkela_buffer_687 (
        .din(new_Jinkela_wire_806),
        .dout(new_Jinkela_wire_807)
    );

    bfr new_Jinkela_buffer_311 (
        .din(new_Jinkela_wire_354),
        .dout(new_Jinkela_wire_355)
    );

    bfr new_Jinkela_buffer_590 (
        .din(new_Jinkela_wire_672),
        .dout(new_Jinkela_wire_673)
    );

    bfr new_Jinkela_buffer_569 (
        .din(new_Jinkela_wire_647),
        .dout(new_Jinkela_wire_648)
    );

    bfr new_Jinkela_buffer_695 (
        .din(new_net_198),
        .dout(new_Jinkela_wire_819)
    );

    bfr new_Jinkela_buffer_299 (
        .din(new_Jinkela_wire_338),
        .dout(new_Jinkela_wire_339)
    );

    bfr new_Jinkela_buffer_688 (
        .din(new_Jinkela_wire_807),
        .dout(new_Jinkela_wire_808)
    );

    bfr new_Jinkela_buffer_598 (
        .din(new_Jinkela_wire_684),
        .dout(new_Jinkela_wire_685)
    );

    bfr new_Jinkela_buffer_712 (
        .din(_054_),
        .dout(new_Jinkela_wire_838)
    );

    bfr new_Jinkela_buffer_570 (
        .din(new_Jinkela_wire_648),
        .dout(new_Jinkela_wire_649)
    );

    bfr new_Jinkela_buffer_696 (
        .din(new_Jinkela_wire_819),
        .dout(new_Jinkela_wire_820)
    );

    bfr new_Jinkela_buffer_300 (
        .din(new_Jinkela_wire_339),
        .dout(new_Jinkela_wire_340)
    );

    bfr new_Jinkela_buffer_689 (
        .din(new_Jinkela_wire_808),
        .dout(new_Jinkela_wire_809)
    );

    spl2 new_Jinkela_splitter_42 (
        .a(_104_),
        .b(new_Jinkela_wire_705),
        .c(new_Jinkela_wire_706)
    );

    bfr new_Jinkela_buffer_312 (
        .din(new_Jinkela_wire_355),
        .dout(new_Jinkela_wire_356)
    );

    bfr new_Jinkela_buffer_591 (
        .din(new_Jinkela_wire_673),
        .dout(new_Jinkela_wire_674)
    );

    bfr new_Jinkela_buffer_571 (
        .din(new_Jinkela_wire_649),
        .dout(new_Jinkela_wire_650)
    );

    bfr new_Jinkela_buffer_703 (
        .din(new_Jinkela_wire_828),
        .dout(new_Jinkela_wire_829)
    );

    spl2 new_Jinkela_splitter_20 (
        .a(new_Jinkela_wire_340),
        .b(new_Jinkela_wire_341),
        .c(new_Jinkela_wire_342)
    );

    bfr new_Jinkela_buffer_690 (
        .din(new_Jinkela_wire_809),
        .dout(new_Jinkela_wire_810)
    );

    bfr new_Jinkela_buffer_301 (
        .din(new_Jinkela_wire_342),
        .dout(new_Jinkela_wire_343)
    );

    bfr new_Jinkela_buffer_595 (
        .din(new_Jinkela_wire_679),
        .dout(new_Jinkela_wire_680)
    );

    bfr new_Jinkela_buffer_572 (
        .din(new_Jinkela_wire_650),
        .dout(new_Jinkela_wire_651)
    );

    bfr new_Jinkela_buffer_697 (
        .din(new_Jinkela_wire_820),
        .dout(new_Jinkela_wire_821)
    );

    bfr new_Jinkela_buffer_691 (
        .din(new_Jinkela_wire_810),
        .dout(new_Jinkela_wire_811)
    );

    spl2 new_Jinkela_splitter_65 (
        .a(_094_),
        .b(new_Jinkela_wire_918),
        .c(new_Jinkela_wire_919)
    );

    bfr new_Jinkela_buffer_319 (
        .din(new_Jinkela_wire_362),
        .dout(new_Jinkela_wire_363)
    );

    bfr new_Jinkela_buffer_313 (
        .din(new_Jinkela_wire_356),
        .dout(new_Jinkela_wire_357)
    );

    bfr new_Jinkela_buffer_592 (
        .din(new_Jinkela_wire_674),
        .dout(new_Jinkela_wire_675)
    );

    bfr new_Jinkela_buffer_573 (
        .din(new_Jinkela_wire_651),
        .dout(new_Jinkela_wire_652)
    );

    bfr new_Jinkela_buffer_302 (
        .din(new_Jinkela_wire_343),
        .dout(new_Jinkela_wire_344)
    );

    bfr new_Jinkela_buffer_692 (
        .din(new_Jinkela_wire_811),
        .dout(new_Jinkela_wire_812)
    );

    spl2 new_Jinkela_splitter_66 (
        .a(_107_),
        .b(new_Jinkela_wire_928),
        .c(new_Jinkela_wire_929)
    );

    bfr new_Jinkela_buffer_375 (
        .din(N53),
        .dout(new_Jinkela_wire_423)
    );

    bfr new_Jinkela_buffer_574 (
        .din(new_Jinkela_wire_652),
        .dout(new_Jinkela_wire_653)
    );

    bfr new_Jinkela_buffer_698 (
        .din(new_Jinkela_wire_821),
        .dout(new_Jinkela_wire_822)
    );

    bfr new_Jinkela_buffer_303 (
        .din(new_Jinkela_wire_344),
        .dout(new_Jinkela_wire_345)
    );

    bfr new_Jinkela_buffer_624 (
        .din(_049_),
        .dout(new_Jinkela_wire_715)
    );

    spl2 new_Jinkela_splitter_58 (
        .a(_045_),
        .b(new_Jinkela_wire_844),
        .c(new_Jinkela_wire_845)
    );

    bfr new_Jinkela_buffer_314 (
        .din(new_Jinkela_wire_357),
        .dout(new_Jinkela_wire_358)
    );

    bfr new_Jinkela_buffer_596 (
        .din(new_Jinkela_wire_680),
        .dout(new_Jinkela_wire_681)
    );

    spl2 new_Jinkela_splitter_59 (
        .a(_011_),
        .b(new_Jinkela_wire_846),
        .c(new_Jinkela_wire_847)
    );

    bfr new_Jinkela_buffer_575 (
        .din(new_Jinkela_wire_653),
        .dout(new_Jinkela_wire_654)
    );

    bfr new_Jinkela_buffer_699 (
        .din(new_Jinkela_wire_822),
        .dout(new_Jinkela_wire_823)
    );

    bfr new_Jinkela_buffer_778 (
        .din(new_Jinkela_wire_919),
        .dout(new_Jinkela_wire_920)
    );

    bfr new_Jinkela_buffer_304 (
        .din(new_Jinkela_wire_345),
        .dout(new_Jinkela_wire_346)
    );

    bfr new_Jinkela_buffer_713 (
        .din(new_Jinkela_wire_838),
        .dout(new_Jinkela_wire_839)
    );

    bfr new_Jinkela_buffer_599 (
        .din(new_Jinkela_wire_685),
        .dout(new_Jinkela_wire_686)
    );

    bfr new_Jinkela_buffer_704 (
        .din(new_Jinkela_wire_829),
        .dout(new_Jinkela_wire_830)
    );

    bfr new_Jinkela_buffer_320 (
        .din(new_Jinkela_wire_363),
        .dout(new_Jinkela_wire_364)
    );

    bfr new_Jinkela_buffer_576 (
        .din(new_Jinkela_wire_654),
        .dout(new_Jinkela_wire_655)
    );

    bfr new_Jinkela_buffer_700 (
        .din(new_Jinkela_wire_823),
        .dout(new_Jinkela_wire_824)
    );

    bfr new_Jinkela_buffer_305 (
        .din(new_Jinkela_wire_346),
        .dout(new_Jinkela_wire_347)
    );

    bfr new_Jinkela_buffer_770 (
        .din(new_Jinkela_wire_909),
        .dout(new_Jinkela_wire_910)
    );

    bfr new_Jinkela_buffer_315 (
        .din(new_Jinkela_wire_358),
        .dout(new_Jinkela_wire_359)
    );

    bfr new_Jinkela_buffer_597 (
        .din(new_Jinkela_wire_681),
        .dout(new_Jinkela_wire_682)
    );

    bfr new_Jinkela_buffer_577 (
        .din(new_Jinkela_wire_655),
        .dout(new_Jinkela_wire_656)
    );

    bfr new_Jinkela_buffer_701 (
        .din(new_Jinkela_wire_824),
        .dout(new_Jinkela_wire_825)
    );

    bfr new_Jinkela_buffer_306 (
        .din(new_Jinkela_wire_347),
        .dout(new_Jinkela_wire_348)
    );

    spl2 new_Jinkela_splitter_60 (
        .a(_097_),
        .b(new_Jinkela_wire_857),
        .c(new_Jinkela_wire_858)
    );

    bfr new_Jinkela_buffer_607 (
        .din(new_Jinkela_wire_695),
        .dout(new_Jinkela_wire_696)
    );

    bfr new_Jinkela_buffer_705 (
        .din(new_Jinkela_wire_830),
        .dout(new_Jinkela_wire_831)
    );

    bfr new_Jinkela_buffer_404 (
        .din(N115),
        .dout(new_Jinkela_wire_454)
    );

    bfr new_Jinkela_buffer_578 (
        .din(new_Jinkela_wire_656),
        .dout(new_Jinkela_wire_657)
    );

    bfr new_Jinkela_buffer_702 (
        .din(new_Jinkela_wire_825),
        .dout(new_Jinkela_wire_826)
    );

    bfr new_Jinkela_buffer_307 (
        .din(new_Jinkela_wire_348),
        .dout(new_Jinkela_wire_349)
    );

    bfr new_Jinkela_buffer_339 (
        .din(new_Jinkela_wire_384),
        .dout(new_Jinkela_wire_385)
    );

    bfr new_Jinkela_buffer_600 (
        .din(new_Jinkela_wire_686),
        .dout(new_Jinkela_wire_687)
    );

    bfr new_Jinkela_buffer_321 (
        .din(new_Jinkela_wire_364),
        .dout(new_Jinkela_wire_365)
    );

    bfr new_Jinkela_buffer_579 (
        .din(new_Jinkela_wire_657),
        .dout(new_Jinkela_wire_658)
    );

    bfr new_Jinkela_buffer_714 (
        .din(new_Jinkela_wire_839),
        .dout(new_Jinkela_wire_840)
    );

    bfr new_Jinkela_buffer_85 (
        .din(new_Jinkela_wire_92),
        .dout(new_Jinkela_wire_93)
    );

    bfr new_Jinkela_buffer_134 (
        .din(new_Jinkela_wire_147),
        .dout(new_Jinkela_wire_148)
    );

    bfr new_Jinkela_buffer_412 (
        .din(new_Jinkela_wire_461),
        .dout(new_Jinkela_wire_462)
    );

    and_bi _230_ (
        .a(_053_),
        .b(new_Jinkela_wire_812),
        .c(_054_)
    );

    bfr new_Jinkela_buffer_787 (
        .din(new_Jinkela_wire_930),
        .dout(new_Jinkela_wire_931)
    );

    bfr new_Jinkela_buffer_68 (
        .din(new_Jinkela_wire_75),
        .dout(new_Jinkela_wire_76)
    );

    spl2 new_Jinkela_splitter_6 (
        .a(new_Jinkela_wire_133),
        .b(new_Jinkela_wire_134),
        .c(new_Jinkela_wire_135)
    );

    bfr new_Jinkela_buffer_392 (
        .din(new_Jinkela_wire_439),
        .dout(new_Jinkela_wire_440)
    );

    and_bi _231_ (
        .a(_052_),
        .b(new_Jinkela_wire_843),
        .c(N421)
    );

    bfr new_Jinkela_buffer_782 (
        .din(new_Jinkela_wire_923),
        .dout(new_Jinkela_wire_924)
    );

    bfr new_Jinkela_buffer_107 (
        .din(new_Jinkela_wire_118),
        .dout(new_Jinkela_wire_119)
    );

    bfr new_Jinkela_buffer_122 (
        .din(new_Jinkela_wire_135),
        .dout(new_Jinkela_wire_136)
    );

    bfr new_Jinkela_buffer_437 (
        .din(new_Jinkela_wire_488),
        .dout(new_Jinkela_wire_489)
    );

    and_bi _232_ (
        .a(new_Jinkela_wire_845),
        .b(new_Jinkela_wire_992),
        .c(_055_)
    );

    bfr new_Jinkela_buffer_802 (
        .din(new_Jinkela_wire_949),
        .dout(new_Jinkela_wire_950)
    );

    bfr new_Jinkela_buffer_806 (
        .din(_058_),
        .dout(new_Jinkela_wire_954)
    );

    bfr new_Jinkela_buffer_69 (
        .din(new_Jinkela_wire_76),
        .dout(new_Jinkela_wire_77)
    );

    bfr new_Jinkela_buffer_177 (
        .din(new_Jinkela_wire_196),
        .dout(new_Jinkela_wire_197)
    );

    bfr new_Jinkela_buffer_393 (
        .din(new_Jinkela_wire_440),
        .dout(new_Jinkela_wire_441)
    );

    or_bb _233_ (
        .a(_055_),
        .b(new_Jinkela_wire_815),
        .c(new_net_196)
    );

    bfr new_Jinkela_buffer_783 (
        .din(new_Jinkela_wire_924),
        .dout(new_Jinkela_wire_925)
    );

    bfr new_Jinkela_buffer_86 (
        .din(new_Jinkela_wire_93),
        .dout(new_Jinkela_wire_94)
    );

    bfr new_Jinkela_buffer_135 (
        .din(new_Jinkela_wire_148),
        .dout(new_Jinkela_wire_149)
    );

    bfr new_Jinkela_buffer_413 (
        .din(new_Jinkela_wire_462),
        .dout(new_Jinkela_wire_463)
    );

    or_bi _234_ (
        .a(new_Jinkela_wire_994),
        .b(new_Jinkela_wire_906),
        .c(_056_)
    );

    bfr new_Jinkela_buffer_788 (
        .din(new_Jinkela_wire_931),
        .dout(new_Jinkela_wire_932)
    );

    bfr new_Jinkela_buffer_70 (
        .din(new_Jinkela_wire_77),
        .dout(new_Jinkela_wire_78)
    );

    bfr new_Jinkela_buffer_123 (
        .din(new_Jinkela_wire_136),
        .dout(new_Jinkela_wire_137)
    );

    bfr new_Jinkela_buffer_394 (
        .din(new_Jinkela_wire_441),
        .dout(new_Jinkela_wire_442)
    );

    and_bi _235_ (
        .a(new_Jinkela_wire_817),
        .b(new_Jinkela_wire_662),
        .c(_057_)
    );

    bfr new_Jinkela_buffer_784 (
        .din(new_Jinkela_wire_925),
        .dout(new_Jinkela_wire_926)
    );

    bfr new_Jinkela_buffer_114 (
        .din(new_Jinkela_wire_125),
        .dout(new_Jinkela_wire_126)
    );

    bfr new_Jinkela_buffer_161 (
        .din(new_Jinkela_wire_176),
        .dout(new_Jinkela_wire_177)
    );

    bfr new_Jinkela_buffer_464 (
        .din(new_Jinkela_wire_517),
        .dout(new_Jinkela_wire_518)
    );

    or_bb _236_ (
        .a(_057_),
        .b(new_Jinkela_wire_901),
        .c(_058_)
    );

    bfr new_Jinkela_buffer_71 (
        .din(new_Jinkela_wire_78),
        .dout(new_Jinkela_wire_79)
    );

    bfr new_Jinkela_buffer_124 (
        .din(new_Jinkela_wire_137),
        .dout(new_Jinkela_wire_138)
    );

    bfr new_Jinkela_buffer_395 (
        .din(new_Jinkela_wire_442),
        .dout(new_Jinkela_wire_443)
    );

    and_bi _237_ (
        .a(_056_),
        .b(new_Jinkela_wire_954),
        .c(_059_)
    );

    bfr new_Jinkela_buffer_785 (
        .din(new_Jinkela_wire_926),
        .dout(new_Jinkela_wire_927)
    );

    bfr new_Jinkela_buffer_87 (
        .din(new_Jinkela_wire_94),
        .dout(new_Jinkela_wire_95)
    );

    bfr new_Jinkela_buffer_136 (
        .din(new_Jinkela_wire_149),
        .dout(new_Jinkela_wire_150)
    );

    bfr new_Jinkela_buffer_414 (
        .din(new_Jinkela_wire_463),
        .dout(new_Jinkela_wire_464)
    );

    and_bi _238_ (
        .a(new_Jinkela_wire_953),
        .b(_059_),
        .c(_060_)
    );

    bfr new_Jinkela_buffer_789 (
        .din(new_Jinkela_wire_932),
        .dout(new_Jinkela_wire_933)
    );

    bfr new_Jinkela_buffer_72 (
        .din(new_Jinkela_wire_79),
        .dout(new_Jinkela_wire_80)
    );

    bfr new_Jinkela_buffer_125 (
        .din(new_Jinkela_wire_138),
        .dout(new_Jinkela_wire_139)
    );

    spl2 new_Jinkela_splitter_24 (
        .a(new_Jinkela_wire_443),
        .b(new_Jinkela_wire_444),
        .c(new_Jinkela_wire_445)
    );

    or_bb _239_ (
        .a(_060_),
        .b(new_Jinkela_wire_682),
        .c(N432)
    );

    bfr new_Jinkela_buffer_795 (
        .din(new_Jinkela_wire_940),
        .dout(new_Jinkela_wire_941)
    );

    bfr new_Jinkela_buffer_108 (
        .din(new_Jinkela_wire_119),
        .dout(new_Jinkela_wire_120)
    );

    bfr new_Jinkela_buffer_396 (
        .din(new_Jinkela_wire_445),
        .dout(new_Jinkela_wire_446)
    );

    bfr new_Jinkela_buffer_790 (
        .din(new_Jinkela_wire_933),
        .dout(new_Jinkela_wire_934)
    );

    inv _240_ (
        .din(new_Jinkela_wire_631),
        .dout(new_net_194)
    );

    spl2 new_Jinkela_splitter_11 (
        .a(N82),
        .b(new_Jinkela_wire_216),
        .c(new_Jinkela_wire_217)
    );

    spl2 new_Jinkela_splitter_67 (
        .a(_101_),
        .b(new_Jinkela_wire_938),
        .c(new_Jinkela_wire_939)
    );

    bfr new_Jinkela_buffer_88 (
        .din(new_Jinkela_wire_95),
        .dout(new_Jinkela_wire_96)
    );

    bfr new_Jinkela_buffer_126 (
        .din(new_Jinkela_wire_139),
        .dout(new_Jinkela_wire_140)
    );

    bfr new_Jinkela_buffer_438 (
        .din(new_Jinkela_wire_489),
        .dout(new_Jinkela_wire_490)
    );

    spl2 new_Jinkela_splitter_69 (
        .a(_000_),
        .b(new_Jinkela_wire_955),
        .c(new_Jinkela_wire_956)
    );

    bfr new_Jinkela_buffer_137 (
        .din(new_Jinkela_wire_150),
        .dout(new_Jinkela_wire_151)
    );

    bfr new_Jinkela_buffer_415 (
        .din(new_Jinkela_wire_464),
        .dout(new_Jinkela_wire_465)
    );

    bfr new_Jinkela_buffer_791 (
        .din(new_Jinkela_wire_934),
        .dout(new_Jinkela_wire_935)
    );

    spl2 new_Jinkela_splitter_9 (
        .a(N108),
        .b(new_Jinkela_wire_195),
        .c(new_Jinkela_wire_196)
    );

    bfr new_Jinkela_buffer_89 (
        .din(new_Jinkela_wire_96),
        .dout(new_Jinkela_wire_97)
    );

    bfr new_Jinkela_buffer_127 (
        .din(new_Jinkela_wire_140),
        .dout(new_Jinkela_wire_141)
    );

    bfr new_Jinkela_buffer_397 (
        .din(new_Jinkela_wire_446),
        .dout(new_Jinkela_wire_447)
    );

    bfr new_Jinkela_buffer_772 (
        .din(new_Jinkela_wire_911),
        .dout(new_Jinkela_wire_912)
    );

    bfr new_Jinkela_buffer_796 (
        .din(new_Jinkela_wire_941),
        .dout(new_Jinkela_wire_942)
    );

    bfr new_Jinkela_buffer_109 (
        .din(new_Jinkela_wire_120),
        .dout(new_Jinkela_wire_121)
    );

    bfr new_Jinkela_buffer_162 (
        .din(new_Jinkela_wire_177),
        .dout(new_Jinkela_wire_178)
    );

    bfr new_Jinkela_buffer_492 (
        .din(new_Jinkela_wire_547),
        .dout(new_Jinkela_wire_548)
    );

    bfr new_Jinkela_buffer_792 (
        .din(new_Jinkela_wire_935),
        .dout(new_Jinkela_wire_936)
    );

    bfr new_Jinkela_buffer_90 (
        .din(new_Jinkela_wire_97),
        .dout(new_Jinkela_wire_98)
    );

    bfr new_Jinkela_buffer_128 (
        .din(new_Jinkela_wire_141),
        .dout(new_Jinkela_wire_142)
    );

    bfr new_Jinkela_buffer_398 (
        .din(new_Jinkela_wire_447),
        .dout(new_Jinkela_wire_448)
    );

    bfr new_Jinkela_buffer_807 (
        .din(new_Jinkela_wire_956),
        .dout(new_Jinkela_wire_957)
    );

    bfr new_Jinkela_buffer_816 (
        .din(_006_),
        .dout(new_Jinkela_wire_966)
    );

    bfr new_Jinkela_buffer_115 (
        .din(new_Jinkela_wire_126),
        .dout(new_Jinkela_wire_127)
    );

    bfr new_Jinkela_buffer_138 (
        .din(new_Jinkela_wire_151),
        .dout(new_Jinkela_wire_152)
    );

    bfr new_Jinkela_buffer_416 (
        .din(new_Jinkela_wire_465),
        .dout(new_Jinkela_wire_466)
    );

    bfr new_Jinkela_buffer_793 (
        .din(new_Jinkela_wire_936),
        .dout(new_Jinkela_wire_937)
    );

    bfr new_Jinkela_buffer_91 (
        .din(new_Jinkela_wire_98),
        .dout(new_Jinkela_wire_99)
    );

    bfr new_Jinkela_buffer_399 (
        .din(new_Jinkela_wire_448),
        .dout(new_Jinkela_wire_449)
    );

    bfr new_Jinkela_buffer_797 (
        .din(new_Jinkela_wire_942),
        .dout(new_Jinkela_wire_943)
    );

    bfr new_Jinkela_buffer_110 (
        .din(new_Jinkela_wire_121),
        .dout(new_Jinkela_wire_122)
    );

    bfr new_Jinkela_buffer_139 (
        .din(new_Jinkela_wire_152),
        .dout(new_Jinkela_wire_153)
    );

    bfr new_Jinkela_buffer_439 (
        .din(new_Jinkela_wire_490),
        .dout(new_Jinkela_wire_491)
    );

    bfr new_Jinkela_buffer_803 (
        .din(new_Jinkela_wire_950),
        .dout(new_Jinkela_wire_951)
    );

    bfr new_Jinkela_buffer_92 (
        .din(new_Jinkela_wire_99),
        .dout(new_Jinkela_wire_100)
    );

    bfr new_Jinkela_buffer_163 (
        .din(new_Jinkela_wire_178),
        .dout(new_Jinkela_wire_179)
    );

    bfr new_Jinkela_buffer_400 (
        .din(new_Jinkela_wire_449),
        .dout(new_Jinkela_wire_450)
    );

    bfr new_Jinkela_buffer_798 (
        .din(new_Jinkela_wire_943),
        .dout(new_Jinkela_wire_944)
    );

    bfr new_Jinkela_buffer_140 (
        .din(new_Jinkela_wire_153),
        .dout(new_Jinkela_wire_154)
    );

    bfr new_Jinkela_buffer_131 (
        .din(new_Jinkela_wire_144),
        .dout(new_Jinkela_wire_145)
    );

    bfr new_Jinkela_buffer_417 (
        .din(new_Jinkela_wire_466),
        .dout(new_Jinkela_wire_467)
    );

    bfr new_Jinkela_buffer_93 (
        .din(new_Jinkela_wire_100),
        .dout(new_Jinkela_wire_101)
    );

    bfr new_Jinkela_buffer_178 (
        .din(new_Jinkela_wire_197),
        .dout(new_Jinkela_wire_198)
    );

    bfr new_Jinkela_buffer_401 (
        .din(new_Jinkela_wire_450),
        .dout(new_Jinkela_wire_451)
    );

    bfr new_Jinkela_buffer_799 (
        .din(new_Jinkela_wire_944),
        .dout(new_Jinkela_wire_945)
    );

    bfr new_Jinkela_buffer_116 (
        .din(new_Jinkela_wire_127),
        .dout(new_Jinkela_wire_128)
    );

    bfr new_Jinkela_buffer_141 (
        .din(new_Jinkela_wire_154),
        .dout(new_Jinkela_wire_155)
    );

    bfr new_Jinkela_buffer_465 (
        .din(new_Jinkela_wire_518),
        .dout(new_Jinkela_wire_519)
    );

    bfr new_Jinkela_buffer_673 (
        .din(new_Jinkela_wire_790),
        .dout(new_Jinkela_wire_791)
    );

    bfr new_Jinkela_buffer_804 (
        .din(new_Jinkela_wire_951),
        .dout(new_Jinkela_wire_952)
    );

    spl2 new_Jinkela_splitter_4 (
        .a(new_Jinkela_wire_101),
        .b(new_Jinkela_wire_102),
        .c(new_Jinkela_wire_103)
    );

    bfr new_Jinkela_buffer_164 (
        .din(new_Jinkela_wire_179),
        .dout(new_Jinkela_wire_180)
    );

    bfr new_Jinkela_buffer_402 (
        .din(new_Jinkela_wire_451),
        .dout(new_Jinkela_wire_452)
    );

    bfr new_Jinkela_buffer_773 (
        .din(new_Jinkela_wire_912),
        .dout(new_Jinkela_wire_913)
    );

    bfr new_Jinkela_buffer_800 (
        .din(new_Jinkela_wire_945),
        .dout(new_Jinkela_wire_946)
    );

    bfr new_Jinkela_buffer_94 (
        .din(new_Jinkela_wire_103),
        .dout(new_Jinkela_wire_104)
    );

    bfr new_Jinkela_buffer_142 (
        .din(new_Jinkela_wire_155),
        .dout(new_Jinkela_wire_156)
    );

    bfr new_Jinkela_buffer_418 (
        .din(new_Jinkela_wire_467),
        .dout(new_Jinkela_wire_468)
    );

    bfr new_Jinkela_buffer_818 (
        .din(_039_),
        .dout(new_Jinkela_wire_968)
    );

    bfr new_Jinkela_buffer_159 (
        .din(new_Jinkela_wire_174),
        .dout(new_Jinkela_wire_175)
    );

    bfr new_Jinkela_buffer_186 (
        .din(new_Jinkela_wire_207),
        .dout(new_Jinkela_wire_208)
    );

    bfr new_Jinkela_buffer_403 (
        .din(new_Jinkela_wire_452),
        .dout(new_Jinkela_wire_453)
    );

    spl2 new_Jinkela_splitter_12 (
        .a(N56),
        .b(new_Jinkela_wire_227),
        .c(new_Jinkela_wire_228)
    );

    bfr new_Jinkela_buffer_801 (
        .din(new_Jinkela_wire_946),
        .dout(new_Jinkela_wire_947)
    );

    bfr new_Jinkela_buffer_117 (
        .din(new_Jinkela_wire_128),
        .dout(new_Jinkela_wire_129)
    );

    bfr new_Jinkela_buffer_143 (
        .din(new_Jinkela_wire_156),
        .dout(new_Jinkela_wire_157)
    );

    bfr new_Jinkela_buffer_440 (
        .din(new_Jinkela_wire_491),
        .dout(new_Jinkela_wire_492)
    );

    bfr new_Jinkela_buffer_805 (
        .din(new_Jinkela_wire_952),
        .dout(new_Jinkela_wire_953)
    );

    bfr new_Jinkela_buffer_95 (
        .din(new_Jinkela_wire_104),
        .dout(new_Jinkela_wire_105)
    );

    bfr new_Jinkela_buffer_165 (
        .din(new_Jinkela_wire_180),
        .dout(new_Jinkela_wire_181)
    );

    bfr new_Jinkela_buffer_419 (
        .din(new_Jinkela_wire_468),
        .dout(new_Jinkela_wire_469)
    );

    bfr new_Jinkela_buffer_817 (
        .din(new_Jinkela_wire_966),
        .dout(new_Jinkela_wire_967)
    );

    bfr new_Jinkela_buffer_144 (
        .din(new_Jinkela_wire_157),
        .dout(new_Jinkela_wire_158)
    );

    bfr new_Jinkela_buffer_132 (
        .din(new_Jinkela_wire_145),
        .dout(new_Jinkela_wire_146)
    );

    spl2 new_Jinkela_splitter_30 (
        .a(N95),
        .b(new_Jinkela_wire_578),
        .c(new_Jinkela_wire_579)
    );

    spl2 new_Jinkela_splitter_29 (
        .a(N4),
        .b(new_Jinkela_wire_567),
        .c(new_Jinkela_wire_568)
    );

    bfr new_Jinkela_buffer_779 (
        .din(new_Jinkela_wire_920),
        .dout(new_Jinkela_wire_921)
    );

    bfr new_Jinkela_buffer_808 (
        .din(new_Jinkela_wire_957),
        .dout(new_Jinkela_wire_958)
    );

    bfr new_Jinkela_buffer_96 (
        .din(new_Jinkela_wire_105),
        .dout(new_Jinkela_wire_106)
    );

    bfr new_Jinkela_buffer_179 (
        .din(new_Jinkela_wire_198),
        .dout(new_Jinkela_wire_199)
    );

    bfr new_Jinkela_buffer_420 (
        .din(new_Jinkela_wire_469),
        .dout(new_Jinkela_wire_470)
    );

    spl3L new_Jinkela_splitter_70 (
        .a(_077_),
        .b(new_Jinkela_wire_969),
        .d(new_Jinkela_wire_972),
        .c(new_Jinkela_wire_977)
    );

    bfr new_Jinkela_buffer_118 (
        .din(new_Jinkela_wire_129),
        .dout(new_Jinkela_wire_130)
    );

    bfr new_Jinkela_buffer_145 (
        .din(new_Jinkela_wire_158),
        .dout(new_Jinkela_wire_159)
    );

    bfr new_Jinkela_buffer_441 (
        .din(new_Jinkela_wire_492),
        .dout(new_Jinkela_wire_493)
    );

    bfr new_Jinkela_buffer_809 (
        .din(new_Jinkela_wire_958),
        .dout(new_Jinkela_wire_959)
    );

    bfr new_Jinkela_buffer_97 (
        .din(new_Jinkela_wire_106),
        .dout(new_Jinkela_wire_107)
    );

    bfr new_Jinkela_buffer_166 (
        .din(new_Jinkela_wire_181),
        .dout(new_Jinkela_wire_182)
    );

    bfr new_Jinkela_buffer_421 (
        .din(new_Jinkela_wire_470),
        .dout(new_Jinkela_wire_471)
    );

    spl3L new_Jinkela_splitter_75 (
        .a(_040_),
        .b(new_Jinkela_wire_992),
        .d(new_Jinkela_wire_993),
        .c(new_Jinkela_wire_994)
    );

    bfr new_Jinkela_buffer_146 (
        .din(new_Jinkela_wire_159),
        .dout(new_Jinkela_wire_160)
    );

    spl2 new_Jinkela_splitter_10 (
        .a(N1),
        .b(new_Jinkela_wire_206),
        .c(new_Jinkela_wire_207)
    );

    bfr new_Jinkela_buffer_466 (
        .din(new_Jinkela_wire_519),
        .dout(new_Jinkela_wire_520)
    );

    bfr new_Jinkela_buffer_810 (
        .din(new_Jinkela_wire_959),
        .dout(new_Jinkela_wire_960)
    );

    bfr new_Jinkela_buffer_98 (
        .din(new_Jinkela_wire_107),
        .dout(new_Jinkela_wire_108)
    );

    bfr new_Jinkela_buffer_422 (
        .din(new_Jinkela_wire_471),
        .dout(new_Jinkela_wire_472)
    );

    bfr new_Jinkela_buffer_194 (
        .din(new_Jinkela_wire_217),
        .dout(new_Jinkela_wire_218)
    );

    spl2 new_Jinkela_splitter_74 (
        .a(_079_),
        .b(new_Jinkela_wire_982),
        .c(new_Jinkela_wire_983)
    );

    bfr new_Jinkela_buffer_119 (
        .din(new_Jinkela_wire_130),
        .dout(new_Jinkela_wire_131)
    );

    bfr new_Jinkela_buffer_147 (
        .din(new_Jinkela_wire_160),
        .dout(new_Jinkela_wire_161)
    );

    bfr new_Jinkela_buffer_442 (
        .din(new_Jinkela_wire_493),
        .dout(new_Jinkela_wire_494)
    );

    bfr new_Jinkela_buffer_811 (
        .din(new_Jinkela_wire_960),
        .dout(new_Jinkela_wire_961)
    );

    bfr new_Jinkela_buffer_99 (
        .din(new_Jinkela_wire_108),
        .dout(new_Jinkela_wire_109)
    );

    bfr new_Jinkela_buffer_167 (
        .din(new_Jinkela_wire_182),
        .dout(new_Jinkela_wire_183)
    );

    bfr new_Jinkela_buffer_423 (
        .din(new_Jinkela_wire_472),
        .dout(new_Jinkela_wire_473)
    );

    bfr new_Jinkela_buffer_148 (
        .din(new_Jinkela_wire_161),
        .dout(new_Jinkela_wire_162)
    );

    bfr new_Jinkela_buffer_133 (
        .din(new_Jinkela_wire_146),
        .dout(new_Jinkela_wire_147)
    );

    bfr new_Jinkela_buffer_493 (
        .din(new_Jinkela_wire_548),
        .dout(new_Jinkela_wire_549)
    );

    bfr new_Jinkela_buffer_812 (
        .din(new_Jinkela_wire_961),
        .dout(new_Jinkela_wire_962)
    );

    bfr new_Jinkela_buffer_100 (
        .din(new_Jinkela_wire_109),
        .dout(new_Jinkela_wire_110)
    );

    bfr new_Jinkela_buffer_180 (
        .din(new_Jinkela_wire_199),
        .dout(new_Jinkela_wire_200)
    );

    bfr new_Jinkela_buffer_424 (
        .din(new_Jinkela_wire_473),
        .dout(new_Jinkela_wire_474)
    );

    bfr new_Jinkela_buffer_668 (
        .din(new_Jinkela_wire_768),
        .dout(new_Jinkela_wire_769)
    );

    spl2 new_Jinkela_splitter_71 (
        .a(new_Jinkela_wire_969),
        .b(new_Jinkela_wire_970),
        .c(new_Jinkela_wire_971)
    );

    bfr new_Jinkela_buffer_819 (
        .din(new_Jinkela_wire_983),
        .dout(new_Jinkela_wire_984)
    );

    bfr new_Jinkela_buffer_120 (
        .din(new_Jinkela_wire_131),
        .dout(new_Jinkela_wire_132)
    );

    bfr new_Jinkela_buffer_149 (
        .din(new_Jinkela_wire_162),
        .dout(new_Jinkela_wire_163)
    );

    bfr new_Jinkela_buffer_443 (
        .din(new_Jinkela_wire_494),
        .dout(new_Jinkela_wire_495)
    );

    bfr new_Jinkela_buffer_786 (
        .din(new_Jinkela_wire_929),
        .dout(new_Jinkela_wire_930)
    );

    bfr new_Jinkela_buffer_813 (
        .din(new_Jinkela_wire_962),
        .dout(new_Jinkela_wire_963)
    );

    bfr new_Jinkela_buffer_101 (
        .din(new_Jinkela_wire_110),
        .dout(new_Jinkela_wire_111)
    );

    bfr new_Jinkela_buffer_168 (
        .din(new_Jinkela_wire_183),
        .dout(new_Jinkela_wire_184)
    );

    spl2 new_Jinkela_splitter_25 (
        .a(new_Jinkela_wire_474),
        .b(new_Jinkela_wire_475),
        .c(new_Jinkela_wire_476)
    );

    spl4L new_Jinkela_splitter_72 (
        .a(new_Jinkela_wire_972),
        .b(new_Jinkela_wire_973),
        .d(new_Jinkela_wire_974),
        .e(new_Jinkela_wire_975),
        .c(new_Jinkela_wire_976)
    );

    spl2 new_Jinkela_splitter_7 (
        .a(new_Jinkela_wire_163),
        .b(new_Jinkela_wire_164),
        .c(new_Jinkela_wire_165)
    );

    bfr new_Jinkela_buffer_160 (
        .din(new_Jinkela_wire_175),
        .dout(new_Jinkela_wire_176)
    );

    bfr new_Jinkela_buffer_425 (
        .din(new_Jinkela_wire_476),
        .dout(new_Jinkela_wire_477)
    );

    bfr new_Jinkela_buffer_814 (
        .din(new_Jinkela_wire_963),
        .dout(new_Jinkela_wire_964)
    );

    bfr new_Jinkela_buffer_121 (
        .din(new_Jinkela_wire_132),
        .dout(new_Jinkela_wire_133)
    );

    bfr new_Jinkela_buffer_150 (
        .din(new_Jinkela_wire_165),
        .dout(new_Jinkela_wire_166)
    );

    bfr new_Jinkela_buffer_467 (
        .din(new_Jinkela_wire_520),
        .dout(new_Jinkela_wire_521)
    );

    spl2 new_Jinkela_splitter_68 (
        .a(_032_),
        .b(new_Jinkela_wire_948),
        .c(new_Jinkela_wire_949)
    );

    spl4L new_Jinkela_splitter_73 (
        .a(new_Jinkela_wire_977),
        .b(new_Jinkela_wire_978),
        .d(new_Jinkela_wire_979),
        .e(new_Jinkela_wire_980),
        .c(new_Jinkela_wire_981)
    );

    bfr new_Jinkela_buffer_476 (
        .din(new_Jinkela_wire_529),
        .dout(new_Jinkela_wire_530)
    );

    and_ii _143_ (
        .a(new_Jinkela_wire_982),
        .b(new_Jinkela_wire_41),
        .c(_087_)
    );

    or_bb _188_ (
        .a(_014_),
        .b(new_Jinkela_wire_714),
        .c(_015_)
    );

    bfr new_Jinkela_buffer_461 (
        .din(new_Jinkela_wire_514),
        .dout(new_Jinkela_wire_515)
    );

    bfr new_Jinkela_buffer_775 (
        .din(new_Jinkela_wire_914),
        .dout(new_Jinkela_wire_915)
    );

    or_bi _144_ (
        .a(new_Jinkela_wire_970),
        .b(new_Jinkela_wire_329),
        .c(_088_)
    );

    and_ii _189_ (
        .a(new_Jinkela_wire_716),
        .b(new_Jinkela_wire_164),
        .c(_016_)
    );

    bfr new_Jinkela_buffer_498 (
        .din(new_Jinkela_wire_553),
        .dout(new_Jinkela_wire_554)
    );

    or_ii _145_ (
        .a(_088_),
        .b(new_Jinkela_wire_258),
        .c(_089_)
    );

    and_bi _190_ (
        .a(new_Jinkela_wire_566),
        .b(new_Jinkela_wire_628),
        .c(_017_)
    );

    bfr new_Jinkela_buffer_477 (
        .din(new_Jinkela_wire_530),
        .dout(new_Jinkela_wire_531)
    );

    and_ii _146_ (
        .a(new_Jinkela_wire_907),
        .b(new_Jinkela_wire_341),
        .c(_090_)
    );

    or_bb _191_ (
        .a(_017_),
        .b(new_Jinkela_wire_947),
        .c(_018_)
    );

    bfr new_Jinkela_buffer_527 (
        .din(new_Jinkela_wire_590),
        .dout(new_Jinkela_wire_591)
    );

    or_bb _147_ (
        .a(_090_),
        .b(_087_),
        .c(_091_)
    );

    and_ii _192_ (
        .a(new_Jinkela_wire_760),
        .b(new_Jinkela_wire_381),
        .c(_019_)
    );

    bfr new_Jinkela_buffer_478 (
        .din(new_Jinkela_wire_531),
        .dout(new_Jinkela_wire_532)
    );

    and_bi _148_ (
        .a(_086_),
        .b(_091_),
        .c(_092_)
    );

    or_bb _193_ (
        .a(new_Jinkela_wire_740),
        .b(new_Jinkela_wire_801),
        .c(_020_)
    );

    bfr new_Jinkela_buffer_499 (
        .din(new_Jinkela_wire_554),
        .dout(new_Jinkela_wire_555)
    );

    bfr new_Jinkela_buffer_780 (
        .din(new_Jinkela_wire_921),
        .dout(new_Jinkela_wire_922)
    );

    or_bi _149_ (
        .a(new_Jinkela_wire_976),
        .b(new_Jinkela_wire_215),
        .c(_093_)
    );

    and_bi _194_ (
        .a(new_Jinkela_wire_142),
        .b(new_Jinkela_wire_630),
        .c(_021_)
    );

    bfr new_Jinkela_buffer_479 (
        .din(new_Jinkela_wire_532),
        .dout(new_Jinkela_wire_533)
    );

    or_ii _150_ (
        .a(_093_),
        .b(new_Jinkela_wire_577),
        .c(_094_)
    );

    or_bb _195_ (
        .a(_021_),
        .b(new_Jinkela_wire_937),
        .c(_022_)
    );

    bfr new_Jinkela_buffer_512 (
        .din(new_Jinkela_wire_571),
        .dout(new_Jinkela_wire_572)
    );

    and_ii _151_ (
        .a(new_Jinkela_wire_918),
        .b(new_Jinkela_wire_311),
        .c(_095_)
    );

    and_ii _196_ (
        .a(new_Jinkela_wire_694),
        .b(new_Jinkela_wire_444),
        .c(_023_)
    );

    bfr new_Jinkela_buffer_480 (
        .din(new_Jinkela_wire_533),
        .dout(new_Jinkela_wire_534)
    );

    or_bi _152_ (
        .a(new_Jinkela_wire_978),
        .b(new_Jinkela_wire_391),
        .c(_096_)
    );

    and_bi _197_ (
        .a(new_Jinkela_wire_618),
        .b(new_Jinkela_wire_620),
        .c(_024_)
    );

    bfr new_Jinkela_buffer_500 (
        .din(new_Jinkela_wire_555),
        .dout(new_Jinkela_wire_556)
    );

    or_ii _153_ (
        .a(_096_),
        .b(new_Jinkela_wire_588),
        .c(_097_)
    );

    or_bb _198_ (
        .a(_024_),
        .b(new_Jinkela_wire_898),
        .c(_025_)
    );

    bfr new_Jinkela_buffer_481 (
        .din(new_Jinkela_wire_534),
        .dout(new_Jinkela_wire_535)
    );

    bfr new_Jinkela_buffer_776 (
        .din(new_Jinkela_wire_915),
        .dout(new_Jinkela_wire_916)
    );

    and_ii _154_ (
        .a(new_Jinkela_wire_857),
        .b(new_Jinkela_wire_291),
        .c(_098_)
    );

    and_ii _199_ (
        .a(new_Jinkela_wire_683),
        .b(new_Jinkela_wire_475),
        .c(_026_)
    );

    bfr new_Jinkela_buffer_519 (
        .din(new_Jinkela_wire_580),
        .dout(new_Jinkela_wire_581)
    );

    or_bb _155_ (
        .a(_098_),
        .b(_095_),
        .c(_099_)
    );

    or_bb _200_ (
        .a(_026_),
        .b(_023_),
        .c(_027_)
    );

    bfr new_Jinkela_buffer_482 (
        .din(new_Jinkela_wire_535),
        .dout(new_Jinkela_wire_536)
    );

    or_bi _156_ (
        .a(new_Jinkela_wire_980),
        .b(new_Jinkela_wire_268),
        .c(_100_)
    );

    or_bb _201_ (
        .a(new_Jinkela_wire_739),
        .b(_020_),
        .c(_028_)
    );

    bfr new_Jinkela_buffer_501 (
        .din(new_Jinkela_wire_556),
        .dout(new_Jinkela_wire_557)
    );

    or_ii _157_ (
        .a(_100_),
        .b(new_Jinkela_wire_237),
        .c(_101_)
    );

    or_bb _202_ (
        .a(_028_),
        .b(new_Jinkela_wire_664),
        .c(_029_)
    );

    or_bb _165_ (
        .a(_108_),
        .b(_105_),
        .c(_109_)
    );

    spl2 new_Jinkela_splitter_27 (
        .a(new_Jinkela_wire_536),
        .b(new_Jinkela_wire_537),
        .c(new_Jinkela_wire_538)
    );

    and_ii _158_ (
        .a(new_Jinkela_wire_938),
        .b(new_Jinkela_wire_558),
        .c(_102_)
    );

    and_bi _203_ (
        .a(new_Jinkela_wire_967),
        .b(_029_),
        .c(_030_)
    );

    bfr new_Jinkela_buffer_483 (
        .din(new_Jinkela_wire_538),
        .dout(new_Jinkela_wire_539)
    );

    or_ii _159_ (
        .a(new_Jinkela_wire_971),
        .b(new_Jinkela_wire_29),
        .c(_103_)
    );

    inv _204_ (
        .din(new_Jinkela_wire_780),
        .dout(new_net_198)
    );

    bfr new_Jinkela_buffer_513 (
        .din(new_Jinkela_wire_572),
        .dout(new_Jinkela_wire_573)
    );

    and_bi _160_ (
        .a(_103_),
        .b(new_Jinkela_wire_675),
        .c(_104_)
    );

    inv _205_ (
        .din(new_Jinkela_wire_974),
        .dout(new_net_192)
    );

    spl2 new_Jinkela_splitter_28 (
        .a(new_Jinkela_wire_557),
        .b(new_Jinkela_wire_558),
        .c(new_Jinkela_wire_559)
    );

    and_ii _161_ (
        .a(new_Jinkela_wire_705),
        .b(new_Jinkela_wire_185),
        .c(_105_)
    );

    and_bi _206_ (
        .a(new_Jinkela_wire_422),
        .b(new_Jinkela_wire_786),
        .c(_031_)
    );

    bfr new_Jinkela_buffer_794 (
        .din(new_Jinkela_wire_939),
        .dout(new_Jinkela_wire_940)
    );

    bfr new_Jinkela_buffer_484 (
        .din(new_Jinkela_wire_539),
        .dout(new_Jinkela_wire_540)
    );

    or_bi _162_ (
        .a(new_Jinkela_wire_981),
        .b(new_Jinkela_wire_598),
        .c(_106_)
    );

    or_bb _207_ (
        .a(_031_),
        .b(new_Jinkela_wire_759),
        .c(_032_)
    );

    bfr new_Jinkela_buffer_502 (
        .din(new_Jinkela_wire_559),
        .dout(new_Jinkela_wire_560)
    );

    or_bb _166_ (
        .a(_109_),
        .b(new_Jinkela_wire_665),
        .c(_110_)
    );

    or_bi _208_ (
        .a(new_Jinkela_wire_787),
        .b(new_Jinkela_wire_111),
        .c(_033_)
    );

    bfr new_Jinkela_buffer_485 (
        .din(new_Jinkela_wire_540),
        .dout(new_Jinkela_wire_541)
    );

    or_bb _167_ (
        .a(_110_),
        .b(new_Jinkela_wire_727),
        .c(_111_)
    );

    and_bi _209_ (
        .a(_033_),
        .b(new_Jinkela_wire_837),
        .c(_034_)
    );

    and_bi _168_ (
        .a(new_Jinkela_wire_917),
        .b(_111_),
        .c(_112_)
    );

    or_bi _210_ (
        .a(new_Jinkela_wire_676),
        .b(new_Jinkela_wire_948),
        .c(_035_)
    );

    spl3L new_Jinkela_splitter_33 (
        .a(_112_),
        .b(new_Jinkela_wire_619),
        .d(new_Jinkela_wire_622),
        .c(new_Jinkela_wire_627)
    );

    bfr new_Jinkela_buffer_486 (
        .din(new_Jinkela_wire_541),
        .dout(new_Jinkela_wire_542)
    );

    and_bi _169_ (
        .a(new_Jinkela_wire_49),
        .b(new_Jinkela_wire_625),
        .c(_113_)
    );

    and_bi _211_ (
        .a(new_Jinkela_wire_453),
        .b(new_Jinkela_wire_782),
        .c(_036_)
    );

    bfr new_Jinkela_buffer_514 (
        .din(new_Jinkela_wire_573),
        .dout(new_Jinkela_wire_574)
    );

    or_bb _170_ (
        .a(_113_),
        .b(new_Jinkela_wire_991),
        .c(_114_)
    );

    and_ii _212_ (
        .a(_036_),
        .b(new_Jinkela_wire_704),
        .c(_037_)
    );

    bfr new_Jinkela_buffer_487 (
        .din(new_Jinkela_wire_542),
        .dout(new_Jinkela_wire_543)
    );

    or_bb _171_ (
        .a(new_Jinkela_wire_749),
        .b(new_Jinkela_wire_413),
        .c(_115_)
    );

    and_bi _213_ (
        .a(new_Jinkela_wire_781),
        .b(new_Jinkela_wire_769),
        .c(_038_)
    );

    bfr new_Jinkela_buffer_503 (
        .din(new_Jinkela_wire_560),
        .dout(new_Jinkela_wire_561)
    );

    and_bi _172_ (
        .a(new_Jinkela_wire_299),
        .b(new_Jinkela_wire_629),
        .c(_116_)
    );

    or_bb _214_ (
        .a(_038_),
        .b(new_Jinkela_wire_748),
        .c(_039_)
    );

    bfr new_Jinkela_buffer_488 (
        .din(new_Jinkela_wire_543),
        .dout(new_Jinkela_wire_544)
    );

    or_bb _173_ (
        .a(_116_),
        .b(new_Jinkela_wire_866),
        .c(_000_)
    );

    or_bb _215_ (
        .a(new_Jinkela_wire_968),
        .b(new_Jinkela_wire_899),
        .c(_040_)
    );

    bfr new_Jinkela_buffer_520 (
        .din(new_Jinkela_wire_581),
        .dout(new_Jinkela_wire_582)
    );

    and_ii _174_ (
        .a(new_Jinkela_wire_955),
        .b(new_Jinkela_wire_537),
        .c(_001_)
    );

    or_bb _216_ (
        .a(new_Jinkela_wire_993),
        .b(new_Jinkela_wire_813),
        .c(new_net_0)
    );

    bfr new_Jinkela_buffer_489 (
        .din(new_Jinkela_wire_544),
        .dout(new_Jinkela_wire_545)
    );

    and_bi _175_ (
        .a(new_Jinkela_wire_349),
        .b(new_Jinkela_wire_621),
        .c(_002_)
    );

    and_bi _217_ (
        .a(new_Jinkela_wire_80),
        .b(new_Jinkela_wire_777),
        .c(_041_)
    );

    bfr new_Jinkela_buffer_504 (
        .din(new_Jinkela_wire_561),
        .dout(new_Jinkela_wire_562)
    );

    or_bb _176_ (
        .a(_002_),
        .b(new_Jinkela_wire_916),
        .c(_003_)
    );

    or_bb _218_ (
        .a(_041_),
        .b(new_Jinkela_wire_856),
        .c(_042_)
    );

    bfr new_Jinkela_buffer_490 (
        .din(new_Jinkela_wire_545),
        .dout(new_Jinkela_wire_546)
    );

    and_ii _177_ (
        .a(new_Jinkela_wire_827),
        .b(new_Jinkela_wire_102),
        .c(_004_)
    );

    and_bi _219_ (
        .a(new_Jinkela_wire_173),
        .b(new_Jinkela_wire_778),
        .c(_043_)
    );

    bfr new_Jinkela_buffer_515 (
        .din(new_Jinkela_wire_574),
        .dout(new_Jinkela_wire_575)
    );

    or_bb _178_ (
        .a(_004_),
        .b(_001_),
        .c(_005_)
    );

    and_ii _220_ (
        .a(_043_),
        .b(new_Jinkela_wire_726),
        .c(_044_)
    );

    bfr new_Jinkela_buffer_505 (
        .din(new_Jinkela_wire_562),
        .dout(new_Jinkela_wire_563)
    );

    and_bi _179_ (
        .a(new_Jinkela_wire_902),
        .b(_005_),
        .c(_006_)
    );

    or_bi _221_ (
        .a(new_Jinkela_wire_903),
        .b(new_Jinkela_wire_816),
        .c(_045_)
    );

    bfr new_Jinkela_buffer_553 (
        .din(new_net_192),
        .dout(new_Jinkela_wire_632)
    );

    and_bi _180_ (
        .a(new_Jinkela_wire_319),
        .b(new_Jinkela_wire_623),
        .c(_007_)
    );

    and_bi _222_ (
        .a(new_Jinkela_wire_546),
        .b(new_Jinkela_wire_785),
        .c(_046_)
    );

    bfr new_Jinkela_buffer_506 (
        .din(new_Jinkela_wire_563),
        .dout(new_Jinkela_wire_564)
    );

    or_bb _181_ (
        .a(_007_),
        .b(new_Jinkela_wire_927),
        .c(_008_)
    );

    or_bb _223_ (
        .a(_046_),
        .b(new_Jinkela_wire_965),
        .c(_047_)
    );

    bfr new_Jinkela_buffer_516 (
        .din(new_Jinkela_wire_575),
        .dout(new_Jinkela_wire_576)
    );

    and_ii _182_ (
        .a(new_Jinkela_wire_802),
        .b(new_Jinkela_wire_506),
        .c(_009_)
    );

    and_bi _224_ (
        .a(new_Jinkela_wire_484),
        .b(new_Jinkela_wire_788),
        .c(_048_)
    );

    bfr new_Jinkela_buffer_507 (
        .din(new_Jinkela_wire_564),
        .dout(new_Jinkela_wire_565)
    );

    and_bi _183_ (
        .a(new_Jinkela_wire_19),
        .b(new_Jinkela_wire_626),
        .c(_010_)
    );

    or_bb _225_ (
        .a(_048_),
        .b(new_Jinkela_wire_693),
        .c(_049_)
    );

    bfr new_Jinkela_buffer_521 (
        .din(new_Jinkela_wire_582),
        .dout(new_Jinkela_wire_583)
    );

    or_bb _184_ (
        .a(_010_),
        .b(new_Jinkela_wire_798),
        .c(_011_)
    );

    or_ii _226_ (
        .a(new_Jinkela_wire_715),
        .b(new_Jinkela_wire_661),
        .c(_050_)
    );

    bfr new_Jinkela_buffer_508 (
        .din(new_Jinkela_wire_565),
        .dout(new_Jinkela_wire_566)
    );

    and_ii _185_ (
        .a(new_Jinkela_wire_846),
        .b(new_Jinkela_wire_71),
        .c(_012_)
    );

    or_bb _227_ (
        .a(new_Jinkela_wire_867),
        .b(new_Jinkela_wire_844),
        .c(_051_)
    );

    bfr new_Jinkela_buffer_517 (
        .din(new_Jinkela_wire_576),
        .dout(new_Jinkela_wire_577)
    );

    or_bb _186_ (
        .a(_012_),
        .b(_009_),
        .c(_013_)
    );

    or_bb _228_ (
        .a(new_Jinkela_wire_774),
        .b(new_Jinkela_wire_770),
        .c(_052_)
    );

    bfr new_Jinkela_buffer_528 (
        .din(new_Jinkela_wire_591),
        .dout(new_Jinkela_wire_592)
    );

    and_bi _187_ (
        .a(new_Jinkela_wire_193),
        .b(new_Jinkela_wire_624),
        .c(_014_)
    );

    or_bi _229_ (
        .a(new_Jinkela_wire_783),
        .b(new_Jinkela_wire_515),
        .c(_053_)
    );

    bfr new_Jinkela_buffer_38 (
        .din(new_Jinkela_wire_43),
        .dout(new_Jinkela_wire_44)
    );

    bfr new_Jinkela_buffer_242 (
        .din(new_Jinkela_wire_275),
        .dout(new_Jinkela_wire_276)
    );

    bfr new_Jinkela_buffer_380 (
        .din(new_Jinkela_wire_427),
        .dout(new_Jinkela_wire_428)
    );

    bfr new_Jinkela_buffer_522 (
        .din(new_Jinkela_wire_583),
        .dout(new_Jinkela_wire_584)
    );

    bfr new_Jinkela_buffer_632 (
        .din(new_Jinkela_wire_724),
        .dout(new_Jinkela_wire_725)
    );

    bfr new_Jinkela_buffer_744 (
        .din(new_Jinkela_wire_875),
        .dout(new_Jinkela_wire_876)
    );

    bfr new_Jinkela_buffer_76 (
        .din(new_Jinkela_wire_83),
        .dout(new_Jinkela_wire_84)
    );

    bfr new_Jinkela_buffer_265 (
        .din(new_Jinkela_wire_300),
        .dout(new_Jinkela_wire_301)
    );

    bfr new_Jinkela_buffer_357 (
        .din(new_Jinkela_wire_402),
        .dout(new_Jinkela_wire_403)
    );

    bfr new_Jinkela_buffer_536 (
        .din(new_Jinkela_wire_599),
        .dout(new_Jinkela_wire_600)
    );

    bfr new_Jinkela_buffer_580 (
        .din(new_Jinkela_wire_658),
        .dout(new_Jinkela_wire_659)
    );

    bfr new_Jinkela_buffer_616 (
        .din(new_Jinkela_wire_706),
        .dout(new_Jinkela_wire_707)
    );

    bfr new_Jinkela_buffer_39 (
        .din(new_Jinkela_wire_44),
        .dout(new_Jinkela_wire_45)
    );

    bfr new_Jinkela_buffer_243 (
        .din(new_Jinkela_wire_276),
        .dout(new_Jinkela_wire_277)
    );

    bfr new_Jinkela_buffer_434 (
        .din(new_Jinkela_wire_485),
        .dout(new_Jinkela_wire_486)
    );

    bfr new_Jinkela_buffer_523 (
        .din(new_Jinkela_wire_584),
        .dout(new_Jinkela_wire_585)
    );

    bfr new_Jinkela_buffer_633 (
        .din(new_Jinkela_wire_725),
        .dout(new_Jinkela_wire_726)
    );

    bfr new_Jinkela_buffer_645 (
        .din(new_Jinkela_wire_741),
        .dout(new_Jinkela_wire_742)
    );

    bfr new_Jinkela_buffer_51 (
        .din(new_Jinkela_wire_56),
        .dout(new_Jinkela_wire_57)
    );

    bfr new_Jinkela_buffer_249 (
        .din(new_Jinkela_wire_282),
        .dout(new_Jinkela_wire_283)
    );

    bfr new_Jinkela_buffer_358 (
        .din(new_Jinkela_wire_403),
        .dout(new_Jinkela_wire_404)
    );

    bfr new_Jinkela_buffer_529 (
        .din(new_Jinkela_wire_592),
        .dout(new_Jinkela_wire_593)
    );

    bfr new_Jinkela_buffer_581 (
        .din(new_Jinkela_wire_659),
        .dout(new_Jinkela_wire_660)
    );

    bfr new_Jinkela_buffer_601 (
        .din(new_Jinkela_wire_687),
        .dout(new_Jinkela_wire_688)
    );

    bfr new_Jinkela_buffer_40 (
        .din(new_Jinkela_wire_45),
        .dout(new_Jinkela_wire_46)
    );

    bfr new_Jinkela_buffer_244 (
        .din(new_Jinkela_wire_277),
        .dout(new_Jinkela_wire_278)
    );

    bfr new_Jinkela_buffer_381 (
        .din(new_Jinkela_wire_428),
        .dout(new_Jinkela_wire_429)
    );

    bfr new_Jinkela_buffer_524 (
        .din(new_Jinkela_wire_585),
        .dout(new_Jinkela_wire_586)
    );

    bfr new_Jinkela_buffer_746 (
        .din(new_Jinkela_wire_877),
        .dout(new_Jinkela_wire_878)
    );

    spl2 new_Jinkela_splitter_64 (
        .a(_089_),
        .b(new_Jinkela_wire_907),
        .c(new_Jinkela_wire_908)
    );

    bfr new_Jinkela_buffer_282 (
        .din(new_Jinkela_wire_321),
        .dout(new_Jinkela_wire_322)
    );

    bfr new_Jinkela_buffer_359 (
        .din(new_Jinkela_wire_404),
        .dout(new_Jinkela_wire_405)
    );

    bfr new_Jinkela_buffer_608 (
        .din(new_Jinkela_wire_696),
        .dout(new_Jinkela_wire_697)
    );

    bfr new_Jinkela_buffer_158 (
        .din(N73),
        .dout(new_Jinkela_wire_174)
    );

    bfr new_Jinkela_buffer_555 (
        .din(new_Jinkela_wire_633),
        .dout(new_Jinkela_wire_634)
    );

    bfr new_Jinkela_buffer_639 (
        .din(new_Jinkela_wire_733),
        .dout(new_Jinkela_wire_734)
    );

    bfr new_Jinkela_buffer_41 (
        .din(new_Jinkela_wire_46),
        .dout(new_Jinkela_wire_47)
    );

    bfr new_Jinkela_buffer_245 (
        .din(new_Jinkela_wire_278),
        .dout(new_Jinkela_wire_279)
    );

    bfr new_Jinkela_buffer_407 (
        .din(new_Jinkela_wire_456),
        .dout(new_Jinkela_wire_457)
    );

    bfr new_Jinkela_buffer_525 (
        .din(new_Jinkela_wire_586),
        .dout(new_Jinkela_wire_587)
    );

    bfr new_Jinkela_buffer_602 (
        .din(new_Jinkela_wire_688),
        .dout(new_Jinkela_wire_689)
    );

    spl2 new_Jinkela_splitter_47 (
        .a(_018_),
        .b(new_Jinkela_wire_760),
        .c(new_Jinkela_wire_761)
    );

    bfr new_Jinkela_buffer_52 (
        .din(new_Jinkela_wire_57),
        .dout(new_Jinkela_wire_58)
    );

    bfr new_Jinkela_buffer_250 (
        .din(new_Jinkela_wire_283),
        .dout(new_Jinkela_wire_284)
    );

    bfr new_Jinkela_buffer_360 (
        .din(new_Jinkela_wire_405),
        .dout(new_Jinkela_wire_406)
    );

    bfr new_Jinkela_buffer_530 (
        .din(new_Jinkela_wire_593),
        .dout(new_Jinkela_wire_594)
    );

    spl2 new_Jinkela_splitter_43 (
        .a(_015_),
        .b(new_Jinkela_wire_716),
        .c(new_Jinkela_wire_717)
    );

    bfr new_Jinkela_buffer_640 (
        .din(new_Jinkela_wire_734),
        .dout(new_Jinkela_wire_735)
    );

    bfr new_Jinkela_buffer_42 (
        .din(new_Jinkela_wire_47),
        .dout(new_Jinkela_wire_48)
    );

    bfr new_Jinkela_buffer_266 (
        .din(new_Jinkela_wire_301),
        .dout(new_Jinkela_wire_302)
    );

    bfr new_Jinkela_buffer_382 (
        .din(new_Jinkela_wire_429),
        .dout(new_Jinkela_wire_430)
    );

    bfr new_Jinkela_buffer_526 (
        .din(new_Jinkela_wire_587),
        .dout(new_Jinkela_wire_588)
    );

    bfr new_Jinkela_buffer_603 (
        .din(new_Jinkela_wire_689),
        .dout(new_Jinkela_wire_690)
    );

    spl2 new_Jinkela_splitter_48 (
        .a(new_net_0),
        .b(new_Jinkela_wire_770),
        .c(new_Jinkela_wire_771)
    );

    bfr new_Jinkela_buffer_77 (
        .din(new_Jinkela_wire_84),
        .dout(new_Jinkela_wire_85)
    );

    bfr new_Jinkela_buffer_251 (
        .din(new_Jinkela_wire_284),
        .dout(new_Jinkela_wire_285)
    );

    bfr new_Jinkela_buffer_361 (
        .din(new_Jinkela_wire_406),
        .dout(new_Jinkela_wire_407)
    );

    bfr new_Jinkela_buffer_537 (
        .din(new_Jinkela_wire_600),
        .dout(new_Jinkela_wire_601)
    );

    bfr new_Jinkela_buffer_609 (
        .din(new_Jinkela_wire_697),
        .dout(new_Jinkela_wire_698)
    );

    bfr new_Jinkela_buffer_641 (
        .din(new_Jinkela_wire_735),
        .dout(new_Jinkela_wire_736)
    );

    bfr new_Jinkela_buffer_43 (
        .din(new_Jinkela_wire_48),
        .dout(new_Jinkela_wire_49)
    );

    bfr new_Jinkela_buffer_531 (
        .din(new_Jinkela_wire_594),
        .dout(new_Jinkela_wire_595)
    );

    bfr new_Jinkela_buffer_604 (
        .din(new_Jinkela_wire_690),
        .dout(new_Jinkela_wire_691)
    );

    spl2 new_Jinkela_splitter_21 (
        .a(N30),
        .b(new_Jinkela_wire_350),
        .c(new_Jinkela_wire_351)
    );

    bfr new_Jinkela_buffer_646 (
        .din(new_Jinkela_wire_742),
        .dout(new_Jinkela_wire_743)
    );

    bfr new_Jinkela_buffer_749 (
        .din(new_Jinkela_wire_880),
        .dout(new_Jinkela_wire_881)
    );

    bfr new_Jinkela_buffer_53 (
        .din(new_Jinkela_wire_58),
        .dout(new_Jinkela_wire_59)
    );

    bfr new_Jinkela_buffer_252 (
        .din(new_Jinkela_wire_285),
        .dout(new_Jinkela_wire_286)
    );

    bfr new_Jinkela_buffer_362 (
        .din(new_Jinkela_wire_407),
        .dout(new_Jinkela_wire_408)
    );

    bfr new_Jinkela_buffer_582 (
        .din(_013_),
        .dout(new_Jinkela_wire_663)
    );

    bfr new_Jinkela_buffer_625 (
        .din(new_Jinkela_wire_717),
        .dout(new_Jinkela_wire_718)
    );

    bfr new_Jinkela_buffer_634 (
        .din(_099_),
        .dout(new_Jinkela_wire_727)
    );

    bfr new_Jinkela_buffer_103 (
        .din(new_Jinkela_wire_114),
        .dout(new_Jinkela_wire_115)
    );

    bfr new_Jinkela_buffer_267 (
        .din(new_Jinkela_wire_302),
        .dout(new_Jinkela_wire_303)
    );

    bfr new_Jinkela_buffer_383 (
        .din(new_Jinkela_wire_430),
        .dout(new_Jinkela_wire_431)
    );

    bfr new_Jinkela_buffer_532 (
        .din(new_Jinkela_wire_595),
        .dout(new_Jinkela_wire_596)
    );

    bfr new_Jinkela_buffer_605 (
        .din(new_Jinkela_wire_691),
        .dout(new_Jinkela_wire_692)
    );

    bfr new_Jinkela_buffer_647 (
        .din(new_Jinkela_wire_743),
        .dout(new_Jinkela_wire_744)
    );

    bfr new_Jinkela_buffer_54 (
        .din(new_Jinkela_wire_59),
        .dout(new_Jinkela_wire_60)
    );

    bfr new_Jinkela_buffer_253 (
        .din(new_Jinkela_wire_286),
        .dout(new_Jinkela_wire_287)
    );

    bfr new_Jinkela_buffer_363 (
        .din(new_Jinkela_wire_408),
        .dout(new_Jinkela_wire_409)
    );

    bfr new_Jinkela_buffer_538 (
        .din(new_Jinkela_wire_601),
        .dout(new_Jinkela_wire_602)
    );

    bfr new_Jinkela_buffer_610 (
        .din(new_Jinkela_wire_698),
        .dout(new_Jinkela_wire_699)
    );

    bfr new_Jinkela_buffer_750 (
        .din(new_Jinkela_wire_881),
        .dout(new_Jinkela_wire_882)
    );

    bfr new_Jinkela_buffer_78 (
        .din(new_Jinkela_wire_85),
        .dout(new_Jinkela_wire_86)
    );

    bfr new_Jinkela_buffer_408 (
        .din(new_Jinkela_wire_457),
        .dout(new_Jinkela_wire_458)
    );

    bfr new_Jinkela_buffer_533 (
        .din(new_Jinkela_wire_596),
        .dout(new_Jinkela_wire_597)
    );

    bfr new_Jinkela_buffer_316 (
        .din(N66),
        .dout(new_Jinkela_wire_360)
    );

    bfr new_Jinkela_buffer_606 (
        .din(new_Jinkela_wire_692),
        .dout(new_Jinkela_wire_693)
    );

    bfr new_Jinkela_buffer_648 (
        .din(new_Jinkela_wire_744),
        .dout(new_Jinkela_wire_745)
    );

    bfr new_Jinkela_buffer_55 (
        .din(new_Jinkela_wire_60),
        .dout(new_Jinkela_wire_61)
    );

    bfr new_Jinkela_buffer_254 (
        .din(new_Jinkela_wire_287),
        .dout(new_Jinkela_wire_288)
    );

    bfr new_Jinkela_buffer_364 (
        .din(new_Jinkela_wire_409),
        .dout(new_Jinkela_wire_410)
    );

    spl2 new_Jinkela_splitter_34 (
        .a(new_Jinkela_wire_619),
        .b(new_Jinkela_wire_620),
        .c(new_Jinkela_wire_621)
    );

    bfr new_Jinkela_buffer_617 (
        .din(new_Jinkela_wire_707),
        .dout(new_Jinkela_wire_708)
    );

    bfr new_Jinkela_buffer_653 (
        .din(new_Jinkela_wire_751),
        .dout(new_Jinkela_wire_752)
    );

    bfr new_Jinkela_buffer_112 (
        .din(new_Jinkela_wire_123),
        .dout(new_Jinkela_wire_124)
    );

    bfr new_Jinkela_buffer_268 (
        .din(new_Jinkela_wire_303),
        .dout(new_Jinkela_wire_304)
    );

    bfr new_Jinkela_buffer_384 (
        .din(new_Jinkela_wire_431),
        .dout(new_Jinkela_wire_432)
    );

    bfr new_Jinkela_buffer_534 (
        .din(new_Jinkela_wire_597),
        .dout(new_Jinkela_wire_598)
    );

    bfr new_Jinkela_buffer_611 (
        .din(new_Jinkela_wire_699),
        .dout(new_Jinkela_wire_700)
    );

    bfr new_Jinkela_buffer_649 (
        .din(new_Jinkela_wire_745),
        .dout(new_Jinkela_wire_746)
    );

    bfr new_Jinkela_buffer_56 (
        .din(new_Jinkela_wire_61),
        .dout(new_Jinkela_wire_62)
    );

    bfr new_Jinkela_buffer_255 (
        .din(new_Jinkela_wire_288),
        .dout(new_Jinkela_wire_289)
    );

    bfr new_Jinkela_buffer_365 (
        .din(new_Jinkela_wire_410),
        .dout(new_Jinkela_wire_411)
    );

    bfr new_Jinkela_buffer_539 (
        .din(new_Jinkela_wire_602),
        .dout(new_Jinkela_wire_603)
    );

    bfr new_Jinkela_buffer_669 (
        .din(new_Jinkela_wire_771),
        .dout(new_Jinkela_wire_772)
    );

    bfr new_Jinkela_buffer_671 (
        .din(_051_),
        .dout(new_Jinkela_wire_774)
    );

    bfr new_Jinkela_buffer_79 (
        .din(new_Jinkela_wire_86),
        .dout(new_Jinkela_wire_87)
    );

    bfr new_Jinkela_buffer_283 (
        .din(new_Jinkela_wire_322),
        .dout(new_Jinkela_wire_323)
    );

    bfr new_Jinkela_buffer_435 (
        .din(new_Jinkela_wire_486),
        .dout(new_Jinkela_wire_487)
    );

    spl4L new_Jinkela_splitter_35 (
        .a(new_Jinkela_wire_622),
        .b(new_Jinkela_wire_623),
        .d(new_Jinkela_wire_624),
        .e(new_Jinkela_wire_625),
        .c(new_Jinkela_wire_626)
    );

    spl2 new_Jinkela_splitter_37 (
        .a(_047_),
        .b(new_Jinkela_wire_661),
        .c(new_Jinkela_wire_662)
    );

    bfr new_Jinkela_buffer_612 (
        .din(new_Jinkela_wire_700),
        .dout(new_Jinkela_wire_701)
    );

    bfr new_Jinkela_buffer_57 (
        .din(new_Jinkela_wire_62),
        .dout(new_Jinkela_wire_63)
    );

    bfr new_Jinkela_buffer_256 (
        .din(new_Jinkela_wire_289),
        .dout(new_Jinkela_wire_290)
    );

    bfr new_Jinkela_buffer_366 (
        .din(new_Jinkela_wire_411),
        .dout(new_Jinkela_wire_412)
    );

    bfr new_Jinkela_buffer_540 (
        .din(new_Jinkela_wire_603),
        .dout(new_Jinkela_wire_604)
    );

    bfr new_Jinkela_buffer_618 (
        .din(new_Jinkela_wire_708),
        .dout(new_Jinkela_wire_709)
    );

    bfr new_Jinkela_buffer_654 (
        .din(new_Jinkela_wire_752),
        .dout(new_Jinkela_wire_753)
    );

    bfr new_Jinkela_buffer_104 (
        .din(new_Jinkela_wire_115),
        .dout(new_Jinkela_wire_116)
    );

    bfr new_Jinkela_buffer_269 (
        .din(new_Jinkela_wire_304),
        .dout(new_Jinkela_wire_305)
    );

    bfr new_Jinkela_buffer_385 (
        .din(new_Jinkela_wire_432),
        .dout(new_Jinkela_wire_433)
    );

    spl4L new_Jinkela_splitter_36 (
        .a(new_Jinkela_wire_627),
        .b(new_Jinkela_wire_628),
        .d(new_Jinkela_wire_629),
        .e(new_Jinkela_wire_630),
        .c(new_Jinkela_wire_631)
    );

    bfr new_Jinkela_buffer_613 (
        .din(new_Jinkela_wire_701),
        .dout(new_Jinkela_wire_702)
    );

    bfr new_Jinkela_buffer_651 (
        .din(new_Jinkela_wire_747),
        .dout(new_Jinkela_wire_748)
    );

    bfr new_Jinkela_buffer_58 (
        .din(new_Jinkela_wire_63),
        .dout(new_Jinkela_wire_64)
    );

    spl2 new_Jinkela_splitter_17 (
        .a(new_Jinkela_wire_290),
        .b(new_Jinkela_wire_291),
        .c(new_Jinkela_wire_292)
    );

    spl2 new_Jinkela_splitter_23 (
        .a(new_Jinkela_wire_412),
        .b(new_Jinkela_wire_413),
        .c(new_Jinkela_wire_414)
    );

    bfr new_Jinkela_buffer_541 (
        .din(new_Jinkela_wire_604),
        .dout(new_Jinkela_wire_605)
    );

    spl2 new_Jinkela_splitter_44 (
        .a(_061_),
        .b(new_Jinkela_wire_728),
        .c(new_Jinkela_wire_729)
    );

    bfr new_Jinkela_buffer_754 (
        .din(new_Jinkela_wire_885),
        .dout(new_Jinkela_wire_886)
    );

    bfr new_Jinkela_buffer_80 (
        .din(new_Jinkela_wire_87),
        .dout(new_Jinkela_wire_88)
    );

    bfr new_Jinkela_buffer_257 (
        .din(new_Jinkela_wire_292),
        .dout(new_Jinkela_wire_293)
    );

    bfr new_Jinkela_buffer_367 (
        .din(new_Jinkela_wire_414),
        .dout(new_Jinkela_wire_415)
    );

    bfr new_Jinkela_buffer_554 (
        .din(new_Jinkela_wire_632),
        .dout(new_Jinkela_wire_633)
    );

    bfr new_Jinkela_buffer_614 (
        .din(new_Jinkela_wire_702),
        .dout(new_Jinkela_wire_703)
    );

    bfr new_Jinkela_buffer_655 (
        .din(new_Jinkela_wire_753),
        .dout(new_Jinkela_wire_754)
    );

    bfr new_Jinkela_buffer_59 (
        .din(new_Jinkela_wire_64),
        .dout(new_Jinkela_wire_65)
    );

    bfr new_Jinkela_buffer_291 (
        .din(new_Jinkela_wire_330),
        .dout(new_Jinkela_wire_331)
    );

    bfr new_Jinkela_buffer_409 (
        .din(new_Jinkela_wire_458),
        .dout(new_Jinkela_wire_459)
    );

    bfr new_Jinkela_buffer_542 (
        .din(new_Jinkela_wire_605),
        .dout(new_Jinkela_wire_606)
    );

    bfr new_Jinkela_buffer_619 (
        .din(new_Jinkela_wire_709),
        .dout(new_Jinkela_wire_710)
    );

    bfr new_Jinkela_buffer_662 (
        .din(new_Jinkela_wire_762),
        .dout(new_Jinkela_wire_763)
    );

    bfr new_Jinkela_buffer_270 (
        .din(new_Jinkela_wire_305),
        .dout(new_Jinkela_wire_306)
    );

    bfr new_Jinkela_buffer_386 (
        .din(new_Jinkela_wire_433),
        .dout(new_Jinkela_wire_434)
    );

    bfr new_Jinkela_buffer_615 (
        .din(new_Jinkela_wire_703),
        .dout(new_Jinkela_wire_704)
    );

    bfr new_Jinkela_buffer_176 (
        .din(N24),
        .dout(new_Jinkela_wire_194)
    );

    bfr new_Jinkela_buffer_656 (
        .din(new_Jinkela_wire_754),
        .dout(new_Jinkela_wire_755)
    );

    bfr new_Jinkela_buffer_756 (
        .din(new_Jinkela_wire_887),
        .dout(new_Jinkela_wire_888)
    );

    bfr new_Jinkela_buffer_60 (
        .din(new_Jinkela_wire_65),
        .dout(new_Jinkela_wire_66)
    );

    bfr new_Jinkela_buffer_258 (
        .din(new_Jinkela_wire_293),
        .dout(new_Jinkela_wire_294)
    );

    bfr new_Jinkela_buffer_368 (
        .din(new_Jinkela_wire_415),
        .dout(new_Jinkela_wire_416)
    );

    bfr new_Jinkela_buffer_543 (
        .din(new_Jinkela_wire_606),
        .dout(new_Jinkela_wire_607)
    );

    bfr new_Jinkela_buffer_635 (
        .din(new_Jinkela_wire_729),
        .dout(new_Jinkela_wire_730)
    );

    bfr new_Jinkela_buffer_642 (
        .din(_064_),
        .dout(new_Jinkela_wire_737)
    );

    bfr new_Jinkela_buffer_81 (
        .din(new_Jinkela_wire_88),
        .dout(new_Jinkela_wire_89)
    );

    bfr new_Jinkela_buffer_284 (
        .din(new_Jinkela_wire_323),
        .dout(new_Jinkela_wire_324)
    );

    bfr new_Jinkela_buffer_463 (
        .din(new_Jinkela_wire_516),
        .dout(new_Jinkela_wire_517)
    );

    bfr new_Jinkela_buffer_583 (
        .din(new_Jinkela_wire_663),
        .dout(new_Jinkela_wire_664)
    );

    bfr new_Jinkela_buffer_620 (
        .din(new_Jinkela_wire_710),
        .dout(new_Jinkela_wire_711)
    );

    bfr new_Jinkela_buffer_657 (
        .din(new_Jinkela_wire_755),
        .dout(new_Jinkela_wire_756)
    );

    bfr new_Jinkela_buffer_61 (
        .din(new_Jinkela_wire_66),
        .dout(new_Jinkela_wire_67)
    );

    bfr new_Jinkela_buffer_259 (
        .din(new_Jinkela_wire_294),
        .dout(new_Jinkela_wire_295)
    );

    bfr new_Jinkela_buffer_369 (
        .din(new_Jinkela_wire_416),
        .dout(new_Jinkela_wire_417)
    );

    bfr new_Jinkela_buffer_544 (
        .din(new_Jinkela_wire_607),
        .dout(new_Jinkela_wire_608)
    );

    bfr new_Jinkela_buffer_626 (
        .din(new_Jinkela_wire_718),
        .dout(new_Jinkela_wire_719)
    );

    bfr new_Jinkela_buffer_663 (
        .din(new_Jinkela_wire_763),
        .dout(new_Jinkela_wire_764)
    );

    bfr new_Jinkela_buffer_105 (
        .din(new_Jinkela_wire_116),
        .dout(new_Jinkela_wire_117)
    );

    bfr new_Jinkela_buffer_271 (
        .din(new_Jinkela_wire_306),
        .dout(new_Jinkela_wire_307)
    );

    bfr new_Jinkela_buffer_387 (
        .din(new_Jinkela_wire_434),
        .dout(new_Jinkela_wire_435)
    );

    bfr new_Jinkela_buffer_556 (
        .din(new_Jinkela_wire_634),
        .dout(new_Jinkela_wire_635)
    );

    bfr new_Jinkela_buffer_621 (
        .din(new_Jinkela_wire_711),
        .dout(new_Jinkela_wire_712)
    );

    bfr new_Jinkela_buffer_658 (
        .din(new_Jinkela_wire_756),
        .dout(new_Jinkela_wire_757)
    );

    bfr new_Jinkela_buffer_62 (
        .din(new_Jinkela_wire_67),
        .dout(new_Jinkela_wire_68)
    );

    bfr new_Jinkela_buffer_260 (
        .din(new_Jinkela_wire_295),
        .dout(new_Jinkela_wire_296)
    );

    bfr new_Jinkela_buffer_370 (
        .din(new_Jinkela_wire_417),
        .dout(new_Jinkela_wire_418)
    );

    bfr new_Jinkela_buffer_545 (
        .din(new_Jinkela_wire_608),
        .dout(new_Jinkela_wire_609)
    );

    spl3L new_Jinkela_splitter_49 (
        .a(_030_),
        .b(new_Jinkela_wire_776),
        .d(new_Jinkela_wire_779),
        .c(new_Jinkela_wire_784)
    );

    bfr new_Jinkela_buffer_771 (
        .din(new_Jinkela_wire_910),
        .dout(new_Jinkela_wire_911)
    );

    bfr new_Jinkela_buffer_82 (
        .din(new_Jinkela_wire_89),
        .dout(new_Jinkela_wire_90)
    );

    bfr new_Jinkela_buffer_410 (
        .din(new_Jinkela_wire_459),
        .dout(new_Jinkela_wire_460)
    );

    bfr new_Jinkela_buffer_622 (
        .din(new_Jinkela_wire_712),
        .dout(new_Jinkela_wire_713)
    );

    bfr new_Jinkela_buffer_308 (
        .din(new_Jinkela_wire_351),
        .dout(new_Jinkela_wire_352)
    );

    bfr new_Jinkela_buffer_584 (
        .din(_102_),
        .dout(new_Jinkela_wire_665)
    );

    bfr new_Jinkela_buffer_659 (
        .din(new_Jinkela_wire_757),
        .dout(new_Jinkela_wire_758)
    );

    bfr new_Jinkela_buffer_63 (
        .din(new_Jinkela_wire_68),
        .dout(new_Jinkela_wire_69)
    );

    bfr new_Jinkela_buffer_261 (
        .din(new_Jinkela_wire_296),
        .dout(new_Jinkela_wire_297)
    );

    bfr new_Jinkela_buffer_371 (
        .din(new_Jinkela_wire_418),
        .dout(new_Jinkela_wire_419)
    );

    spl2 new_Jinkela_splitter_32 (
        .a(new_Jinkela_wire_609),
        .b(new_Jinkela_wire_610),
        .c(new_Jinkela_wire_611)
    );

    bfr new_Jinkela_buffer_627 (
        .din(new_Jinkela_wire_719),
        .dout(new_Jinkela_wire_720)
    );

    bfr new_Jinkela_buffer_664 (
        .din(new_Jinkela_wire_764),
        .dout(new_Jinkela_wire_765)
    );

    bfr new_Jinkela_buffer_113 (
        .din(new_Jinkela_wire_124),
        .dout(new_Jinkela_wire_125)
    );

    bfr new_Jinkela_buffer_272 (
        .din(new_Jinkela_wire_307),
        .dout(new_Jinkela_wire_308)
    );

    bfr new_Jinkela_buffer_388 (
        .din(new_Jinkela_wire_435),
        .dout(new_Jinkela_wire_436)
    );

    bfr new_Jinkela_buffer_546 (
        .din(new_Jinkela_wire_611),
        .dout(new_Jinkela_wire_612)
    );

    bfr new_Jinkela_buffer_623 (
        .din(new_Jinkela_wire_713),
        .dout(new_Jinkela_wire_714)
    );

    bfr new_Jinkela_buffer_660 (
        .din(new_Jinkela_wire_758),
        .dout(new_Jinkela_wire_759)
    );

    bfr new_Jinkela_buffer_64 (
        .din(new_Jinkela_wire_69),
        .dout(new_Jinkela_wire_70)
    );

    bfr new_Jinkela_buffer_262 (
        .din(new_Jinkela_wire_297),
        .dout(new_Jinkela_wire_298)
    );

    bfr new_Jinkela_buffer_372 (
        .din(new_Jinkela_wire_419),
        .dout(new_Jinkela_wire_420)
    );

    bfr new_Jinkela_buffer_557 (
        .din(new_Jinkela_wire_635),
        .dout(new_Jinkela_wire_636)
    );

    bfr new_Jinkela_buffer_643 (
        .din(_074_),
        .dout(new_Jinkela_wire_738)
    );

    bfr new_Jinkela_buffer_670 (
        .din(new_Jinkela_wire_772),
        .dout(new_Jinkela_wire_773)
    );

    bfr new_Jinkela_buffer_83 (
        .din(new_Jinkela_wire_90),
        .dout(new_Jinkela_wire_91)
    );

    bfr new_Jinkela_buffer_285 (
        .din(new_Jinkela_wire_324),
        .dout(new_Jinkela_wire_325)
    );

    bfr new_Jinkela_buffer_436 (
        .din(new_Jinkela_wire_487),
        .dout(new_Jinkela_wire_488)
    );

    bfr new_Jinkela_buffer_585 (
        .din(_070_),
        .dout(new_Jinkela_wire_666)
    );

    bfr new_Jinkela_buffer_628 (
        .din(new_Jinkela_wire_720),
        .dout(new_Jinkela_wire_721)
    );

    bfr new_Jinkela_buffer_665 (
        .din(new_Jinkela_wire_765),
        .dout(new_Jinkela_wire_766)
    );

    spl2 new_Jinkela_splitter_3 (
        .a(new_Jinkela_wire_70),
        .b(new_Jinkela_wire_71),
        .c(new_Jinkela_wire_72)
    );

    bfr new_Jinkela_buffer_263 (
        .din(new_Jinkela_wire_298),
        .dout(new_Jinkela_wire_299)
    );

    bfr new_Jinkela_buffer_373 (
        .din(new_Jinkela_wire_420),
        .dout(new_Jinkela_wire_421)
    );

    bfr new_Jinkela_buffer_547 (
        .din(new_Jinkela_wire_612),
        .dout(new_Jinkela_wire_613)
    );

    bfr new_Jinkela_buffer_644 (
        .din(_027_),
        .dout(new_Jinkela_wire_739)
    );

    bfr new_Jinkela_buffer_774 (
        .din(new_Jinkela_wire_913),
        .dout(new_Jinkela_wire_914)
    );

    bfr new_Jinkela_buffer_273 (
        .din(new_Jinkela_wire_308),
        .dout(new_Jinkela_wire_309)
    );

    bfr new_Jinkela_buffer_65 (
        .din(new_Jinkela_wire_72),
        .dout(new_Jinkela_wire_73)
    );

    bfr new_Jinkela_buffer_389 (
        .din(new_Jinkela_wire_436),
        .dout(new_Jinkela_wire_437)
    );

    bfr new_Jinkela_buffer_558 (
        .din(new_Jinkela_wire_636),
        .dout(new_Jinkela_wire_637)
    );

    bfr new_Jinkela_buffer_629 (
        .din(new_Jinkela_wire_721),
        .dout(new_Jinkela_wire_722)
    );

    bfr new_Jinkela_buffer_666 (
        .din(new_Jinkela_wire_766),
        .dout(new_Jinkela_wire_767)
    );

    bfr new_Jinkela_buffer_106 (
        .din(new_Jinkela_wire_117),
        .dout(new_Jinkela_wire_118)
    );

    bfr new_Jinkela_buffer_292 (
        .din(new_Jinkela_wire_331),
        .dout(new_Jinkela_wire_332)
    );

    bfr new_Jinkela_buffer_374 (
        .din(new_Jinkela_wire_421),
        .dout(new_Jinkela_wire_422)
    );

    bfr new_Jinkela_buffer_548 (
        .din(new_Jinkela_wire_613),
        .dout(new_Jinkela_wire_614)
    );

    bfr new_Jinkela_buffer_636 (
        .din(new_Jinkela_wire_730),
        .dout(new_Jinkela_wire_731)
    );

    spl4L new_Jinkela_splitter_51 (
        .a(new_Jinkela_wire_779),
        .b(new_Jinkela_wire_780),
        .d(new_Jinkela_wire_781),
        .e(new_Jinkela_wire_782),
        .c(new_Jinkela_wire_783)
    );

    bfr new_Jinkela_buffer_84 (
        .din(new_Jinkela_wire_91),
        .dout(new_Jinkela_wire_92)
    );

    bfr new_Jinkela_buffer_274 (
        .din(new_Jinkela_wire_309),
        .dout(new_Jinkela_wire_310)
    );

    bfr new_Jinkela_buffer_411 (
        .din(new_Jinkela_wire_460),
        .dout(new_Jinkela_wire_461)
    );

    spl2 new_Jinkela_splitter_38 (
        .a(_069_),
        .b(new_Jinkela_wire_667),
        .c(new_Jinkela_wire_668)
    );

    bfr new_Jinkela_buffer_630 (
        .din(new_Jinkela_wire_722),
        .dout(new_Jinkela_wire_723)
    );

    bfr new_Jinkela_buffer_667 (
        .din(new_Jinkela_wire_767),
        .dout(new_Jinkela_wire_768)
    );

    bfr new_Jinkela_buffer_66 (
        .din(new_Jinkela_wire_73),
        .dout(new_Jinkela_wire_74)
    );

    bfr new_Jinkela_buffer_286 (
        .din(new_Jinkela_wire_325),
        .dout(new_Jinkela_wire_326)
    );

    bfr new_Jinkela_buffer_390 (
        .din(new_Jinkela_wire_437),
        .dout(new_Jinkela_wire_438)
    );

    bfr new_Jinkela_buffer_549 (
        .din(new_Jinkela_wire_614),
        .dout(new_Jinkela_wire_615)
    );

    spl2 new_Jinkela_splitter_45 (
        .a(_019_),
        .b(new_Jinkela_wire_740),
        .c(new_Jinkela_wire_741)
    );

    spl2 new_Jinkela_splitter_53 (
        .a(_084_),
        .b(new_Jinkela_wire_789),
        .c(new_Jinkela_wire_790)
    );

    bfr new_Jinkela_buffer_130 (
        .din(new_Jinkela_wire_143),
        .dout(new_Jinkela_wire_144)
    );

    spl2 new_Jinkela_splitter_18 (
        .a(new_Jinkela_wire_310),
        .b(new_Jinkela_wire_311),
        .c(new_Jinkela_wire_312)
    );

    bfr new_Jinkela_buffer_509 (
        .din(new_Jinkela_wire_568),
        .dout(new_Jinkela_wire_569)
    );

    bfr new_Jinkela_buffer_559 (
        .din(new_Jinkela_wire_637),
        .dout(new_Jinkela_wire_638)
    );

    spl2 new_Jinkela_splitter_39 (
        .a(_034_),
        .b(new_Jinkela_wire_676),
        .c(new_Jinkela_wire_677)
    );

    bfr new_Jinkela_buffer_631 (
        .din(new_Jinkela_wire_723),
        .dout(new_Jinkela_wire_724)
    );

    bfr new_Jinkela_buffer_67 (
        .din(new_Jinkela_wire_74),
        .dout(new_Jinkela_wire_75)
    );

    bfr new_Jinkela_buffer_275 (
        .din(new_Jinkela_wire_312),
        .dout(new_Jinkela_wire_313)
    );

    bfr new_Jinkela_buffer_391 (
        .din(new_Jinkela_wire_438),
        .dout(new_Jinkela_wire_439)
    );

    bfr new_Jinkela_buffer_550 (
        .din(new_Jinkela_wire_615),
        .dout(new_Jinkela_wire_616)
    );

    bfr new_Jinkela_buffer_637 (
        .din(new_Jinkela_wire_731),
        .dout(new_Jinkela_wire_732)
    );

    spl2 new_Jinkela_splitter_50 (
        .a(new_Jinkela_wire_776),
        .b(new_Jinkela_wire_777),
        .c(new_Jinkela_wire_778)
    );

    bfr new_Jinkela_buffer_781 (
        .din(new_Jinkela_wire_922),
        .dout(new_Jinkela_wire_923)
    );

    and_ii _164_ (
        .a(new_Jinkela_wire_928),
        .b(new_Jinkela_wire_134),
        .c(_108_)
    );

    bfr new_Jinkela_buffer_6 (
        .din(new_Jinkela_wire_5),
        .dout(new_Jinkela_wire_6)
    );

    bfr new_Jinkela_buffer_187 (
        .din(new_Jinkela_wire_208),
        .dout(new_Jinkela_wire_209)
    );

    bfr new_Jinkela_buffer_206 (
        .din(new_Jinkela_wire_231),
        .dout(new_Jinkela_wire_232)
    );

    spl2 new_Jinkela_splitter_8 (
        .a(new_Jinkela_wire_184),
        .b(new_Jinkela_wire_185),
        .c(new_Jinkela_wire_186)
    );

    bfr new_Jinkela_buffer_20 (
        .din(new_Jinkela_wire_23),
        .dout(new_Jinkela_wire_24)
    );

    bfr new_Jinkela_buffer_202 (
        .din(new_Jinkela_wire_225),
        .dout(new_Jinkela_wire_226)
    );

    bfr new_Jinkela_buffer_151 (
        .din(new_Jinkela_wire_166),
        .dout(new_Jinkela_wire_167)
    );

    bfr new_Jinkela_buffer_7 (
        .din(new_Jinkela_wire_6),
        .dout(new_Jinkela_wire_7)
    );

    bfr new_Jinkela_buffer_213 (
        .din(new_Jinkela_wire_240),
        .dout(new_Jinkela_wire_241)
    );

    bfr new_Jinkela_buffer_207 (
        .din(new_Jinkela_wire_232),
        .dout(new_Jinkela_wire_233)
    );

    bfr new_Jinkela_buffer_169 (
        .din(new_Jinkela_wire_186),
        .dout(new_Jinkela_wire_187)
    );

    spl2 new_Jinkela_splitter_5 (
        .a(N43),
        .b(new_Jinkela_wire_112),
        .c(new_Jinkela_wire_113)
    );

    bfr new_Jinkela_buffer_8 (
        .din(new_Jinkela_wire_7),
        .dout(new_Jinkela_wire_8)
    );

    bfr new_Jinkela_buffer_152 (
        .din(new_Jinkela_wire_167),
        .dout(new_Jinkela_wire_168)
    );

    bfr new_Jinkela_buffer_237 (
        .din(N63),
        .dout(new_Jinkela_wire_269)
    );

    bfr new_Jinkela_buffer_181 (
        .din(new_Jinkela_wire_200),
        .dout(new_Jinkela_wire_201)
    );

    bfr new_Jinkela_buffer_21 (
        .din(new_Jinkela_wire_24),
        .dout(new_Jinkela_wire_25)
    );

    bfr new_Jinkela_buffer_208 (
        .din(new_Jinkela_wire_233),
        .dout(new_Jinkela_wire_234)
    );

    bfr new_Jinkela_buffer_153 (
        .din(new_Jinkela_wire_168),
        .dout(new_Jinkela_wire_169)
    );

    bfr new_Jinkela_buffer_9 (
        .din(new_Jinkela_wire_8),
        .dout(new_Jinkela_wire_9)
    );

    bfr new_Jinkela_buffer_214 (
        .din(new_Jinkela_wire_241),
        .dout(new_Jinkela_wire_242)
    );

    bfr new_Jinkela_buffer_209 (
        .din(new_Jinkela_wire_234),
        .dout(new_Jinkela_wire_235)
    );

    bfr new_Jinkela_buffer_28 (
        .din(new_Jinkela_wire_31),
        .dout(new_Jinkela_wire_32)
    );

    spl2 new_Jinkela_splitter_13 (
        .a(N102),
        .b(new_Jinkela_wire_238),
        .c(new_Jinkela_wire_239)
    );

    bfr new_Jinkela_buffer_154 (
        .din(new_Jinkela_wire_169),
        .dout(new_Jinkela_wire_170)
    );

    bfr new_Jinkela_buffer_10 (
        .din(new_Jinkela_wire_9),
        .dout(new_Jinkela_wire_10)
    );

    bfr new_Jinkela_buffer_170 (
        .din(new_Jinkela_wire_187),
        .dout(new_Jinkela_wire_188)
    );

    bfr new_Jinkela_buffer_22 (
        .din(new_Jinkela_wire_25),
        .dout(new_Jinkela_wire_26)
    );

    bfr new_Jinkela_buffer_210 (
        .din(new_Jinkela_wire_235),
        .dout(new_Jinkela_wire_236)
    );

    bfr new_Jinkela_buffer_155 (
        .din(new_Jinkela_wire_170),
        .dout(new_Jinkela_wire_171)
    );

    spl2 new_Jinkela_splitter_0 (
        .a(new_Jinkela_wire_10),
        .b(new_Jinkela_wire_11),
        .c(new_Jinkela_wire_12)
    );

    bfr new_Jinkela_buffer_215 (
        .din(new_Jinkela_wire_242),
        .dout(new_Jinkela_wire_243)
    );

    bfr new_Jinkela_buffer_182 (
        .din(new_Jinkela_wire_201),
        .dout(new_Jinkela_wire_202)
    );

    bfr new_Jinkela_buffer_11 (
        .din(new_Jinkela_wire_12),
        .dout(new_Jinkela_wire_13)
    );

    bfr new_Jinkela_buffer_211 (
        .din(new_Jinkela_wire_236),
        .dout(new_Jinkela_wire_237)
    );

    spl2 new_Jinkela_splitter_46 (
        .a(_114_),
        .b(new_Jinkela_wire_749),
        .c(new_Jinkela_wire_750)
    );

    bfr new_Jinkela_buffer_156 (
        .din(new_Jinkela_wire_171),
        .dout(new_Jinkela_wire_172)
    );

    bfr new_Jinkela_buffer_45 (
        .din(new_Jinkela_wire_50),
        .dout(new_Jinkela_wire_51)
    );

    bfr new_Jinkela_buffer_221 (
        .din(new_Jinkela_wire_250),
        .dout(new_Jinkela_wire_251)
    );

    bfr new_Jinkela_buffer_171 (
        .din(new_Jinkela_wire_188),
        .dout(new_Jinkela_wire_189)
    );

    bfr new_Jinkela_buffer_23 (
        .din(new_Jinkela_wire_26),
        .dout(new_Jinkela_wire_27)
    );

    bfr new_Jinkela_buffer_216 (
        .din(new_Jinkela_wire_243),
        .dout(new_Jinkela_wire_244)
    );

    bfr new_Jinkela_buffer_157 (
        .din(new_Jinkela_wire_172),
        .dout(new_Jinkela_wire_173)
    );

    bfr new_Jinkela_buffer_12 (
        .din(new_Jinkela_wire_13),
        .dout(new_Jinkela_wire_14)
    );

    bfr new_Jinkela_buffer_229 (
        .din(new_Jinkela_wire_260),
        .dout(new_Jinkela_wire_261)
    );

    spl2 new_Jinkela_splitter_16 (
        .a(N76),
        .b(new_Jinkela_wire_270),
        .c(new_Jinkela_wire_271)
    );

    bfr new_Jinkela_buffer_188 (
        .din(new_Jinkela_wire_209),
        .dout(new_Jinkela_wire_210)
    );

    bfr new_Jinkela_buffer_29 (
        .din(new_Jinkela_wire_32),
        .dout(new_Jinkela_wire_33)
    );

    bfr new_Jinkela_buffer_217 (
        .din(new_Jinkela_wire_244),
        .dout(new_Jinkela_wire_245)
    );

    bfr new_Jinkela_buffer_172 (
        .din(new_Jinkela_wire_189),
        .dout(new_Jinkela_wire_190)
    );

    bfr new_Jinkela_buffer_13 (
        .din(new_Jinkela_wire_14),
        .dout(new_Jinkela_wire_15)
    );

    bfr new_Jinkela_buffer_222 (
        .din(new_Jinkela_wire_251),
        .dout(new_Jinkela_wire_252)
    );

    bfr new_Jinkela_buffer_183 (
        .din(new_Jinkela_wire_202),
        .dout(new_Jinkela_wire_203)
    );

    bfr new_Jinkela_buffer_24 (
        .din(new_Jinkela_wire_27),
        .dout(new_Jinkela_wire_28)
    );

    bfr new_Jinkela_buffer_218 (
        .din(new_Jinkela_wire_245),
        .dout(new_Jinkela_wire_246)
    );

    bfr new_Jinkela_buffer_173 (
        .din(new_Jinkela_wire_190),
        .dout(new_Jinkela_wire_191)
    );

    bfr new_Jinkela_buffer_14 (
        .din(new_Jinkela_wire_15),
        .dout(new_Jinkela_wire_16)
    );

    bfr new_Jinkela_buffer_246 (
        .din(N99),
        .dout(new_Jinkela_wire_280)
    );

    bfr new_Jinkela_buffer_238 (
        .din(new_Jinkela_wire_271),
        .dout(new_Jinkela_wire_272)
    );

    bfr new_Jinkela_buffer_219 (
        .din(new_Jinkela_wire_246),
        .dout(new_Jinkela_wire_247)
    );

    bfr new_Jinkela_buffer_111 (
        .din(N47),
        .dout(new_Jinkela_wire_123)
    );

    bfr new_Jinkela_buffer_15 (
        .din(new_Jinkela_wire_16),
        .dout(new_Jinkela_wire_17)
    );

    bfr new_Jinkela_buffer_174 (
        .din(new_Jinkela_wire_191),
        .dout(new_Jinkela_wire_192)
    );

    bfr new_Jinkela_buffer_223 (
        .din(new_Jinkela_wire_252),
        .dout(new_Jinkela_wire_253)
    );

    bfr new_Jinkela_buffer_184 (
        .din(new_Jinkela_wire_203),
        .dout(new_Jinkela_wire_204)
    );

    bfr new_Jinkela_buffer_25 (
        .din(new_Jinkela_wire_28),
        .dout(new_Jinkela_wire_29)
    );

    bfr new_Jinkela_buffer_230 (
        .din(new_Jinkela_wire_261),
        .dout(new_Jinkela_wire_262)
    );

    bfr new_Jinkela_buffer_638 (
        .din(new_Jinkela_wire_732),
        .dout(new_Jinkela_wire_733)
    );

    bfr new_Jinkela_buffer_175 (
        .din(new_Jinkela_wire_192),
        .dout(new_Jinkela_wire_193)
    );

    bfr new_Jinkela_buffer_16 (
        .din(new_Jinkela_wire_17),
        .dout(new_Jinkela_wire_18)
    );

    bfr new_Jinkela_buffer_224 (
        .din(new_Jinkela_wire_253),
        .dout(new_Jinkela_wire_254)
    );

    bfr new_Jinkela_buffer_189 (
        .din(new_Jinkela_wire_210),
        .dout(new_Jinkela_wire_211)
    );

    bfr new_Jinkela_buffer_30 (
        .din(new_Jinkela_wire_33),
        .dout(new_Jinkela_wire_34)
    );

    bfr new_Jinkela_buffer_185 (
        .din(new_Jinkela_wire_204),
        .dout(new_Jinkela_wire_205)
    );

    bfr new_Jinkela_buffer_17 (
        .din(new_Jinkela_wire_18),
        .dout(new_Jinkela_wire_19)
    );

    bfr new_Jinkela_buffer_225 (
        .din(new_Jinkela_wire_254),
        .dout(new_Jinkela_wire_255)
    );

    bfr new_Jinkela_buffer_195 (
        .din(new_Jinkela_wire_218),
        .dout(new_Jinkela_wire_219)
    );

    bfr new_Jinkela_buffer_46 (
        .din(new_Jinkela_wire_51),
        .dout(new_Jinkela_wire_52)
    );

    bfr new_Jinkela_buffer_231 (
        .din(new_Jinkela_wire_262),
        .dout(new_Jinkela_wire_263)
    );

    bfr new_Jinkela_buffer_190 (
        .din(new_Jinkela_wire_211),
        .dout(new_Jinkela_wire_212)
    );

    bfr new_Jinkela_buffer_31 (
        .din(new_Jinkela_wire_34),
        .dout(new_Jinkela_wire_35)
    );

    bfr new_Jinkela_buffer_226 (
        .din(new_Jinkela_wire_255),
        .dout(new_Jinkela_wire_256)
    );

    bfr new_Jinkela_buffer_203 (
        .din(new_Jinkela_wire_228),
        .dout(new_Jinkela_wire_229)
    );

    bfr new_Jinkela_buffer_74 (
        .din(new_Jinkela_wire_81),
        .dout(new_Jinkela_wire_82)
    );

    bfr new_Jinkela_buffer_264 (
        .din(N8),
        .dout(new_Jinkela_wire_300)
    );

    spl2 new_Jinkela_splitter_14 (
        .a(N17),
        .b(new_Jinkela_wire_248),
        .c(new_Jinkela_wire_249)
    );

    bfr new_Jinkela_buffer_191 (
        .din(new_Jinkela_wire_212),
        .dout(new_Jinkela_wire_213)
    );

    bfr new_Jinkela_buffer_32 (
        .din(new_Jinkela_wire_35),
        .dout(new_Jinkela_wire_36)
    );

    bfr new_Jinkela_buffer_227 (
        .din(new_Jinkela_wire_256),
        .dout(new_Jinkela_wire_257)
    );

    bfr new_Jinkela_buffer_196 (
        .din(new_Jinkela_wire_219),
        .dout(new_Jinkela_wire_220)
    );

    bfr new_Jinkela_buffer_47 (
        .din(new_Jinkela_wire_52),
        .dout(new_Jinkela_wire_53)
    );

    bfr new_Jinkela_buffer_232 (
        .din(new_Jinkela_wire_263),
        .dout(new_Jinkela_wire_264)
    );

    bfr new_Jinkela_buffer_192 (
        .din(new_Jinkela_wire_213),
        .dout(new_Jinkela_wire_214)
    );

    bfr new_Jinkela_buffer_33 (
        .din(new_Jinkela_wire_36),
        .dout(new_Jinkela_wire_37)
    );

    bfr new_Jinkela_buffer_228 (
        .din(new_Jinkela_wire_257),
        .dout(new_Jinkela_wire_258)
    );

    spl2 new_Jinkela_splitter_19 (
        .a(N11),
        .b(new_Jinkela_wire_320),
        .c(new_Jinkela_wire_321)
    );

    bfr new_Jinkela_buffer_193 (
        .din(new_Jinkela_wire_214),
        .dout(new_Jinkela_wire_215)
    );

    bfr new_Jinkela_buffer_34 (
        .din(new_Jinkela_wire_37),
        .dout(new_Jinkela_wire_38)
    );

    bfr new_Jinkela_buffer_233 (
        .din(new_Jinkela_wire_264),
        .dout(new_Jinkela_wire_265)
    );

    bfr new_Jinkela_buffer_197 (
        .din(new_Jinkela_wire_220),
        .dout(new_Jinkela_wire_221)
    );

    bfr new_Jinkela_buffer_48 (
        .din(new_Jinkela_wire_53),
        .dout(new_Jinkela_wire_54)
    );

    bfr new_Jinkela_buffer_239 (
        .din(new_Jinkela_wire_272),
        .dout(new_Jinkela_wire_273)
    );

    bfr new_Jinkela_buffer_204 (
        .din(new_Jinkela_wire_229),
        .dout(new_Jinkela_wire_230)
    );

    bfr new_Jinkela_buffer_35 (
        .din(new_Jinkela_wire_38),
        .dout(new_Jinkela_wire_39)
    );

    bfr new_Jinkela_buffer_234 (
        .din(new_Jinkela_wire_265),
        .dout(new_Jinkela_wire_266)
    );

    bfr new_Jinkela_buffer_198 (
        .din(new_Jinkela_wire_221),
        .dout(new_Jinkela_wire_222)
    );

    bfr new_Jinkela_buffer_75 (
        .din(new_Jinkela_wire_82),
        .dout(new_Jinkela_wire_83)
    );

    bfr new_Jinkela_buffer_247 (
        .din(new_Jinkela_wire_280),
        .dout(new_Jinkela_wire_281)
    );

    spl2 new_Jinkela_splitter_63 (
        .a(_044_),
        .b(new_Jinkela_wire_903),
        .c(new_Jinkela_wire_904)
    );

    bfr new_Jinkela_buffer_212 (
        .din(new_Jinkela_wire_239),
        .dout(new_Jinkela_wire_240)
    );

    bfr new_Jinkela_buffer_36 (
        .din(new_Jinkela_wire_39),
        .dout(new_Jinkela_wire_40)
    );

    bfr new_Jinkela_buffer_235 (
        .din(new_Jinkela_wire_266),
        .dout(new_Jinkela_wire_267)
    );

    spl2 new_Jinkela_splitter_15 (
        .a(N50),
        .b(new_Jinkela_wire_259),
        .c(new_Jinkela_wire_260)
    );

    bfr new_Jinkela_buffer_199 (
        .din(new_Jinkela_wire_222),
        .dout(new_Jinkela_wire_223)
    );

    bfr new_Jinkela_buffer_49 (
        .din(new_Jinkela_wire_54),
        .dout(new_Jinkela_wire_55)
    );

    bfr new_Jinkela_buffer_240 (
        .din(new_Jinkela_wire_273),
        .dout(new_Jinkela_wire_274)
    );

    bfr new_Jinkela_buffer_205 (
        .din(new_Jinkela_wire_230),
        .dout(new_Jinkela_wire_231)
    );

    spl2 new_Jinkela_splitter_2 (
        .a(new_Jinkela_wire_40),
        .b(new_Jinkela_wire_41),
        .c(new_Jinkela_wire_42)
    );

    bfr new_Jinkela_buffer_236 (
        .din(new_Jinkela_wire_267),
        .dout(new_Jinkela_wire_268)
    );

    bfr new_Jinkela_buffer_759 (
        .din(new_Jinkela_wire_892),
        .dout(new_Jinkela_wire_893)
    );

    bfr new_Jinkela_buffer_200 (
        .din(new_Jinkela_wire_223),
        .dout(new_Jinkela_wire_224)
    );

    bfr new_Jinkela_buffer_37 (
        .din(new_Jinkela_wire_42),
        .dout(new_Jinkela_wire_43)
    );

    bfr new_Jinkela_buffer_290 (
        .din(N21),
        .dout(new_Jinkela_wire_330)
    );

    bfr new_Jinkela_buffer_241 (
        .din(new_Jinkela_wire_274),
        .dout(new_Jinkela_wire_275)
    );

    bfr new_Jinkela_buffer_102 (
        .din(new_Jinkela_wire_113),
        .dout(new_Jinkela_wire_114)
    );

    bfr new_Jinkela_buffer_220 (
        .din(new_Jinkela_wire_249),
        .dout(new_Jinkela_wire_250)
    );

    bfr new_Jinkela_buffer_129 (
        .din(N79),
        .dout(new_Jinkela_wire_143)
    );

    bfr new_Jinkela_buffer_745 (
        .din(new_Jinkela_wire_876),
        .dout(new_Jinkela_wire_877)
    );

    bfr new_Jinkela_buffer_201 (
        .din(new_Jinkela_wire_224),
        .dout(new_Jinkela_wire_225)
    );

    bfr new_Jinkela_buffer_248 (
        .din(new_Jinkela_wire_281),
        .dout(new_Jinkela_wire_282)
    );

    bfr new_Jinkela_buffer_50 (
        .din(new_Jinkela_wire_55),
        .dout(new_Jinkela_wire_56)
    );

    bfr new_Jinkela_buffer_444 (
        .din(new_Jinkela_wire_495),
        .dout(new_Jinkela_wire_496)
    );

    bfr new_Jinkela_buffer_706 (
        .din(new_Jinkela_wire_831),
        .dout(new_Jinkela_wire_832)
    );

    bfr new_Jinkela_buffer_347 (
        .din(new_Jinkela_wire_392),
        .dout(new_Jinkela_wire_393)
    );

    bfr new_Jinkela_buffer_426 (
        .din(new_Jinkela_wire_477),
        .dout(new_Jinkela_wire_478)
    );

    bfr new_Jinkela_buffer_322 (
        .din(new_Jinkela_wire_365),
        .dout(new_Jinkela_wire_366)
    );

    bfr new_Jinkela_buffer_707 (
        .din(new_Jinkela_wire_832),
        .dout(new_Jinkela_wire_833)
    );

    spl2 new_Jinkela_splitter_31 (
        .a(N37),
        .b(new_Jinkela_wire_589),
        .c(new_Jinkela_wire_590)
    );

    bfr new_Jinkela_buffer_340 (
        .din(new_Jinkela_wire_385),
        .dout(new_Jinkela_wire_386)
    );

    bfr new_Jinkela_buffer_427 (
        .din(new_Jinkela_wire_478),
        .dout(new_Jinkela_wire_479)
    );

    bfr new_Jinkela_buffer_323 (
        .din(new_Jinkela_wire_366),
        .dout(new_Jinkela_wire_367)
    );

    bfr new_Jinkela_buffer_715 (
        .din(new_Jinkela_wire_840),
        .dout(new_Jinkela_wire_841)
    );

    bfr new_Jinkela_buffer_445 (
        .din(new_Jinkela_wire_496),
        .dout(new_Jinkela_wire_497)
    );

    bfr new_Jinkela_buffer_708 (
        .din(new_Jinkela_wire_833),
        .dout(new_Jinkela_wire_834)
    );

    bfr new_Jinkela_buffer_428 (
        .din(new_Jinkela_wire_479),
        .dout(new_Jinkela_wire_480)
    );

    bfr new_Jinkela_buffer_324 (
        .din(new_Jinkela_wire_367),
        .dout(new_Jinkela_wire_368)
    );

    bfr new_Jinkela_buffer_718 (
        .din(new_Jinkela_wire_847),
        .dout(new_Jinkela_wire_848)
    );

    bfr new_Jinkela_buffer_468 (
        .din(new_Jinkela_wire_521),
        .dout(new_Jinkela_wire_522)
    );

    bfr new_Jinkela_buffer_709 (
        .din(new_Jinkela_wire_834),
        .dout(new_Jinkela_wire_835)
    );

    bfr new_Jinkela_buffer_433 (
        .din(N14),
        .dout(new_Jinkela_wire_485)
    );

    bfr new_Jinkela_buffer_341 (
        .din(new_Jinkela_wire_386),
        .dout(new_Jinkela_wire_387)
    );

    bfr new_Jinkela_buffer_429 (
        .din(new_Jinkela_wire_480),
        .dout(new_Jinkela_wire_481)
    );

    bfr new_Jinkela_buffer_325 (
        .din(new_Jinkela_wire_368),
        .dout(new_Jinkela_wire_369)
    );

    bfr new_Jinkela_buffer_716 (
        .din(new_Jinkela_wire_841),
        .dout(new_Jinkela_wire_842)
    );

    bfr new_Jinkela_buffer_446 (
        .din(new_Jinkela_wire_497),
        .dout(new_Jinkela_wire_498)
    );

    bfr new_Jinkela_buffer_710 (
        .din(new_Jinkela_wire_835),
        .dout(new_Jinkela_wire_836)
    );

    bfr new_Jinkela_buffer_348 (
        .din(new_Jinkela_wire_393),
        .dout(new_Jinkela_wire_394)
    );

    bfr new_Jinkela_buffer_430 (
        .din(new_Jinkela_wire_481),
        .dout(new_Jinkela_wire_482)
    );

    bfr new_Jinkela_buffer_326 (
        .din(new_Jinkela_wire_369),
        .dout(new_Jinkela_wire_370)
    );

    bfr new_Jinkela_buffer_735 (
        .din(_050_),
        .dout(new_Jinkela_wire_867)
    );

    bfr new_Jinkela_buffer_494 (
        .din(new_Jinkela_wire_549),
        .dout(new_Jinkela_wire_550)
    );

    bfr new_Jinkela_buffer_711 (
        .din(new_Jinkela_wire_836),
        .dout(new_Jinkela_wire_837)
    );

    bfr new_Jinkela_buffer_342 (
        .din(new_Jinkela_wire_387),
        .dout(new_Jinkela_wire_388)
    );

    bfr new_Jinkela_buffer_431 (
        .din(new_Jinkela_wire_482),
        .dout(new_Jinkela_wire_483)
    );

    bfr new_Jinkela_buffer_327 (
        .din(new_Jinkela_wire_370),
        .dout(new_Jinkela_wire_371)
    );

    bfr new_Jinkela_buffer_717 (
        .din(new_Jinkela_wire_842),
        .dout(new_Jinkela_wire_843)
    );

    bfr new_Jinkela_buffer_447 (
        .din(new_Jinkela_wire_498),
        .dout(new_Jinkela_wire_499)
    );

    bfr new_Jinkela_buffer_376 (
        .din(new_Jinkela_wire_423),
        .dout(new_Jinkela_wire_424)
    );

    bfr new_Jinkela_buffer_432 (
        .din(new_Jinkela_wire_483),
        .dout(new_Jinkela_wire_484)
    );

    bfr new_Jinkela_buffer_719 (
        .din(new_Jinkela_wire_848),
        .dout(new_Jinkela_wire_849)
    );

    bfr new_Jinkela_buffer_328 (
        .din(new_Jinkela_wire_371),
        .dout(new_Jinkela_wire_372)
    );

    bfr new_Jinkela_buffer_767 (
        .din(new_Jinkela_wire_904),
        .dout(new_Jinkela_wire_905)
    );

    bfr new_Jinkela_buffer_469 (
        .din(new_Jinkela_wire_522),
        .dout(new_Jinkela_wire_523)
    );

    bfr new_Jinkela_buffer_727 (
        .din(new_Jinkela_wire_858),
        .dout(new_Jinkela_wire_859)
    );

    bfr new_Jinkela_buffer_736 (
        .din(new_net_196),
        .dout(new_Jinkela_wire_868)
    );

    bfr new_Jinkela_buffer_343 (
        .din(new_Jinkela_wire_388),
        .dout(new_Jinkela_wire_389)
    );

    bfr new_Jinkela_buffer_448 (
        .din(new_Jinkela_wire_499),
        .dout(new_Jinkela_wire_500)
    );

    bfr new_Jinkela_buffer_720 (
        .din(new_Jinkela_wire_849),
        .dout(new_Jinkela_wire_850)
    );

    bfr new_Jinkela_buffer_329 (
        .din(new_Jinkela_wire_372),
        .dout(new_Jinkela_wire_373)
    );

    bfr new_Jinkela_buffer_760 (
        .din(new_Jinkela_wire_893),
        .dout(new_Jinkela_wire_894)
    );

    bfr new_Jinkela_buffer_738 (
        .din(new_net_194),
        .dout(new_Jinkela_wire_870)
    );

    bfr new_Jinkela_buffer_349 (
        .din(new_Jinkela_wire_394),
        .dout(new_Jinkela_wire_395)
    );

    bfr new_Jinkela_buffer_449 (
        .din(new_Jinkela_wire_500),
        .dout(new_Jinkela_wire_501)
    );

    bfr new_Jinkela_buffer_721 (
        .din(new_Jinkela_wire_850),
        .dout(new_Jinkela_wire_851)
    );

    bfr new_Jinkela_buffer_330 (
        .din(new_Jinkela_wire_373),
        .dout(new_Jinkela_wire_374)
    );

    bfr new_Jinkela_buffer_470 (
        .din(new_Jinkela_wire_523),
        .dout(new_Jinkela_wire_524)
    );

    bfr new_Jinkela_buffer_728 (
        .din(new_Jinkela_wire_859),
        .dout(new_Jinkela_wire_860)
    );

    bfr new_Jinkela_buffer_747 (
        .din(new_Jinkela_wire_878),
        .dout(new_Jinkela_wire_879)
    );

    bfr new_Jinkela_buffer_344 (
        .din(new_Jinkela_wire_389),
        .dout(new_Jinkela_wire_390)
    );

    bfr new_Jinkela_buffer_450 (
        .din(new_Jinkela_wire_501),
        .dout(new_Jinkela_wire_502)
    );

    bfr new_Jinkela_buffer_722 (
        .din(new_Jinkela_wire_851),
        .dout(new_Jinkela_wire_852)
    );

    bfr new_Jinkela_buffer_331 (
        .din(new_Jinkela_wire_374),
        .dout(new_Jinkela_wire_375)
    );

    bfr new_Jinkela_buffer_652 (
        .din(new_Jinkela_wire_750),
        .dout(new_Jinkela_wire_751)
    );

    bfr new_Jinkela_buffer_495 (
        .din(new_Jinkela_wire_550),
        .dout(new_Jinkela_wire_551)
    );

    bfr new_Jinkela_buffer_737 (
        .din(new_Jinkela_wire_868),
        .dout(new_Jinkela_wire_869)
    );

    bfr new_Jinkela_buffer_451 (
        .din(new_Jinkela_wire_502),
        .dout(new_Jinkela_wire_503)
    );

    bfr new_Jinkela_buffer_723 (
        .din(new_Jinkela_wire_852),
        .dout(new_Jinkela_wire_853)
    );

    bfr new_Jinkela_buffer_332 (
        .din(new_Jinkela_wire_375),
        .dout(new_Jinkela_wire_376)
    );

    bfr new_Jinkela_buffer_471 (
        .din(new_Jinkela_wire_524),
        .dout(new_Jinkela_wire_525)
    );

    bfr new_Jinkela_buffer_661 (
        .din(new_Jinkela_wire_761),
        .dout(new_Jinkela_wire_762)
    );

    bfr new_Jinkela_buffer_729 (
        .din(new_Jinkela_wire_860),
        .dout(new_Jinkela_wire_861)
    );

    bfr new_Jinkela_buffer_462 (
        .din(N105),
        .dout(new_Jinkela_wire_516)
    );

    bfr new_Jinkela_buffer_345 (
        .din(new_Jinkela_wire_390),
        .dout(new_Jinkela_wire_391)
    );

    bfr new_Jinkela_buffer_452 (
        .din(new_Jinkela_wire_503),
        .dout(new_Jinkela_wire_504)
    );

    bfr new_Jinkela_buffer_724 (
        .din(new_Jinkela_wire_853),
        .dout(new_Jinkela_wire_854)
    );

    bfr new_Jinkela_buffer_333 (
        .din(new_Jinkela_wire_376),
        .dout(new_Jinkela_wire_377)
    );

    bfr new_Jinkela_buffer_510 (
        .din(new_Jinkela_wire_569),
        .dout(new_Jinkela_wire_570)
    );

    spl2 new_Jinkela_splitter_61 (
        .a(_081_),
        .b(new_Jinkela_wire_889),
        .c(new_Jinkela_wire_890)
    );

    bfr new_Jinkela_buffer_350 (
        .din(new_Jinkela_wire_395),
        .dout(new_Jinkela_wire_396)
    );

    bfr new_Jinkela_buffer_453 (
        .din(new_Jinkela_wire_504),
        .dout(new_Jinkela_wire_505)
    );

    bfr new_Jinkela_buffer_725 (
        .din(new_Jinkela_wire_854),
        .dout(new_Jinkela_wire_855)
    );

    bfr new_Jinkela_buffer_334 (
        .din(new_Jinkela_wire_377),
        .dout(new_Jinkela_wire_378)
    );

    bfr new_Jinkela_buffer_472 (
        .din(new_Jinkela_wire_525),
        .dout(new_Jinkela_wire_526)
    );

    bfr new_Jinkela_buffer_730 (
        .din(new_Jinkela_wire_861),
        .dout(new_Jinkela_wire_862)
    );

    bfr new_Jinkela_buffer_377 (
        .din(new_Jinkela_wire_424),
        .dout(new_Jinkela_wire_425)
    );

    spl2 new_Jinkela_splitter_26 (
        .a(new_Jinkela_wire_505),
        .b(new_Jinkela_wire_506),
        .c(new_Jinkela_wire_507)
    );

    bfr new_Jinkela_buffer_726 (
        .din(new_Jinkela_wire_855),
        .dout(new_Jinkela_wire_856)
    );

    bfr new_Jinkela_buffer_335 (
        .din(new_Jinkela_wire_378),
        .dout(new_Jinkela_wire_379)
    );

    bfr new_Jinkela_buffer_454 (
        .din(new_Jinkela_wire_507),
        .dout(new_Jinkela_wire_508)
    );

    bfr new_Jinkela_buffer_748 (
        .din(new_Jinkela_wire_879),
        .dout(new_Jinkela_wire_880)
    );

    spl2 new_Jinkela_splitter_62 (
        .a(_037_),
        .b(new_Jinkela_wire_899),
        .c(new_Jinkela_wire_900)
    );

    bfr new_Jinkela_buffer_739 (
        .din(new_Jinkela_wire_870),
        .dout(new_Jinkela_wire_871)
    );

    bfr new_Jinkela_buffer_351 (
        .din(new_Jinkela_wire_396),
        .dout(new_Jinkela_wire_397)
    );

    bfr new_Jinkela_buffer_496 (
        .din(new_Jinkela_wire_551),
        .dout(new_Jinkela_wire_552)
    );

    bfr new_Jinkela_buffer_731 (
        .din(new_Jinkela_wire_862),
        .dout(new_Jinkela_wire_863)
    );

    bfr new_Jinkela_buffer_336 (
        .din(new_Jinkela_wire_379),
        .dout(new_Jinkela_wire_380)
    );

    bfr new_Jinkela_buffer_0 (
        .din(N86),
        .dout(new_Jinkela_wire_0)
    );

    bfr new_Jinkela_buffer_473 (
        .din(new_Jinkela_wire_526),
        .dout(new_Jinkela_wire_527)
    );

    bfr new_Jinkela_buffer_757 (
        .din(new_Jinkela_wire_890),
        .dout(new_Jinkela_wire_891)
    );

    spl2 new_Jinkela_splitter_1 (
        .a(N69),
        .b(new_Jinkela_wire_20),
        .c(new_Jinkela_wire_21)
    );

    bfr new_Jinkela_buffer_405 (
        .din(new_Jinkela_wire_454),
        .dout(new_Jinkela_wire_455)
    );

    bfr new_Jinkela_buffer_455 (
        .din(new_Jinkela_wire_508),
        .dout(new_Jinkela_wire_509)
    );

    bfr new_Jinkela_buffer_26 (
        .din(N34),
        .dout(new_Jinkela_wire_30)
    );

    bfr new_Jinkela_buffer_337 (
        .din(new_Jinkela_wire_380),
        .dout(new_Jinkela_wire_381)
    );

    bfr new_Jinkela_buffer_732 (
        .din(new_Jinkela_wire_863),
        .dout(new_Jinkela_wire_864)
    );

    bfr new_Jinkela_buffer_1 (
        .din(new_Jinkela_wire_0),
        .dout(new_Jinkela_wire_1)
    );

    bfr new_Jinkela_buffer_518 (
        .din(new_Jinkela_wire_579),
        .dout(new_Jinkela_wire_580)
    );

    bfr new_Jinkela_buffer_535 (
        .din(N112),
        .dout(new_Jinkela_wire_599)
    );

    bfr new_Jinkela_buffer_740 (
        .din(new_Jinkela_wire_871),
        .dout(new_Jinkela_wire_872)
    );

    bfr new_Jinkela_buffer_352 (
        .din(new_Jinkela_wire_397),
        .dout(new_Jinkela_wire_398)
    );

    bfr new_Jinkela_buffer_456 (
        .din(new_Jinkela_wire_509),
        .dout(new_Jinkela_wire_510)
    );

    bfr new_Jinkela_buffer_733 (
        .din(new_Jinkela_wire_864),
        .dout(new_Jinkela_wire_865)
    );

    bfr new_Jinkela_buffer_2 (
        .din(new_Jinkela_wire_1),
        .dout(new_Jinkela_wire_2)
    );

    bfr new_Jinkela_buffer_378 (
        .din(new_Jinkela_wire_425),
        .dout(new_Jinkela_wire_426)
    );

    bfr new_Jinkela_buffer_474 (
        .din(new_Jinkela_wire_527),
        .dout(new_Jinkela_wire_528)
    );

    bfr new_Jinkela_buffer_18 (
        .din(new_Jinkela_wire_21),
        .dout(new_Jinkela_wire_22)
    );

    bfr new_Jinkela_buffer_353 (
        .din(new_Jinkela_wire_398),
        .dout(new_Jinkela_wire_399)
    );

    bfr new_Jinkela_buffer_457 (
        .din(new_Jinkela_wire_510),
        .dout(new_Jinkela_wire_511)
    );

    bfr new_Jinkela_buffer_44 (
        .din(N92),
        .dout(new_Jinkela_wire_50)
    );

    bfr new_Jinkela_buffer_734 (
        .din(new_Jinkela_wire_865),
        .dout(new_Jinkela_wire_866)
    );

    bfr new_Jinkela_buffer_761 (
        .din(new_Jinkela_wire_894),
        .dout(new_Jinkela_wire_895)
    );

    bfr new_Jinkela_buffer_3 (
        .din(new_Jinkela_wire_2),
        .dout(new_Jinkela_wire_3)
    );

    bfr new_Jinkela_buffer_497 (
        .din(new_Jinkela_wire_552),
        .dout(new_Jinkela_wire_553)
    );

    bfr new_Jinkela_buffer_766 (
        .din(_115_),
        .dout(new_Jinkela_wire_902)
    );

    bfr new_Jinkela_buffer_491 (
        .din(N60),
        .dout(new_Jinkela_wire_547)
    );

    bfr new_Jinkela_buffer_741 (
        .din(new_Jinkela_wire_872),
        .dout(new_Jinkela_wire_873)
    );

    bfr new_Jinkela_buffer_354 (
        .din(new_Jinkela_wire_399),
        .dout(new_Jinkela_wire_400)
    );

    bfr new_Jinkela_buffer_458 (
        .din(new_Jinkela_wire_511),
        .dout(new_Jinkela_wire_512)
    );

    bfr new_Jinkela_buffer_73 (
        .din(N27),
        .dout(new_Jinkela_wire_81)
    );

    bfr new_Jinkela_buffer_765 (
        .din(new_Jinkela_wire_900),
        .dout(new_Jinkela_wire_901)
    );

    bfr new_Jinkela_buffer_4 (
        .din(new_Jinkela_wire_3),
        .dout(new_Jinkela_wire_4)
    );

    bfr new_Jinkela_buffer_379 (
        .din(new_Jinkela_wire_426),
        .dout(new_Jinkela_wire_427)
    );

    bfr new_Jinkela_buffer_475 (
        .din(new_Jinkela_wire_528),
        .dout(new_Jinkela_wire_529)
    );

    bfr new_Jinkela_buffer_742 (
        .din(new_Jinkela_wire_873),
        .dout(new_Jinkela_wire_874)
    );

    bfr new_Jinkela_buffer_19 (
        .din(new_Jinkela_wire_22),
        .dout(new_Jinkela_wire_23)
    );

    bfr new_Jinkela_buffer_355 (
        .din(new_Jinkela_wire_400),
        .dout(new_Jinkela_wire_401)
    );

    bfr new_Jinkela_buffer_459 (
        .din(new_Jinkela_wire_512),
        .dout(new_Jinkela_wire_513)
    );

    or_ii _163_ (
        .a(_106_),
        .b(new_Jinkela_wire_122),
        .c(_107_)
    );

    bfr new_Jinkela_buffer_5 (
        .din(new_Jinkela_wire_4),
        .dout(new_Jinkela_wire_5)
    );

    bfr new_Jinkela_buffer_406 (
        .din(new_Jinkela_wire_455),
        .dout(new_Jinkela_wire_456)
    );

    bfr new_Jinkela_buffer_511 (
        .din(new_Jinkela_wire_570),
        .dout(new_Jinkela_wire_571)
    );

    bfr new_Jinkela_buffer_743 (
        .din(new_Jinkela_wire_874),
        .dout(new_Jinkela_wire_875)
    );

    bfr new_Jinkela_buffer_758 (
        .din(new_Jinkela_wire_891),
        .dout(new_Jinkela_wire_892)
    );

    bfr new_Jinkela_buffer_27 (
        .din(new_Jinkela_wire_30),
        .dout(new_Jinkela_wire_31)
    );

    bfr new_Jinkela_buffer_356 (
        .din(new_Jinkela_wire_401),
        .dout(new_Jinkela_wire_402)
    );

    bfr new_Jinkela_buffer_460 (
        .din(new_Jinkela_wire_513),
        .dout(new_Jinkela_wire_514)
    );

    bfr new_Jinkela_buffer_815 (
        .din(new_Jinkela_wire_964),
        .dout(new_Jinkela_wire_965)
    );

    bfr new_Jinkela_buffer_820 (
        .din(new_Jinkela_wire_984),
        .dout(new_Jinkela_wire_985)
    );

    bfr new_Jinkela_buffer_777 (
        .din(_092_),
        .dout(new_Jinkela_wire_917)
    );

    bfr new_Jinkela_buffer_821 (
        .din(new_Jinkela_wire_985),
        .dout(new_Jinkela_wire_986)
    );

    bfr new_Jinkela_buffer_822 (
        .din(new_Jinkela_wire_986),
        .dout(new_Jinkela_wire_987)
    );

    bfr new_Jinkela_buffer_823 (
        .din(new_Jinkela_wire_987),
        .dout(new_Jinkela_wire_988)
    );

    bfr new_Jinkela_buffer_769 (
        .din(new_Jinkela_wire_908),
        .dout(new_Jinkela_wire_909)
    );

    bfr new_Jinkela_buffer_824 (
        .din(new_Jinkela_wire_988),
        .dout(new_Jinkela_wire_989)
    );

    bfr new_Jinkela_buffer_650 (
        .din(new_Jinkela_wire_746),
        .dout(new_Jinkela_wire_747)
    );

    bfr new_Jinkela_buffer_825 (
        .din(new_Jinkela_wire_989),
        .dout(new_Jinkela_wire_990)
    );

    bfr new_Jinkela_buffer_762 (
        .din(new_Jinkela_wire_895),
        .dout(new_Jinkela_wire_896)
    );

    bfr new_Jinkela_buffer_826 (
        .din(new_Jinkela_wire_990),
        .dout(new_Jinkela_wire_991)
    );

    bfr new_Jinkela_buffer_751 (
        .din(new_Jinkela_wire_882),
        .dout(new_Jinkela_wire_883)
    );

    and_bi _142_ (
        .a(_082_),
        .b(_085_),
        .c(_086_)
    );

    and_bi _120_ (
        .a(new_Jinkela_wire_567),
        .b(new_Jinkela_wire_206),
        .c(_064_)
    );

    and_bi _118_ (
        .a(new_Jinkela_wire_195),
        .b(new_Jinkela_wire_238),
        .c(_062_)
    );

    and_bi _119_ (
        .a(new_Jinkela_wire_728),
        .b(new_Jinkela_wire_818),
        .c(_063_)
    );

    or_bi _117_ (
        .a(new_Jinkela_wire_194),
        .b(new_Jinkela_wire_350),
        .c(_061_)
    );

    and_bi _121_ (
        .a(new_Jinkela_wire_578),
        .b(new_Jinkela_wire_382),
        .c(_065_)
    );

    and_bi _125_ (
        .a(new_Jinkela_wire_20),
        .b(new_Jinkela_wire_269),
        .c(_069_)
    );

    or_bb _124_ (
        .a(_067_),
        .b(new_Jinkela_wire_737),
        .c(_068_)
    );

    and_bi _122_ (
        .a(new_Jinkela_wire_216),
        .b(new_Jinkela_wire_270),
        .c(_066_)
    );

    or_ii _134_ (
        .a(new_Jinkela_wire_973),
        .b(new_Jinkela_wire_359),
        .c(_078_)
    );

    bfr new_Jinkela_buffer_752 (
        .din(new_Jinkela_wire_883),
        .dout(new_Jinkela_wire_884)
    );

    or_bb _123_ (
        .a(_066_),
        .b(_065_),
        .c(_067_)
    );

    and_bi _126_ (
        .a(new_Jinkela_wire_112),
        .b(new_Jinkela_wire_589),
        .c(_070_)
    );

    or_bb _127_ (
        .a(new_Jinkela_wire_666),
        .b(new_Jinkela_wire_667),
        .c(_071_)
    );

    and_bi _128_ (
        .a(new_Jinkela_wire_227),
        .b(new_Jinkela_wire_259),
        .c(_072_)
    );

    and_bi _129_ (
        .a(new_Jinkela_wire_248),
        .b(new_Jinkela_wire_320),
        .c(_073_)
    );

    or_bb _130_ (
        .a(_073_),
        .b(_072_),
        .c(_074_)
    );

    or_bb _131_ (
        .a(new_Jinkela_wire_738),
        .b(_071_),
        .c(_075_)
    );

    or_bb _132_ (
        .a(_075_),
        .b(new_Jinkela_wire_775),
        .c(_076_)
    );

    bfr new_Jinkela_buffer_763 (
        .din(new_Jinkela_wire_896),
        .dout(new_Jinkela_wire_897)
    );

    and_bi _133_ (
        .a(new_Jinkela_wire_800),
        .b(_076_),
        .c(_077_)
    );

    and_bb _135_ (
        .a(_078_),
        .b(new_Jinkela_wire_736),
        .c(_079_)
    );

    bfr new_Jinkela_buffer_753 (
        .din(new_Jinkela_wire_884),
        .dout(new_Jinkela_wire_885)
    );

    or_bi _136_ (
        .a(new_Jinkela_wire_979),
        .b(new_Jinkela_wire_247),
        .c(_080_)
    );

    or_ii _137_ (
        .a(_080_),
        .b(new_Jinkela_wire_205),
        .c(_081_)
    );

    or_bb _138_ (
        .a(new_Jinkela_wire_889),
        .b(new_Jinkela_wire_610),
        .c(_082_)
    );

    or_bi _139_ (
        .a(new_Jinkela_wire_975),
        .b(new_Jinkela_wire_279),
        .c(_083_)
    );

    or_ii _140_ (
        .a(_083_),
        .b(new_Jinkela_wire_226),
        .c(_084_)
    );

    and_ii _141_ (
        .a(new_Jinkela_wire_789),
        .b(new_Jinkela_wire_11),
        .c(_085_)
    );

endmodule
